��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��.�2ָi1f�Rןx5~?��77`*����V5�[%�W��[+
.�������S��Vz�!a�Vx�� j���ͳ-��e�y�U�5�0��!�%�D~K� �S��T(��]��DA�E�J�q����T���� ���oѨ�p��0#;pqp�4�yX���0�U�1������	�Yt���a�xl
Gd�},�Y����ӣE>@ůX#pa(]Ȥ����g"]wQ��U�] O1���2���.���dؐ����X�E�DY����4�ah�Xj�Nݔ��Ur-W��,B��Q�o��,Q�O������ĺx�&���Ak�c�&�P�^?]~r7��?������e$��?>� d�Q���x��$�
u��5��8�h7��LY�w�s�2ޏ���.CT�:�g^���B(����{��4+j�=7s�����!�]e����Jf�d�bS �9D{,2c��_�ʲ���數�A�I�	tA����6�w�`B�\�
{��2{� �{��&ۧ�9$�WF��OⵗM
=�Mv{�+\,���?=�a��H��M�@y~	YHu�:�;�N�׿�U�&l>�9�7�^1c���J�4y�v��6��*jݔO����Z ����!CL�w��h\��y=����}��ϫ��D�{�N퉾<��V�G�4��P�1\�Q4�P�{��V ���?�l�o�f��-��J��Y�a-3��ne�M�!,�B��>�1���O��w���۹�U%P�H�Q_�¶UM
3�o��FR�?�����<�.C���.]I���c���L/h�����Y �+�P�H��G}L�䦟�0r���g�cv.�D��9A��$�����9^YQ�C)XpŘ��@$$k������>-�-In�C���V��-�����V��kxcM�^��-��X���em9�+��s�r��X���N���*���'���8�=�ͫh᥉�J�M�'�X��4�Ti��-yAL�o�8�^�?�E�I�)W`����Z-��v����*����A����K�ͮ�B��3�X̴�TV<��h6�p�|AMN�"�s��#�I#l;]��1T����w���O��ۓ;m��U�5� *5w��� �y���>i�����m�p��v/�Ras�D��u?
�LF�N�f�j}�_�b�`qI%[�$Y��F���8�0�`�^�U�F��Q,0>�Bݘ��{��'SĶ�)����D���M�Z�S��|T&�r��n�����[�;q�����7���8�̆'b>yޙ�
�Λ-CH8S�@+c��Ǧ����&i|�*AI˒.�c_=(t)�5�ƴ;:Y8�d��+�m�घ	��!S���uDnJ�b����I�7�E�.�����Y���I����B<�x�_�xH$w�=��B.n/���i�b4��7*��"��(A��Ҙ��	A_D�E���W?j		Q����Y�[��*�����="�%�G6ʌY5ls,��ŕd+��Uw�֗��~����*��'f츅�28as��S�����S��E=��\�<`/�Uc�D�4Y�;� �P`0��"[���,�
�A�+��7N��i�����9�{��숱&������������w:NE�߱̑q�+7�p��������홧2�)GZလ'�!������x�Y�y?6>���({r�4���ǁ�_%i�RV�U ���@���L��E�g��;�T6O����>�<�����uK�j�9�qWVa�<O���I�=¼U�H-�'I�Ef����t�M��8A��e�jF���̈��9��B�B'����G�w>l�.�3�tse(^��:�Yȶ���49²�F�@Tyt�8�@c:	�s���g�o�X�-�3`8��6<��9�m̸@��^��G�^�'�u��/���+Z��.~�2�cDm�IL�D��2��x4+�(V��7S8 A`��������Yxᣠ\&���_���C�va�Sf�iP�6[28�a�܀+]$qa�i�� �zO�D�ؚ���:�
�����(S[i@bT����B")��X�=Ɵ�@q�,��B	�L��;�� �M��<���h���b��l滖*s�(G뇮�G���ӡ��Żn���E�&�.�nA+:���噫p�*�g�����F�9��p �ݺJ����Wďqb��Qr�՚��������F�� �o2n�^X5�=�8���o����7B)0� 	&��?�n��U�;�tu�`����d^����0h��E@1+�����*����H~��|��s;�ѡ��'��jD��A�M�fl��>�04Z8S�AA<�ߑAi��d�Č��������N���t�
�`6����#����X1���"�Ka,yz�cל_ҫ�9����J�֛�԰%��U��!B��?����'�q>�_��L�����G�/�؂��Us��MP���f6��EFՎES�J���_�]SM������z��
�-�BV��uxն��~*�d���RN���>q��H1Y�����m��Ǎq�\�vZ��Om�N6��y��0�Z�T͂%N��@��ԇ�y��JW�N�;������p�i��̵�]��9�6%���+o�t�#��֙-mm���p�]g>��'�1��:�,�V`[��t��A�O��@H�^R�3��G�/���Dհ�|�\�:3���E���m~>r��9�®����_k;Q�9�Н�ؾ7��@p��n�Ş,~���i5�RN��J����d�ζ�{�MI�Y�