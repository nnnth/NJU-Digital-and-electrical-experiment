��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��H�2��M*e�b��a�/\�?hcVU�թ0�{��:�����=N����TV8�㥔i �jV������[-���NC%��Jga��������%%�rhp�;
!��/�������'�YU��։����b�/�0���<L;�-����i�нC��.Yg��g��s8�Smcj�^�/�3�'��l��ykm&�=�s�ۼ�;������<L��̛p^�<�u����*�A};E��sz2=�y�_S���N&H�45/�������7NQ<��-�;�>bQW�%�x�U��22����#��Z\�KHW��^qT't���2��,=}y������g�n�֯���r�$��`�׻��{l�L�������&?��iLZ����f=H�"�0���_c�C�qj��BVX����py#-��<��J K+�&Wov����F�/��㵱��.k_"@<�у5��T	w��<���(;����G��Ta���,B��E���Hwq��t>M����c�`3Ǐ���������v �������F�7ַS M��ZǪ��W}�ި�ݢQ��U$s��l�H��Ov����,�b
Ҵ���Y�b���%(�����}{�l`#�p���6A�@le@Sq�����Vk����S�G٤I-v=�2}t0��c�t�_j4&о���Ӆ/�Kw��UJO��\��zy�Vy��$%�SZ�|d2�t�Y����'w��}�_B!�q���3�F��t�@�(�*:����]�|�1+��p=%��#���u�A��,&��y�bz���g��� tG�� X�k*Xϕo�4>�`i0KE:B(�D�s5Q׽�8��Ȱ�t)wiE�|��d2��S��7�W'�4v���񚫥���H��iV�j�������tp�"��)�b>�h����.�b��]�`��S�g�J{�T�;,*l���@��l��mKw-���
�-~5>�Y��&�JĪ;[��X��˙1[2d�|����;	,��k/~-.5��Fg2��c�Jw �Rh@��O|�C,$���W����^�=�h��7\�ꯟ?�~�A������ׁ�'G(^��Og���hP��a:��"��T����$�CIz���P�U�cU!�2�4Ut%���)}hŖ��J�dQO�KZ�u��Ρ\���#2�����f��8�L�7[~y��x�JQG�}�©�;k��yC-���zn�s�>h��V��V���\X"[Hh ���?s�I�<��V0ĸ%@�ts��aFm,$r�i�T���}Ug��&@N�vV�`6GI|?~����W �9
lȨ��LkT�=�%�ʮ���?RdD��3��j���#��7�R�cY���Y9?>�I���hΦ8�`�{��I��<�5�JRE���B��p���ճbG'���+�5V���!^8�N��y��S�C'��h=tSģ2Oe�^]�9!�F�b��(��';g���	\��]S���g���]o��k�cz����n�>/��w+V�%�e����W>�=������1{��F��x��C@��+$<2g��0���,��tw s��,���P[O�B�aTEy��y:�=,9�C��75�'�M(N���g����P�Cd��?�Ԉ�A��3LVR[�ܴӻ�w\��c����㺳Z��p="H�Kp�K�(K2T���>t����7��T���j����x��Y{�0�oVZF�t&�&v	z��aZ�!c�= ��R-T>�3��� ;&�BE�Kal�P+G/���dܞ����_sK�Q�����B�
E�<��3�EJ�>����V�k�Q�g�U�묯X�m��}�p*���{2S���,g�`����V��赒J�Q��`Zn�oK����ƭA���H{�uy0�D�^�u�f�ZXҶr�u�yvI�e4��`7�߭ȼ��;�9�1��
T�����Q;qt��ǈ=X�}w=���8� �£�����q�b`K_����O��-*ŋ�����&��w�BP���	�͕)p�t*Ui�����i'"��P�_B.
!������BE��ٍ�B/_
w��`�C ��|�N
�B|�,�b����+p�+8_�BBo^�ǲs�o�<.?0��&�w�( ��g��]\h�����((�v���R�ހ�{L\����ϙ��E�-A����,��1�;����4����K����j��$a��8���
T�_�qj���@ֆd���y���S5k���/Ō�k�b�8�������`��o�g@/���AS����7�N{��u՜�a:{T��f������Ŋ�Qs-��m���/���a4�6����s�?J�R>5um����E`���'_�$9֡��m\�m��+��t�����?�Eސ��{(�F�`���it�j�z�b��k��ߪ`s��)�s���?��J(+��lk_L���Q��=�5�t۱.(����j����s���:Fv-�^����>��	��C��}�S�jjb�k2-]���v�K������"�c�>φݩh'C� �(LL�����3��مlq�@����� �Ή�n!ӭz�Rf�#�T����0�u����]��CӤZ����T.���G��E�=�C�7���gbָ��R�h��7:�8<^�-��?u`� 7�2l��pA�)�K@o�Ä�-��|��7�Hr�$o�9�w��׷��Ž��t���K�%쓖ʔ]&�6�n�.t���c���&�o����N�q�l7Mb���r�QT��?Di|��鈏w��/��⊪��a���6�xl���%���AY3(Ʉ+ˑ����*�|r�������&�b����o�9�u}��z�g��|g���|��V5�I�/���Җ��b�x�bd��!�r�Yb�5~<�~�[����J��W�v�ؙ)���q�Ɓ����O�aw��<rdO�b����M�SR-e������h.!�d�����OQ���7u�Ȩ$��P�q^�b{�+�B�W\�!�چ��M��x�0b��Ӳ��]�  ��װML|�5>8�����@�>�#��9�'��G
X�z=����m�D�=��|��n��������R���~ �Ɗ�N�>�W�զ���u@�R��b`]�d]��26	��Dt���4!9ﴡ���-�u���[͗0�a%�����8�T�M��R��T�|GC�ěG���æ���k�������(�D�1�@�y�j�.|��:z>�
�r�I��:�,�)X!��d��7a53��g2�d���Q�4љT��^%��ȚƱl�������m���iq���^�?��k�����o���,�n�:c�����Q�&�l��O;�}�^վh-Z"���7�P�^�/כB�з�޷���m�����V�h���	��%9{��9��}�Anb6�Y�/z�Ɩ#��Gu!Wgy�dcq�.��[�Ҽ�6Ux5���J��_��<���j��
�)掸��V+ �{~F�w��;)z.&���hb�@+Kz��v��qB���N�hD*MNR,p�Am�
����Э�ٺ} /s9�YI&>���c�(���~Q���>�4�k}�,�&|�%�ǭ$|���Z_I�䍢�÷��I�@3_�ڻ$p*Ń�D�k�2��U<��� �����+��FKQ�erw�le�>���jv`�F$�%�ll���� DV;����� i^�N�������ݤ�S}�z�7-�G�E�\�(;��1O)'V��ߎ(��bkKi�)6�[��>��j�o����g��[���3|��E��WE��ִ)z(�sM[�n �O�����Ǚ�� �Wet��ٴ�/�j\�3�}S3b�/�jꓫ�J�g֊e�'�eΨ�{5�`�! �+7��#^a**��C�Ma� K�� Y��
�7��W�[�T�;���I����Ui0�>7��x�JhG�O&8W<[Q�[(���{�1��^^5s��P!m��m7�A�2=t:�֝p��fxx���U��v4@a-(��y��=�Y�8�a${��쒲��)U/�[m4'�f����K�`���\�z6��Kbi�W�_˿���I���]�\!�	�� ���B`�]�3ы���kn�&��xT�
юY�ޣ�RuTRH�X'�J���{�b�~C���6�v����q��Y@%�6�WEy�*�������*��M�i57��d�|"���qx������z��G�3Ĥ��"��*�SzI]Z9��o�����w�$��ix��:\P�� ܜ6�ة��qB�B��Q�Kݲ0,�Q4�wN<�e���]�ێ�!DJ��r�A��O5R�#�G�P�:����#�T籢>b^o����e�Me2�(��J�}o-��h�H�(��u�7�Â��e&�Nx���}4x�O_�p�0���W'\�"�=���M�(���<����7䩌5�=n�0����|��h <.!'�c�������U��N�ż
�(����!���Ŷi�5͛�����<z��TYؗq4��_�̎�$���A�.��)~pH�:IR���@���W�v��K�'��^e�ggP��Y�GPp��^�����t�ő|�f�����`����ɤA�n1��Fg�*�c;eR��!�[NaOf�6&�c�i��~lt$q�D���_΀��r���eNF���2/#B�lK�,i���3�`�˒�P�}5�ʘ=-�jSk"]��Wɶ6��\׊��0]��vk��OO.i���=�!�G[���j�{�lǟ��X�t�gEW���㍀2D.*]w}'���C�/N�}�z���`
�M�B����]�TC���g��r�%_���1���%��٬<a��)d�B���3�'���@]�k �;�ʋ�©�M���rd
_J7+�b����n�is� c ���F����@o-����A���2=2��G�yq3�]m�]�=�Gc�e�V����[t8:��PY~	��!$��j�i��Y����*�>���A�;��4"���h�b���e5�0F�U�H��ѐ�_#��Dd"G��Ɛ� ��E)��	ï	/���d��ZZ����{Yf�WL˘D�Y�7c:�=D��}�P���M�ˏXB�/\XF,%觾�3H��>���D!+fIP;���i��J�c�9N�o~닒�t��7Ō;���7��&�  P|��\ur��$M�V�С�V��	���%�n��]Q���6�����̷��~� ���*��ֶ�T�c�-��O�oBE��.����1�WRg��h�Q\��E�E�9�i��`�R��-��L�-� �k�+4�"�b��������c"��e�b���%���M,S"�pu/Z�H�!���`>�3�!���x�6,DK5���"_?'����>@�w�����;���?��4W.]���Z-n�D��p����5QIY�_,b'K��<V��X7�s�<u �D0ᓝYtrĊݦv��07@��S,���E�Aٻ��+`�����������`��w����x�ި��Uep�ߋy��Q,ɦ�Zs�>T�������Ć��q�(a�j`73� ���Dʹ/+���y8��:��t�H��̥\c�"�5j�Ic�p���c���X����A�z/�UO���g_vþ��Z�$��v�U&�֟3����x�bƳjv����X��x�ܓ1ɫ
jwI��#u��J�z��(S��kw�:4Du�&����󪑋��|����dH�?A��{)�X�cѹ�xl]�$i���a�6K����46����9
���ޠ���,<\4>�T9�ǲ�����������.)��-���kM|+�L�Y� �J����������)��!�l(�ˀ��!UǼ��=9�F~��,���(۞��J;ς"vjX�P�m�Ru"��u (C�Q���o��l4���n����L�[@S�D&����W�X���Q��%2Ϲ�� �z�^��m��G���8�w	Qa�os־�+|��w?��ݸ�ä���`�ۨ�Z�����]QM[�$�	��C�E,���gI$;E��[�����6�"����vM��/�vREg?<Ϻ� ��s�+ ��\�F�'�Eّ��R�54���{�Z2�(��J:ϳ�;��ⵇ�=��c���p�oϑ;f���nyͩV����K��J�2;԰>��J��a��(���h��Fv�j$��'V1�D����$��j��.(����8Y<�q���S�ɱ�a]E��P�@Lس6�9�;���D����G�٢t�͔$��S��{�/(Ojk���eNI��u�Uv$�K��*%���v7�}F/,,�-�"��+Q(���z�����X��CĄs	�oE'b�)xeO�O�R������=Uõ��˹� �����P����5.$��74s%�Qcu�ޗG:��5e��4���p��b[��� BQy���쇣��Ė�Tˎ� ��OO}
t] ��kv�ΥK��F;c;���~.���Jr?P2�,>�PK�Y���u����J1�Z�������'y֊ٳJt:�Jj�TE 9oQ����I�:9�Kw��hG�A�Ԗ����2�ԛ+F�EM�5��խ=H�;��t]�!�>XoH�&�����Rt���M����)��VnvE����H[8�ޝ0l�*"�ڌo�	���yH-����p�:���j~_Id��6��֑o����:d�2q�#RE)Jĕ���%M#�ZV�L3�>�%m�q�c�I�"T$�no����m��J�ʟ�_���mv��A_��
�#����b��*�⨦�Wk{Ud����T��]�B�E&Z�k�kK��85������foSZyN�}�.�r��($�.5��$�`D�E�j��j#�v�I�!�?�\�::�3:�s.XZ"*E)��s���>�F��=Ż��t �b@[<���)���rQ�����3���A������E�*A���}���q�v����my�G6�)3ƙS���!���s��2�s>(Քt��-��@ۀ��C�)�j,��z4�RtN)�vZ�f�Y����*����Z���8>�0ы��Q��j-��v�.�g�������mQ����*���=2AA����\�$�,fr�!��Z�J�#R�SRZ>��\��󄰡6�5
�3�؉�l|�k�����щLz�C���֖pp����֓�:LdЪ 諈x=�`�̙kBnMڻ:��P@����A���2�v4	)��m��&���XE�?����u��GJr��j�����eT�Ռ�r�P/�B��<��++$�� ��Y5jd�y߬���/J��an�=�b��K�	O����.B|�_����#nO+����%k��_4����垥{T�%�[hƀ�(<A}]r�*���o�Yo�_$e��2��O�k�몸�Tݞ��?L-�%QL�M�z�r}�L���G.x��P˥��QN��˾��;y�xb�r���/
I�Mm��OM�<d]�#
�u�NiG9�Z�@ֻ�[^��dD59�{���~Hs�7�Kӝ�' �l�(J��I������}	u%8�c��B��
96��]MV%ߥ������7�Y��fֶh��J5Q�)9U��^à������Ϣ��l�^�'�����	���=8Q�szR�\����(�����I�;�И�X��tW�_��4Cm1Je����0ݾ,H����`Py3�f�YZy���� �H��~ɮ��w����^�=�#�iIxdX r�0���ǐkj�q_h�˛%��G������>�˨�q��jn?� n\-	�+�gM��*�=�C�U���j�WV-���%� 	���=�k�4�?�-v�P��)b7\!�n	ʃ�!�3f���>r�L.f�����L�fqa���B2MKo���إ�'���E!P��}�����#��W'	lN��}v�����WJP)�7j'�Hϲ�-w�H"��.!�k˦�Ŀ�Ca.^Bc`�3���3�Hv��Տk��qv��q���C�\�N�$G�E�pE���DN�x);�Ҹ��ײ����$���lj~��8*GǮ���N�qW�G�3����-�w���Q3���坁�D��rq=L���o��2)ce��)����$�!�n���!p+I��$k���lf���L�t�m�[��]�IBn`���y�>�I�%X�5Z��3�;e�i⪎-p����5|r�W^�?Re���n���l��s��!���,�@ho�D��#Nw��|��V/`N0����k*n��?��+S����U�f�0�ljr!�QP�Zw"�1<�0{Teu�5L ;ʦ�F:L�cWVr��TwspNB�q��D��ι�$�]^ ]�Ґ��
�O>��&xk̡��9k2�a$'Ϻ�9$�i�9�<\d���@@��Քإ�8@��Z@<�;���I;B��	zZ�$h��-�2��-��\�-ݞ>����J.k�_�JƼ��Һ�$��:+��0�pV�Yg��#��݁���?�4E��z��I)��	>�ִ��i�!�ĉ�6�6>�!7.@��F������*��$A۞���t�v�|�:I��E0���Lx@	�+�if�e�{x�ihϡ,)�vjM�� i�%E(��%�tv�w�r`
�d
����-�@;���M��� �RNJ_%`AF7��Z�$yHe�o�,��K ��0NДb�q۰���4鳒�U�諡���������B������@%���S�_��F�����[�D���s?���$J�� ��E[��uw��2���)��z��r�p6�U9J����t��ӏN���(�^�,/��E�?/�8��# H�(-�� �xI��	2�[�%��"/�K��`�Y\�쵸J��b������E����g��C�{u����32l����K�lTax�}.S�bt����W������/mӋJ�L��������Y��%����3$��#3��Ws=H�"��pWK<�{���q$�<��ࠈ�lh=꣌����y�L�;�Jk�7�<�:EŮ.�����$Zg���h�Z����*�dQ�66h��ˁ�^o�7�T�;�A]}9X�� D��4�{7����O}�Wֵ����/)�#0$���H2LD(��HT3N�E��[z��Ϻ�!� ^���p�D��w"��^:8r�+aU��I�̛�Σ�8�E�)�h�­k�@N�Jm*r�L�AH[�,0�e�'��G�Ǩ���tP��~�W%�&L�'_�Wu�(�[���> �M~jբ�T����1�~��	����V8�~Uy���(g�ǒ�t�
z�y����̀#�K��*ʣ/f�7��86��;;�c�;뢃��L
��:����Z~�M�(�
���A��_�|@�˓�6��P�����J���C��.t�Z|҇&�Ͷ��2TV�dE�
9(�&���\l�Hc����p�2�?�b����/�޿�EF��5�T%����і�b�}�|r��M�}k�\��C`'�k=��c�~#����г�,�ԝ��h�x �q$L�ʾ Ȕ1��̩nY��Z�g�ln'��9�Z��@l��JB�����%J���mi�l��ۥ��E�6WȚf-aK��G�a7�&R�E�EN�咙��'V���,���+"7�I{R�6�bZD�臿��1��i�a�\�-��}Kb�j�v)p ,!T��AOF��:�S�+��Ȧ�`�V�eFٷ� ���Yy���b�$�+�_���"^���I/gz��){��ݴ�}�d8�bh"62rG@%����N�(Pg�8�$	OCtH���
ޟ����iT����7�ˠ��`u�FV��޻=��Tp#56䇕�ּ2]�R�R�lm��jy���sx�FKQ7�o���K� {���I�0P9��ե[��V��H�!�[��?1��[C�ȕ��Ĩ���6?�gz��?]A9Nָ;��}�e��s6�l�r_��5�� ӹ�z@ĉf��������;ҼI-�	;���~;g����5��������Q�Z��LΔ�:]7��'�{g�}�� ԯ7�J�"cM�T�8��J'W�a���YS�j/�ce~'�Z�%���=҇����ݰ8$^���C�H�=�W����W��A���ȯi�=�ԫ1�*�����$�ҳ���<2@7*���0�OJ������j9����-�Z�f��� ���F�wM'�!�p�_^&�5�P^�-��.�g��е&�L༿���ƽ#6��U���E]�zJ<˳��[=�f���+/p�(uL��i+��8��c?P�MH6ѩ@�]P���rsR�k�	��q�o�PK��{:~��*����¨�H��ʉ�z���Z�m�f{���`�û���e�b���m�/����iu����MhBwĽ�y�[��湸=��-NQ��nn�nIֽ+��sm�M��/VZ}=��� ��ɀr���ΐ�{?��נ 7��o�έ:s��F�2���	i��wA�������N�i���e	3�:�ᦅKDăZ��ݚ���nq��9X�ᳲ����V��S�5�_�6�pU�`�%��Iw��3��~�#C�@�׎-%�q��u�x3a���Ͳ� ����3�겲@l�+��9��r_�5{h1/��LSl�If�J�����2�.�QLC԰��no�ퟶʃo�r�������4[�Ӹ.)&��/�夔tF@�PS*��*<d����y�~$]�Ԋ�<ُ&p�� ,{~C�s�1���4��q�G�S��<}�Ā��4q������˃���x䵴,��2����:�����ÅoA�Q;^��/h��W{�31��T1�o7� ���)��Ҹ�LG�p>�L8$�e��O�"Y�mi�Ω	����\�;�s�nG�%�{�t)�T26�����U�F�`�	#	�S�$�h�����s=��|!�_J����Y�l�өR[�6ͱÎ�w3�Nۿ zE��!���~�X>��)tʹ��-��|�ʔ-�f��p 2�\����=��&���d;�`��=�&OI��Jd߈=��p�Z`Vd��ε���#Y����՛�7��uS�1X��MD�+(J�1�]u��ﵺe�nN1-�@��DWHRV!SN���+��������������p���bMi5�� �vI��`d>M��Qd��2]1��d�vQ�A��PA� xUpp�(�hl�!k�x�+�� ��!�z����0L�/d�մ���k�bт-s�-�d#О��|�]��4m��K����`|�����Hr��V\��@%a����&��r��텆a��Y��V�K��}:� ���Թ����~"���ojJ�C�b��W��Ja��Afى{��@i����d�d��tL(��"�՘�L{�r��n��Ŀ�C�4
�Y�}ե��b���HzY�M^O�����I����A�S�qF%�񁎃�
�Z&B�M�w@ÈarT�>g��Kn���j<�̺�zQ��M�.��+�]�-�4�z=�шX��meygI�J[ #xu�E~d���A���s�Y�V:r��S >�x�M"�,�&'�h�����Ě�`�5){�-M��ǜ�a��ϵ�3Z�x+���Yb���^I(�E;�Y a�jQץ4�)\e�G�z��.<.���ɟ+�	a5<�T�/��U]9�J �$�ֱ@:����h@�&�{�� /�*�K�M�%7'&�ĿkLmt�ﾊ`�)I|���]��.��rxʮB��V��τ�@���!~%YP^��\����Mv��_�H�?B6_��)�bo��+8���c�fﴚ2��Q3琹�8��}��"�N{EM�eΞ� 0H߀x���'�hO��jK���S��q�S�i�F1�|������x���~+�ШYq�8���O%�G ��p�+C)�?���D��'�٢��u��Ӏ�?����(���&���5U�tic�;D�'���H�m��/^��)�؆�c��Y����N����q8w6��գQm3�8N� ;���|n�Ǡ��h�K"T�F��!����|��.4����j�x����U���!����[��]D��X~�e�|�^W<`����|O�ҺWF`&�kE,h�\cW6i�pt�2����`�M��a�g�JG��dx�^�&	�D]
�QF��1�S�e��)��[Y�W��g�>�$ڗf�p�lS��V����]�L7��&v����{G'���m�co�(@.=3kYD��R��],� ����o��O7#��>��-�+��g���68h�f�c`�D�Yv^�� �����c S�0����ξ���I㹉���?�D�,.��|Y���n�xѸ�M>��w�;V7�.����"`4e ۤ�JP�m�L�bkh�/]�3};�~��I�</��,����߮)���WX���<��e�lmed�DU��!����!�A,��wo^���y��5;8�*����fv�����cq����/^�ı�����ը	=`�~
���xF�wlmiI�yX끸��S�$7t��Vb�3;�ܷ�r�&I>;�5/wI Є�'8 @�)#�xP�ۙ߄,0^����u>�u�/�mh]wJ���,J�f��u=�S�tb؇��T����[:����)?�ɓ������vpm���J�TcB�D�"�j`P&&[2<I�FK���F��~L��g�@��&\���Y���o�u�z=YL���,����ES+0[��;#i0�\ȹ��9($�V//��%�}mgE���8���f� ��������<�1�\����;���kc���X�0؂J{:z�7���&��u=̦H���#����M��8���O�"n�~(p-f���"uz7N���K��,�k"kE�&�����l�2P�R���lO)��O�񙐣n�»�{b��o���k3����&�p��B�ݖq�������!�UH�I�tݳ�����ۻ�����������G�E)���m���5�o����p���
|��Q�=;$��4����ͬ�� ��vˍ$m�I��de2s.�Z�^��y�z�h\�UMG��!����7G`�+_qt��(�`b>�B���7^�`�&�_�VG��:�����`!�\UOM�SMj��}���$����!�}���c������ �8����+Y��D���e���k�M�sq�ND,ۊ9�8ưI��y��#C���m�i����=c|��˼bj} Js#����՞C}��T�RL����K�?+F�����7p��B��9�@ Wt�.�v�H����%.�����oKQ�+@��QB�c��t%;��]�֗;f!^�#���!�>�^p����ԣ�B;�'oՀ�T
T;�]��R�,��˅��c�5/��ɟQ����*p��՛�j?���'�����6�Rl��q�U�Q�Re�V��Y4t����?7�� z��巍�����f���%/��c#}\�{��4����r�����t��tW�Vb+e�L�@�i�Ž8,|�4M���
�"
���^Ac�Ʀ��3�j�Vv�U�Q��vl����LA&4���iwI�9��YcEΒqj:X0C@�=M�X^_�z��̔�3��
O����6AZ/��2;�N!.ٯ/7n�/д[OZ��󸕞r%p�THu��f��J�-/a�D���Z�-�WB0����y�b����?b������N��a�p�
�c����Ύ{��Xr]B"�����ղ2EPHD�S��qqsc{���~\�{����'��LP��Hx����@�KS�?�|�������&�9�Ȯqu}Ͷ4�f�����>yQ	D�XWf���r�ؙ�e��Tו6j8y��=�n�S���i��I(�͜zL[���ێ�G;�N���&W+������� x��``�Vh���܇65��ַ-�{��ԸE���b�B�Z��C��ܓ0��%y �>�M�a�E�`�z9��4��p��h��AbP&x���'�.�i)Ge�Qtf��'�<~ ngFʛ������ b5֑���1��[%�t~	�o�7]�3�������>qFǸ՜���jb���y�!Lu	Lq4����g��������-��ati�!�����	;X6L����n��Ij�3kQ���!bP�ʌp,y<�����K홏��j꺲�>�z�uF3��~S�MW�!�f;��<�wN�%��Ҏ�h�k��]�^Px�^�=�"ޚd�.�H�hAʖa����sLt�d�K��<�w�c"iHrK��K�q�Oޞ�5�pw����&���s�c�}��帳�8�/�Zm�kCw�����$�����v��(�E���n��t���'�*k�
���#0���i�AM�êx+����Ⱥ4t�ߵ�F����H���yU�]�o�G�pJ�\�I8�ŵ@.��r�:C�"`$�o�6�ҕ�K��G&5���u
�Ud������j�:
l�M���MF���5*ҡ����f�w��t��h�'^H�H%� ����k�v���0ۍ�M��W]:��aR����9�S��Hƽ�����D��)��.�ۃ�,�xK��J\Y�-��5���cG�}��⼪>NYZ��v\ޖ_k`>�l��岍�����$N�KL��!�u^������\6���t�y 8��)��� '�@d��v�������.��0���@����p�$��s9�~�T+P��?�\	�09o���y�6L]Yq����dE�#����w����R�Ϧ�x�_�LӶ�m�Hi�w�L^��Я�P������|ݻP6qD+J��8$��2_�5����Ӻ��6p�EH��T�<�ȹ_�'�R�JR�� �m�%�.�e��j��h]P����oWNf��s��\x����p�� ��=
�'�a,�P�⩸��Sh >��[j�g6vV���n��d}랟��Cs	H�� ��O"Л'�'S��#Fb@��U����<�ƮH��KK Qz��`�Z1���^~z��	XDy�?N��{i��)-vE#p��߰��}j��q�F�^J�l|4���j�s��澜�����|aX��W T�QN{�8E3���2�{ɒ`�$�K��n�@�V!����̿Y�H�!ǻ�H{��j��@�߈����8q�ZBRz	���V�d��|n��ijǍ��{�o���ܷ���$�����#>�Ml���ν�t8�,_�(��o�*G�o���虌��kB�)� �
�i���^�)Y�ף\�6���CG
&5P9��`�BT莾U%ؖ������~i��Td�O��� �LY���%�!%(�pѺH� �;QVi� ?��ا��y�ě��=��#�z-�����8�F����d�J��a�gI��'�z K�VY�#�`�~�9Z� �Y�q�e���z��lV]d1������m�t�c?��H�0�[�؞���