��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`����.vr��nw�%�{�� ��}D��x��0���<999�X��'JV���p�Q�1U��̈́i��zB��x��4�p��GC�cd�H�)��s��Ģ͍�mB��@|Y/U8��4b��͢��%���#�a�$�Ry��� "�]}Q�������������4����?��_�(f_�|lh5��J���!�R�;]U�(9���p�A/�эrfzU!Ԧ����sV
��FK���}}��d%_�h���������.B��.)�>��b)�&�Hޛ��[sș��(�i	w�y�n�K����xB]��v�B���QB��IHl���2�V<�k�b7��P2��l�k)�z�������f��:HR杮�`��<����`㬐������-N����Uy�>gGs"�\m��g��<B���]�WP����eݐi�_v`������p'Ɵy��?;)�$ʡ���5�� �Ce�ڎ�Kz|�_'����Yb�Ӥ~�[��D��n�����y�+�6P�U��3'�z��ŝ2tg�`1�U=���mL�����S�[$m��E�CH �$���J2#��3'FS���=�;|����
�� ��,����
�N��]�[<�G[[���a-�p"J=��V��M��)�o�"Rz3��\��r\���J,&��fE+����f?�;��f	��^A&���b!��%�{ �r-�{`�5����T��|w��s�������ٖy��1{��<��?Ηxrg���NigZ=��VGA2W�=[��R�*O��C��}i�$��,�&�$N�L��U�K-�0Q�Hb�\+��m����m�[���uoq�$.i���Y�˩�)�^�lZU��I %���
�+�K�C�������F�[o�z�Aa�6���;'��W����!_�r3��,؎�)=y'��	�9���NK���)�s���l�?N���|��Ix@��._ф��f����Lf�#�,ӗ���)�2\�t4&�J5)}����H̭����Ǡ�*�pߕ=�*����C��	�p�hfE�Rd+����ӌy�&�6�)w`���$�2��n��Y���g��tä�wP�yQ�ڴ��Kp\�ȃ=H�ƞ�7���E�j�b��q,�������>S,ɢ���F
�覸ɃϖRN�`9�����)ᵚ�)AN�C���;��ھ 3���*D���kwJ�*fD���l9�L�/�����I6�����`zԯ�S�^����
~�b��<˨EXH��-����邎�`��t�s*�k(�!�[�Euv�t�8e����PgmG��m{���	�G���A
/�R��^�/YgW_2[�UUpc=/a�)�E5�M� �7��Q�-���s�<����e��s?A­�%[�w��¬��D��-ص�\�ޤ�Q)A~Rg�j\2(A�]#�]�����(�k	�j�G�J:��0���>�y��*vJ9.vO����4\��қ/x�ϖ��r�*�T��BK��SG��'���2u($k
������l5��r�Ƿ���7C�@���S`f��5�'U�D��� |���,���pے�7���_��R'Tԋ:^�O�U�Ɉ���/��1Ԏ��C(�Iߝ��}~o��������R��K��|5y1?bXp�"�<G[ʀv@\�]A��<3�\{��2aL���U��k�D�[w�;
��%C2g�����؏QR�t�l F%/�%e��	l�^��Mw�+���(�~З@�]Ao�H���:�BB�_����Y9��*��U�I�e˷��@'U��b�,)s�q#| /A�n�Q͒�"��-&���	0��	R�'L�n�e�( �S��BL�P��#�$�TTUՐ�{hj�~q�>��{�ʷ�NC��S���O��j���=�nH�C�j׮ke^�� ,��A�H��g8���K�8�ޏ��Z #-�xA��ux����eV��n,m�O3*��[��~��ۜ�������b8�%M޹�<�\�a&L��͖��$��;P�t��#g�$�ll;�O��j����:[��9�-�1$�Rd}z��"t:�B��19���O���.��(ǚ�d���?��&v����GS��r�k�d�	�z�7/���1�E^`r����i���	(KGy��g';W|Ex�N�