��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�q���4]oHe��zL!�[fY���f~�2�����z�S���Y3��1��";�Z��xp�����T�<k�x��UEX�T,�ߪ�+h��M7�87d/S:P�O#�7��� �A������`H��EzC�r"�������Z�e�����e�6�K~H��70l�k�-L#�Ea��Q�JIJN���1�u�0��?W���]T�W`K}RR�����̮x=��TN��P���q�o��WM�	�����������j�;E8���r�)��yKa�'�,��4.1C��{�OV���a�_3	qvߠU�2.hz��t�o�S���r��������G�ZZ�2���H
�
�,�{���Bs�iRY���8S���5;��<<�o�S���������u���_�
�;�y�Y�p�m�3ס�|��8(�%��_��VX���:��P���ņ�ڴ)K�1FV�j��T�Vy7��PZ'�{@.�K��/��fr��j�r�3���;�F/Y����T5�@��H��
���W~��s�z���~����V�Z��BĞ�ӏj�X�X�Rbv��*4���c\&j������x��,��O���>���
���ͦ(0R�(iy{�����a�;d�O"�]jq�	E��^���z�>�	"W⊦�\z���2a2U�����l�X���A�4� g:�2�^Y���m6(���3�d}B�W������ϗ�5'�8]D�c�Ј]R�W����O�q���]gL�U��1b�����m Hd!�"X0E���#�	^�H�����b SB�gO(���������K�u~�ʩ�gF��V��Դ��j�n��X�Y�H�U��]���]iNE
�������_���!�w��8�����H�sߋ���Cn1c�2o$������R�3X����P���*a&���E�����b�����7�p�;���+ �{��c-��.�Xf��c<����IJ��l�V��4`g�y�]�U�$'9�xK�Z��f�+�6�v�����z*�Q�'�o`CY~������L_E�d��G鏴a���Y���C1��&�T����grN��0A�t�0�B^ʽ��$%;2R���w�:�$�&5Z�"�	��#�ܼ W>�+fJ�	�uS:����v��)}`�Cj�x-��J]��+C��2Q,IO���w>9v�y���{)�`�̡ɚ� ty���������X��uڣP\]��tG�*�k#����v�����U�<�����'5!����[=��xh�M"h���#/�C�b7!�D!�`�yR�{=k��;&L�mJ�/A#TΕ�`m��&��s��4ud5�DG"� ߱�G���GMDC7pMBo>�ҌͩۇsU��D�����K^O.�oK]���̶oZ���Ay!�7�Þ2�6�T�X����M-C���8�&TC��=f^$骿7�ަB4�`���/��
3�\0�N�����܇d�����q��u��=��Å������+7JHL��b�!>Y0c
q:<S���8���}����w�B�9&B�\�R�v|�VQ��	"%]nH����sCO��pq�8-��$��·��)�N�L��¢湡!�������zv���џ�ǘA�,�	�/c5n�]���xR�WJ�+����0������͉O�-뉺x�[������(� �A�H�]���h����[�"�[�V �u����o\ӁK~t"j��a��h�J�:=��+!���R�I�d����d.���kQ0�/�aH$�����x:	/ܛ_��m�[R�CUV�8�&�[t�In|���j����H��N��^R���v����b�^�[g����z<�C�����~9ۙ������Ψ�ګ~�Ľ��ҏB��j�O��P��F���:x�����X�>U�V�I�ڞ'���¤����GS��1U���c��y�s���4�)	
��-K��Y@���3�S�>e׽���GR;�vP���C��=�B��.�U/HI����(-z;�^�����JȔ�>{� _~��E�^K3!��;�g�ǆ>�0���J@Z�A�Ia��\�G� r( .�;��N�D���k��E8pN"�SӜs�t_[���^��w�b�z�B��8�.��xK�NhS���Q�NmX;f���7�Ͼ�Pj�/]�S%J��-�F�՞�1�΀v|�dI| ���#I�����;�K{Btjm��_Y���X���dQ)�1�#�E+X�R�f�ɟ�7�iE�k��-ݜ6'ՐfBz�qy�2A�0ߍn&�Zy
Qy2L�RWypfl4L���#�X�6dD9FgxW5j����=�W��>B�Nv����?���-�O��n7AC����̣��L	��H8�>���{�h���AM�v��[�a��̕V��e�57P �X��sdC�p�x$��V��:+~��W�β�].S��B_���V^Q���f7��J�c�������39�b2'&|�s�VC����VrW�Nx�d�����3��{����R��=&�So@��� ���]�Vj�E�Wv��,x�V/��e��${o����˜芞�}X�u��	�~�r��dL'�-ΨR^�i��h��*������2_G$ɲGl�������O��y�p��+�9�MR,�QҒ�il�ĥ����J������b�3�da�4��3Tm�+Gg �BO� JA3�RslھZs�9Xm����"�B���=)��l�� Yz2�q��-z��f�O~����v�[G��Ue	,��z|~8$����`)"@�MV�͗6�J�9�lg@(���]\@�����MD�1S��8u��S'���/�s}gzl��-�ɻ�i�Ӻ�_r��_�~&w��~�}�b֋�|�Kvj�KH����9MqG�󎢂���;H��c�y��\�W��.���."�{j��Y�K��U7�*�g�O��N�-�@�Q#Ȗ�1�"����7����;w�+.7C�xL	%��t�K4]lZ�ѐCr���o�@~����[6Q�\u@��'�	s�#����;�ꋏ���f��٠Id�3+]�G����vi�AF�6�����Q���0�;��"#PD��)1��snr���A�8^�+ʠ�l�A�ţ�� �z4n�YOw�6��s�=u&3I�:�]	V��T�!����^�N�Ld,��W��Ti !܎�{���QX�;��6[F�q���|!��͊@V;������A#n�L`IOiE�w	ӝ�ܩ�@�����������^��K ߗ]�X c��~�'I�=���X��
w�Eѭ�wX�"���{�g-�q�@l�[q��	���?-2%��E �\Δ���Z�S`a�l�_M�vm������Z8"#�ǡ?$R�d��2�xl[ؐ�a[ae(��\6�}J !�K��]r.!��TW�>��{�0"���u�  zzd�at«2��P��4V�ƣ������tq�Q>�<���b��?��}+�����<}1�3G5\����n�]洣�7�Lbexx�oa�ʍ��9&��|)��6���m���h���U�C�4��:�c��P�2� M^�j~�[�Iha�����y�GcN��k.��y�Һ�	>��=���Mw�s���J�"c� �Ly8��ĻU��V�;������ɫbE�[8VU@�`Z=���п�� W��5��84M���jk�D�X?#L��>��>x�H�A��)[)a�*F�	�];o�np����j?p�Y;���ȗF�a��4O�6Fϵ�V��=#]��^GA�E��0��y>��t���f�� ���ki�Mՙ(����V\����-2O!��*i��?o�������*���`��a�y<��%^���+�hё�^��sܹT?U����v)6��2b$:>�]$���73}�qL�k�zzͩ'��N*����Sq�vV�⿼M�^�Oo>O�|�+k��S���Q����pj��,aH���Nϔ��ة�
��L�K/���TK�d���X����-�X�	A�K��8������80(�o��ɶ������V��7Y��'�b�Y����knv���p8�D�*��/N������"�{A �Ĺ�쯷��l���Rh��=�[2�;4S9#i1�v^VM:3�\ڮ�y�f�^G�Tqi�EJ���甞t�
(���R�=;�~��t۾h\��2W���J����%���.�(��Bm-�{+<������O���W&NAf�?���~1�d�Τ�
�7�7���P���ͮ���j�[��T��>�Á\��)!�L,�a��t)�]�T���y�TN+�&�=Њ��$)z�]���-�ߺ�e��T "r�-�冪���3�_��+��Z�!? ~���RF��F��p0�y����%vᨆ?+�\r��c�*���L�f��j_�7	�R���჊o�m��ޥ`���"-&J�9�]��.�]���0�_��X��y � eh/��X�j��e�W��N�����ݥfݿ�.ߞ�y�L���L��l�\�N9��I�O��d�wr��>z�߉xM.͒�L$L���nGٮ=��"A3;z����im�H d4����l�*7�.f��׷Ih�p�b��2�<S=�LԥQ�
kS]�a"t/��$
����!(�+tj�b?����GC$�[{�Z�k�[�k��e��9���Cޣj��2�A�D1��ٚ�,7�%���Ą����t4���fS�by����)mΨ�5h��#t����퇏���]��?��`q�c��d�=TT��R�E�[���m���Q2ꐚ�|����l�������H-*����\�X^)�pz�D׉����()TB�"�7�W*�c��fwSS0]+�Έ��B��v���蓠qb[G��V���W�ʥ&�{*pir�?{�9�=<�3������i�M��>2xD�Kb6���	o�� ��Wt��Q��`�*&���'<����R���}�p��m[�P,愽�"�V"���_S��ѡD����)����i��L�E����J]zh���.��W�U��w�G�����V���4.�W}�I��J?�̶�.V�$kx �m8�u4�iwӟ��Xۍ��};UͲB�$�*wZ���Pg���WY�7����*�E��ɸk���	�D�j����>�GS��9��ᆏs�O�\"H؇,��q�L ��ڦ���޺W��`�T��՛d��l�{���gӵr1 ����I(�A���>z"}ciMk1��Xv,6���9�i� ���v��X�ԛ��t���vYC5�?}���Q�{����_�@p���.��jz������p�����&y�����7�����J2%����W�̯~�S�gB�/�s9��	�����$נּI�bn��Q������E�[z��߿^k7TQ(��	Yc-�e�* h�q/4Q%���-L�h��jtlM6�ΠA`��eC�(I�;x~�v�dc��cܨ��4&N�^U8-9�m�p:�g͟%�p�N �r�p�D�['��������",	��� o�l9eO���h�p��Y�5�\�i�Wc���z�Ey!�LȆW�E_^#�'ĵ�V�H*��Rl�Udff�M�Ö���3)�(�ң�G�aa�{�{�m3��W�*�w@��D�8�R��t\�ݷ �[�@�>�r���ϐ�#c8�]�M��)�8�%�R�� y6�A���Y���K�8_0ǻō>jĥ��;8��x6.�}	�-*DK��U3�ͺ�@� ��1h�s,��!�N��򔞭nF��=T��<�J��m�T0�AO��K.�E����Yq|B&��4�iL�܋����gd����7��q/)�;������.�Бa�-�z���yh�����6����,��{�1iQӇ��-�p�o�[�7��?��|��i(��
����\I$��|ď�<-R��$>�j2P��:��ث6�F+yy��8��pk��C#~�캆�-�w�hӨ���؝���w� �<�bW�<~G�"��nS܊����"���5Io�����+��w�+�0����VI�p���;�v]Co��A�dC�#_�j��@9�"�v�[�V����~�� �4�8�p��iJ˕*?'�(D�O�#_���o�a�f�I���OpG��e�ef���ظs��]����H����j�	��_1�V�W� ��Q�����?�Ci�/a��F%��x^�ǣ��\(�Z�c�eW�7�}�j��)���TP�e�3���GЩ*�🡇���@z�� C�w�e�*�
�
0���F�qTY*r3݋Z��ZLx}�ޱϦ��0��p�\<M�	
�I6j��Kǳ���.M?3t^����B;�՞�)�m��uz���A>�F��dH9�0�����֚րMx@��Xgm:L/����}���5Jt:�b�6Cq�6��C��;��+Y� �{�v]I�N��t��d2� :7"ˣ�^�Cg_��f�Q�b���p8|v.�݃,�y�ɐ�,��p4��Cm$�$�֝�'v4�γk<B�ND. ϟ��_@8>��I�a���jey+��o�����\'PZ�"����
���}�����bn��Aٽ����Jv�`K�ܠ)��v�i=��]�^Q�^:�%w����Hq9���~Loi|�~�_�;#'�����oF*ϖ�������|��j!?�S��C�)���G쪥�t>���5g�= C�^�m��0��!�AjC4�����m�|tEٜe�3'�+ex��c��P2ڨ����ȁ>4�&%2���<^��A����H���\2I�	���j�6V��u���A9���p�U�!d�TvdA���j,\��F2��YI�j´�^ݿՒCT��r�@oR=�X��*3³�����M�G�3�n�\:��)�������h)6�� ��M�1t.o���]�R��R����)��2��,��z���nze��_:?Hi{����U��'�C�"��S�[wS~���5�ug7y���6T�iU)t�+�yLI@+`3N��YaV��x��'����?�Z=W5���dT�!}�-fpob������L�ߋ���B��:��<��`4�4s�~~���g�Q����8%2#vO�E8����LC'�,'Oo_���ޅQ<����{�Զ��]�	^ �:b.���T�kN�z�ɤ��;i���eTu�7"�־*�EI�>������l��kn3n���])���������p�C|�hV���a�K�hޭl��n^EMJ�*9�e�)�X(�Ӽ&��{�贃F�/CA��}D�+�#&u��b�*1zfK�k-�h�arTٽ��+�7��c�, �Ʉ>F��L�㰷E���3GM]�Q�`S�Œ�G3�����E�q3HsW/r��{� o����!�������K>��d� �/��7ٮ@>�kM�l�!��"·J�SEз`�С/EpN�.ǒɓr	~���]�0�{i�~�������l�Q(�n��Ն���Qa�q!T��%꧋:���4t��2�#J�X�/�C^�{��k�9l[���-D�y�18 %Na�	����ζ���Ό|��6m��/���V|b�iU� K �BU������쳲��0��{�~ϣ�j�r��G���<ZF��VPfNP��.Dn���6�|�r�Sd4�3�s� ��Rr,�0:�w��q֤m�)uxl���(nC��kP����L����Ã�|�ra�0�����T?����XW�h�d29����
���
Sb�0�2��	~�H�%x����j�dC&�zSf��;j����37u44C�mTĈL��r�~p߳;��$�K^�� y
��r��v.�_5�W�Oq��YI��kxI�k:���ހG��"�	�/|��ۃa��v��]K��(��KaX���݁(o��pǽ���e�p��oG�_=�#�7�2f��⹤#/�-|�1�~�MƬG�r_ϻ!���k��	c2K���[�
����uQ�t��:o�ꭄ��o&ۙ��h�{����!��8�'������F9��ic+<�m���YJu_��tU�@�E�����v�o�7X��V8'_��ܤ��Z�_	��Ӊ�0(��([��q����Ys���`z�iwJ���z3�iwD��9$y�mT!}N���ޞ7^��<bbW�����M&�*�45-���N5��v��0��nSD�+����BQ'�s�&�4�I~�{�^��e��ь^���1�W�i����q���]�$p��#1�S�F�#
�� �]���F�P?u�h�ma9 �ć"Vs3ta�4�kR���R��� �N%�;��q���zV`<�TEڈ0{�7���Z�<�#w�F��h����dG�I����S��:��+qe�,6��ۑ)���->TYs��U��+��f${Ȟ���Y��5�Py��8>�/��>r�B��R�v&v���b��%]c�sR�d����ߘ�������g>�%���	8k�e������UC�#�OD_��a:(�rS\U:h��iM�)���F���lOF���G>�����j�u\��\ ���~��A�� 	��;tf��� 'W�U�h�[!NŲ����e��!�J�ZD���%PB�^6,"1JQ8�����9��~�O[�#dh���s@�;���$k�\\�` �j�;xE�ƊODr�@!5�bO��~wH�Ax�Y�
G�2�8���K�X:!ZE�,+��I�\��JRK�8K����lq�J)��%%�3g�Cجp���Ar�p~`�)�����r�^(-�Y?m��V�K�-��I��QC�����\�>��<��\;�ڳ!a5=,-8o$,�"�	�e����ϙI>��4蜔��:+�G C	��J�C�k�H��SYm`,@iÕ,�cO�hi��-�A���a���0A���)��꺎M,�)[�+�^��su�Ԗ:ߍp4;���Y�䶠�Y��O@8��>'�G0{oOńn����,M�^����%��k��ʥ�*�O��q�i+�0����ˀ�[�JZpVZ��$��a�ouRMK��MkF��	�M79�r34C���Iv߯���H4���Dc�t�⠌�܂\R�-;��f\̩�@�P{�Y�������p5��t*�@�v!�ZU�}Ī�u�bT�n���9���/Qw6�3��Q�8�db� ��'�W���^n�iƖ�k��5��:��F�I��/���5��x�vY|�C>eh)��$JX������qr�����#M��W��[r�Z-G���`߹M��n}�Kn骚���ӽ�{��0������8��|t��,&��4�}A������?�]]PN���<���*Y-�s��|8�X�/���KƮ+8�&���O`�}��$��[�w4W�<J�o� ov��  �D�����Օwɘ�B�||�y��)�c~-�}ĵx����Mよd_�|R*�x��fH��C�	O
`��~�aiQ^(�bnt!�ؘ����L��
>�����ƒ��w1v� ������-�����~�I##��]*y���������?FEf��D��=O`63�����s}/C��iTa9������>�#X�����$%��J��蒿~�ќ�H��%ġrND��8^3L?���������G�s)~��E29G83��	DZ5��M����G&�HL����04f�?�	BHe�þ����C�t���S��uw�e��>��
�;;��	1��N$~�`�����k�ʼï3|���Cx:�5��U�+�VÉ񡛭���V��'�\���ֺ�����K��2��F���=Ē��-��� T�Ҁ�����-���S=a�]�4.^R*���
�VN�
�����Z"�����j�p�a��I�LĒ2�,���%jN�4D�U�Oa��#���*�etG�!<f��$�!`t9NyQ��ӖO$�׉���\�i�
�qC�����yG�}0��y�>�W�Qt>���#�[���f���s!�ݙ�R�C�7d�������?�
����ap9�R��T��9P��:s%m��K�d���/�6���Dz��e6mqDu�)��J������̟�J u�����s ���o���Zk��{W��ALч�ZV��i�\�e.���Ѹ��>-2�]6_Êa�)�Ah�����ؖw�IQP�֑��)"�����=��bڊ|`�qL�b6�m{]n��#n����&LP�4���/+=\L^`eCsYB����"'�f�Z��)J����~�a^�\��D��x�6B�e��\�Z\�do�l�@�
��U(��@��t� ���A87������ �>xe�_c.1S�}XHɬ'�nn�	���A��_�F���ӊ<r?[��({���X����Y�L�V$p.
ʼ���觚K7�*��Z�ҟ/7+x�l0���W!���Hh��Us���~��ʑm��3㍾���7��c�Ed�B�� t���m��ST��ﳺag�HΧ���"=އb{Y'W�Qj������=%Uk�$��ՏA[��B'��@1'<Lz����V�ΜR�_Հ���1�+mdz��hQ<]:z�����r�(�X������=��H����@��^��©?�)|���iX�B���FD�8H�T�h.v۱#�,I}k ��X��0Ħe�[=E�}#���fLr�����1���'�����BSF���Yj8��D�%�+:�� ZBr�YΣ�-��2�=��+ڜ��PC���=ڛ|+hp���&�q\G�ܢ��q�E;��� b7��|a�_$�^�݅v�~��c�|�"<��
1�<���LyW40��"���MX�Eo�$�q�T'R� '8�]�#����5�����æ�2�;9o�af�_@5����.�� �aeC;,��1���/�C�we��ʉ�W�boc�1���g%k�`�d�'�Z�u7p��[Ɓ�]�P7_� �,�S$�O.���x<��� ��/]F��틏[�� ɕ|�ZKTZ���f�é{��ٺ,a���k>`㱀�@�>,;��q{!  Zr�6�f�rQ� ������ ��N.�qO~���V����D�EF�C��:�o�N:z���8b��m^�e[�_@��E��	��"��2�����(Ǎԇ���z��{��?!%k>Oiu/�K����N;�mI�'8A���i�
*}�	nI���f38��ll\Z؏7![V#���m8����7B!��1��P@n��KTa���%�r�D�w1�H��4Ʋ�Ee��D�*cޑ��&����e�qfX��J�gY�-�ַh,	�K��a�'�x?����"Y+*�� ���u)�so�m�m��0�����`�:O�|W�媨�AP��|�%'�7:�7�A;��*l�ih�y���ܖGq��)�s��P�]��������3鷷���ҙ)�5;
TƷ,p��k���3��p��an�\WS��=e���;ߙ���Y��]�>9Ȕ =,+������>���s遉��nq#E�ma$�f��\Oh�M ��䉐�n�wY�-$�b�ov�����C�?���Y��f| q��{`#��}`��'����E��m���d|nPlg5j��P�NS�S>��"Qό�R�e���\eɿRR��8ų�D9��1]i~��E�P���'�!��E\�/rvء�]2X�D�S��=z�����rN�ub�K��=ƳN���y�|�Đ­�
�{�o�KG#B�tDf���#p�1����@�Q�臨Ά_�m��$��=�IV�5q���:�^k �n�����!�Ǟ�fr�08_�xq+�;�ʃ�Q��s��S�wL�JV���A6a����m�N�������`���=�����?f�֊�`�ts�~蓆��Ͳ˶0ݛ�{�'��|�`�5����)M|v����0� 1b�mA;�	I�\�N��(�ۋZ�C��ipl�)�/�XV���]mK�O9`���}k���j�oS����lr���.��:�Wa��L�q��Q}4�*$g���SD��9�tt�f���6�����6�P��u-F��y��7�����v�(�ul�Nt�c��|��DT�W6�8���`������yпP	��ĩ|�d��X� Z{YAhiܞ1t�f��D*��g"I���y Y��-D�*��!M�o��V��0oa��@-J���]9��DT �,��ߣ���xy�㍘�� >��q�Q\�ɕ��!�t�d�PJ�g�O�:����>����2g(U���	��(�Opu���C7OW�.�������i��Q�Z��+&]���V�3�mF�4Z��p0#ϋ��QI?��֭E_��×Sdv�-��;C���5��1ǵ�V\N�_WK�1qإ�C���� �����]��ȫ�G�\"h��f_��d�;2��grI�IF���XP���	<"��֥~߁��X`�_�Ogd�f�H�'�P��//�WVj�����rw�����pp��J��le>��[=<�𾂱|�B�|�|f;�)�p�6S�ZWg�A:�p���s�}�T�U撁����-̮������@�����~�uN6<�8Ot%��V����J��Ó�<�R�߿Y�t�g�L�<o"����}g�y�Z�|��n���1Ǐxp��oX�J'X�H���j)���7:�C+����rb���z4:´�t�Zg�3��hYڿ��C\�|�\����f������)��A�@r��u`���~����oq]˛϶8h�7�9.�g�Jf�2f;V����#o]�"I�RsF����1�|E�0��!j������"K;G� U ��k]�{�f��ǰ!���V�a)t��0��D�S)�VW�_'y&N�8�1��kp�Qx��]ߦ2t?O�v���5-=�>�ہ��Gv�tQ�G��ZW0��L| We<6��J&51Elh�YĘ�4(L����V��6}��}�Y��^ !��. �	ElP�O;t�zg@�ں�iz삱�ZN� ���[�b����61����@�Gc�pev�^yf$��\]w���ډ+[�"�q�D�ٟجb���}0�϶�����;� �?��
>�h��{���0G�M0���:��B� �ڨ	���Ԍs�:'���O9���w �D�	�j���cT*Z�J��Si��ݭu��om�s�z�	��ܓčJD)�1B[����0�&����`�/�INU*)���r�����wZ�� �H�1|�&���{��i��g`"@Q� ]ؑ=Wh�QˌGy*�,�?�4�w�ڭ�e�q)��>%�s�����P-�Ma.5��[��W|<l�E�>�
�4�ߎ
.��hy��Φ��9�J-���ĨA�j�	�0a���؏�޻�ׯW�L�Y�Gw�'1��v�͠
X�|����a&��+Ο��[�0v�3�+RU2ëoʅ)�:�~�\9߃-�&�����"����U��tؕ:��8���|R�P�I�Bk�,��`�a^4����H���')L��.�����E�%����B��)�Aq���
6=/�bn:�f%� KH� �!�6�m�L�Au��-�U�u�BpЙ�����6ϭ3��tIj(R�[;��@%�Y�`��K%?��,S}Sf��8���+�))�){�6q3�i������&�ݛ�����N�ܿ��W�>Nj7�m�.�
�4���~66�8/9�gM�ɬ�^�X��Щx���Tq�w�ܹXe�
�a
��������f��e�8J0�ߖ����)������������ՏH/͹����%�6#7�W$7�
*��?J�ñ�@����k�@��:!ĻK6���=���۴���.�4I�rBe.�J��	M��&O@k�F� rRw��
�Q��rT����ZO�V�%��z}��L[���Ӫd�W�m���9|�RaS�4�㱉��mo�T�f.B �O���Ka"�F���G�t�u��p�l�s��s�&I�jhV#��0���!�+vU�D(8r�,7|��#�N�Z�4�w�����<���_[o���yv�8;�BcSf�*��9
?h< �R�0���wQoL��'�_�h�A YYl�|�'����%���e ���F/��e�7���6���H�� �+ho�u꺝�@��E�dj*�=mI�(�^�E[�%1�������a8���a]�22��L7^�u'�;��\�~���U��,?3�����~s�P~�F�D�����6PHL��� �+~�Js���_����EaG���_�o�\a��̻�P�dg��Q1馑0��e�Au��%�$�f��b)��p&�j/�\~`���һ�k�K]���c���Ѡ��d���u94{�f�8m�.H��h��IR?�Z:lÜW�I+M��e�!>E���q~O�e���!�ia���@�v�ｚC��ɴ�@_t�He���4��(j�E>��{������E����Y���R���E�֬ZD��UN���P��H8.��� ��#�`dK��6sv��C4oܯ���G
��(N��e޿�5�~��(@]�t�[O�� ��r9�!֔J�����5���㘸��
P(RL�L�y��;\��i���㼽�{>̠�w<<�o_Vt��O�2�(B��AQ��f�ǿ�gy�$(��KZ*Jg�k�U�|蕠���O���y�ڨ����:��c>9���a�z��A�J�Tq&��K(Ƒ/���+1̈@L�E��r�ޫ�a��$e���Ȁ2,\w��
3�!����xbWJ�0�ؤV�m!�@\jo!g��!褏���-���,��gk��V1|".:(��|�UJ�=�.Vm�V��oy�5����#�����4K���cJݚs�&�-l�آ�R���#HE�"LE���ʨC�X��vՄ�D�����x�'����I���/U���@v�N&b�����"׎��Q���_?��WvA��f��hR�ppJφ�l��)������V8zv�� ZmC��^�;d0�,�
�\v}ů�;��<�ޔn�^�)��h�
�{Ѥ�������,~Fs��"�m�q�SF���?/,��5��؃_H��2d�jh'*�q��[}�s"w��no9��Ey���+� 5�b������Z�y/����YM*w�d�+���R�تV���2 RG�d�"t�yŎ=�.Z���b��B�;$1Ke>a��^0e�)&�fy��%�M�8�s�i�RE0?ݐ�Efo~�5�|�_��ֶ��+�e<>&�^���O ����eW:1��]]��z�Xa7m��	Dkߑ��?��`.�Od�'�)�%���Rv��s+I�2ي���Sr��'4���a3�{��>���I����3��>@���/��0^�F\���@�w�ٞ����8��w����y�8*��^�P6��rum{%8Oʧ]�Z�c����J_8i�?�X��$J(S�Ձ�!D��!KHuG�M�j%�����o�U~����v��5�@����ܛ���X��c1�w�����q��_D�W&:)gU(C���:�O���^
:�_ռx^ٝ�g�fB?�vQ܂��F
��<��ϗ1x��.=E)=�.��;��1�� �"N�󜶦M
�n���C?��{�Ң�

��)�XD�1�oy��� �5�Cu!9ْ[^�e�Ce���=�,��8SPO�=k�H��"��޹��!�,�>Et\2�w��tR"9���]6p�o;Vj��b�h�Ͳ*��W�:�fl��P
�|���� ��XxI�X{�i}�,���1N���J��F��d�Hm]V��ŝ�����s��þ~n'	�}�1}�f�%�c��XQ����P%"���oK�T�w4�E-��T=�aF�7/2O�/[ի� 	��"��*�na�L:
 �
\�7u�z�kՑ���U7Đ�'G|�c�jd���TU�<A]5{�)�����T��c�z_\�����͐��,Ob2Q�F����хg�Hy~����7���K�0�����X ��2�B�j���v;Nϙ$�3$�G���
@�ߒ�gൈ.wn�?���D��o�zv��Bn�@2~�n�b��8�^0�PnMЇ��e�5(���N����C��.;=�6�4�^�=ct���|���M:bď��X�!2q�+ؔ��*^������=	��d0���=7����^ۚ�\����{���m�	��r���Ɨ|7�4'3���R~MAmvf�o)���a��gv9�6A��
�*��?��͘���38CF�՞$���O�v�h���������W�~��N���pf�>���"�$|�rqN>Ժ�ڿ1�9B�&�Jh���8vI�g�(��)x�rR!���\�*5$�.]%��hL����ُ��s6[6;Q���-h�,`j�h�c�{Xa>��H-��/9��|M|@J �u����Kv��+L�\�ev�9"�L#X3��7vE��-
�w�_z筇����EO��J/:�S�;��+�y����f��#�7�]��(�����c�V�R^�fב�i���4yw�2"�_�{w��Ze$����@���U��,-ϰŌZ�|�Z6&��Y�R����8�=���+`F�j�XP���U��0am<���n�%��x�]�����QE��If�S�K{ 20�B5���h�9 /��Wֺ���=��å��%�J��(��,ЫS�� YL!Q����Yl�)��9�xܛ>.��U���ȉ�r Qu����OR�ۉ9҆���v8����41J����,���<oṈ��f�9B���%t��+kOq��u��@�����9 ����Dj{/7�aؚV:��y	�u�5�޺~�w�l�.5d�G$!}$�G0�eF��s� �%}�t:X�Uؿ̻���=�U�l�uNϔ�t&����2��_�P6i��x�����͖o�����F��s< "�+��N�S�;W���Q>��4͞�;����%�g� =�-Ԍ�c2�3j�]ޖ�I ��
�덽�9S�$_���1v�y�,k�%;z]���d'�Jo-;�Aَ!�m��1o~K�@��)b��¹H_.JPI���VB��S�R�� �.�*y�cg02�֨���t�#��R܏R�yN�2�� <?�S��ޣ��1�1n��vk�a��,�W/�߉�JU��#K�[�8a�\����(D{�4;ڞ�����-R���/�[jiu�\0����g� ���˽�|�i髹O�d��+���*U�2i@=Y�������W��D�",�=��U'|�[��G�h3��;���WvU�ӱo2weA��$�A� J-2���tǊ�:w}��_���3�����[���?���M��:���棔.Q��~���ec�q�/D�w��!�}4�ޞs�#o�C�1���o�n�)�sj��HN���팷c"�ߤv�ѡ^��4�v7��7���A��y#]�L�*n�ɶQ��`�9M��&RD"��꼄�a�<�\�%�D�C_�F�n�-uf��a�R8^n �v��>ɰ����a?�ˊ�X1͔������\?5i��O7�k��a��r>w�)B\��k��)#T���A�n{���pwе�^�7=�o��#�xS�}�T�+�I�J���X���!��ћr��@�����/NTo�Pj����%˹dq��6&�t|8�H[�X��>P���Օh&�F.��iPG~�n���F�<99��P�!	�@V1����ڬ� �v���pj�7K��O%;r����ھ�H� ��9���]�dk3��uk;��+c��ऴ�L��`����޹��g�������S� 
��]�-�eGS�9�,g�=��d![��*@lq��n��ҡ����	��H9��#	�[UM 踎���5si�bw��qD4�9���G_lj7��0�A��Ñ�PP=���vo���ȝHf��co^�L<t�d�Z9�ӛ)�k�����M���Pv�!���N2Q�xȒ��8D�%y�)lK#���]^4��a�Y���A^Z��bo������%i�]#;��`w��`)K~�<n(~���L�>�r|�k୼���=�h=V�_���.�B�A��(��}T%���N�d;�g?�k��'��ŗ���.�<->�=~�f�!h_���Y��>!�$۴�0i=�����;�"@�*6Y-A0�;ZB U��2��C�j��G_.ep��aµ��x����,4����2�"ggo(�@
%'�f�Ov��̗.�I5)H��T�wGS�̺/�J�D�-O�wh�T�����E�@�p�e�3h]�S�4�b��������V���cи���õrg�`e��ߺ������~[�Wr��X��p�9���sGS�Da�P�Lm��D V�.L�9����V,�V�#�*�<�J�>��)Kr��_+b|��Y��C�Fڼi����CN�B�.�
���no�,Q��Z�*�?2p	��*��<���Q5�P�mP�\*��)�A$ëƈBw���lR��WUǰ £�q^��~�M#U�0�(�o СHZ��ފ�]v��� �|�,ݓ��e|ʹ���4^ЄW�I0~3uA�acm�깲�Z����^b��Ш�����&�n����_%t.%��"�ЄdlQfqW,��Z����X⛓�f��J;��������w�n�ie2������a*�22"���^ ��:�9a�鉶Ew��TI���o�ZT�����Ҋ��_��\��.�X���bi��9�c�e�G���Ɗ�X)��v��jm(����l8�W�ئp�3���{��=� ����
ԗ��I��ǈXb3&[ߞ1ȓ}��|�C��G��۹J�=�=�!��!gCƸ\d;n��uMF�)l����|S%��	�~�|�7ۭ��Iu�j�7ـKX�������c��N��I/��&�J�Iߴ����N�l�I'#^J��kE%��x,
�2:���i[�HY�A�"6�����:�\�����[{�����v����.��<KN�㙻c>�b3G��H�6��p1�2��So���p�|���P1j~`���.�bw~���᭪̹x�c����c	��a�1uV����T�9�pO#�P�u1Ɲ��G�,��3E��p],�z�M�E�XZ�转+E�tw�������C�2*\�_��%��+1�sf�O��U�XL�<�԰�f;������_3bEq�Qn�q��p�N��.x�n}���*�g�x�,�'�0�.�'���I��h���C�=�X���Pn�m����� ^�(y�8`�Ny�Fi�vK��&�������Q����f���H�KE�;�;N�H!i���s (����!H�K��Q��]k���mZ��3��=_#��d[��q·�g&��F����>E��Iu�����mA�ȹ%qv�W�D:��8���i�?ҟ~K��cc����sb�^���X[1.2����U�典H����;����'9��}*�'�I�%��c��bR��3��*��������1�M�6�q0 �5XZ�8ȫ&��M4 7��1�]׉|f����/sy�w�7�Eǔ��ӻl�{��L�?�"C���"eǜ�|x:g�$"���#��۰�����>��!��^�;� �h^˧�bxe�{Ղl�}�^g�q��_�,i���i�[�%sw4�����0i����Q�6h��;"��]��ڞ�v�<��L6v�u�^0��1G�\	z�n~�h6;UM-l[s�chm0F����3�领�1��Ot�I�;��~J�u�̒ ٨.�-����B�(K�K��U������ʳ!���LAPF-^Wk}�(���j�.���5}��շ�(�@�(xL2g�'�Ɯ�Aq�=aX������	��;����'0I�pF�ZsN��$t����?+!/ߌZ��|-X�gK����J�THs�[��ܦ�B�ݸ����Y�t,��p�,]d�5���:�;�H����05+F8r�FXH����#��3�ft���U�VMƼ�5����� *g���ũ/N�tǀN�ګ���B`u��̡z�
$��]@1�`Ɗa�޸eE ]h����O^�ݴE�i~��&�TE�{;:�0�Ʃ���
�Wq�֬X��V/'�N<7g��^H7���0ZE,�C��A�lȐn]��J���d�H��"�`�]����h-0'�`q�-,Bxau˳a&�TȳEj�+�h�Q�MBq��δ/{�}Jb�`<����J�,��uD�^��9�!h�(�eЧ�P�\ɂ��苿���d�������	�	U~b�X�D�� Bgq�V,ᮭ�&]h���#�H���j�\�wd3(�Nޝm�����:���q�IE�}R�ׄ���J���5�:��^$Й
���M%<�#8VɁ�Qb/Nܤpn(��U2�BlY7vd23x�kK�eQM�^���w��y;�E�Ҿ�p�L:��"�7�-(�Z3��)\�f���(�5��U����Ɠ���K�o�*���H�]�ڎ��Ӽ�/��c��-�\�����uP���,=������0�.�]H��1�D�Bs��	R��:�kKq`T���Z�(m�� 8Z�H�Ƣ2�����'�`dp�2n"c}��D\��fjef/H�=L�������W���Ӱ���_)p��wF2<��|�k� `�sX�e�P�40�֧N:U:��l�S����4Q��TnX���m�o��Ҝ��_��S���m�'�O�r�X�I������^���Y�|��s;
O������V�Jꧩ�B:�e��R����Mo�j�2�H�f��BkdiI�^�@�8�� t0�;��匿P��2���u�Gl�<��;���y@s�]�De�w��Ԗ���#3��޽�M-�j��ea]dۜ�T��?�u��oמR Y��rF��n���;�����'F�R1����j���~7p���/�~�N�صk��
� iTe��4N����?E�Z5�,����$^��-�џof�x d��4�������wV;<�/��7�*�@x�X�,I���t�X�*�� Y0�)����č�Y&��Կ���ٺݽ��W��krWD�:�|��i��]�0>�ru<�kփ:5͹xN��*m)��(RG���S����v�oQ�P"=��%;ܴU�~P��
�t[.Ww��H�^(�D��i�+GG���''_�)Y��h�I���S��_Py�D�[n��\��a�ݶD2�KLǫB�ID���[(�z���܊��Q�V������l�6�n�~P�5����6-���N圖�)�;e��?]�T��Nn�j(��ң!�����CX�ј�V�C@f�h�SE�Km�u4ѣUW�,zA؏N��&�� �=@��s�4�x3��h��E�J2�D;m����F{�����f&�3Y/�c�>a�)(5D�/��c´������]��ښA>�\��2���H\�D������T��b\ʑ�8Y�/��,tCgLX]�c�0�O�82�f��q���ߥߞ��:h̥%���nz�cBZ���� 2�Q���@� m�kqJ���~I���� ��ݧu���i�͛�v��(�j��V�!�b��h�3�\ Su������{ E՞t�Y4� �- �?8'��N���oO�׹y�ԝ�}7:p���9;c�#�+��bN��k�p����\���T��mF�8�3*��zȾ�!���x~I���v��&����:o2��q^����Ϧ�\'9
+B�M��:yF��$�w��h�#s�,,1i�5��o����������٨��Wr�b�_E��)ެ�˕�-7�0[�(��X�(�W<�d��'�#Sf�d�x����HZ	��a*&1�G�Zp��!�If�	W��p<�� ؏���5�b#b�d`[�9i|8���QM��wt�b9��Z-xq�	M�9L�[�Q�Dt�t:���[-.��J��xxIG1���nM�㐝�r��/k�[S%7��ӐX��E��7:�=�����P�&.Hu�K}z9���-�;�1 �9�9ʁ�h�����h,¡P�h#�+ޕ��O�ܰ���_@.�������t4�D�j�lp���c$yh��:\�vP�5{�4{��L��>�G�K��*A�t�rg^8x�l4�	*@���h�����UA�d��uag!;2�s����7ز"�p�P(jƍ�|u�+G�=]��F��pɕf�S��|O��PU6ԟZ�G��	M�_<���]V�R^����J�� ��2�y���ܹw,�i��p���4'] ̕��Z∏u��E���|�+q��{��9#�,����M�Eq���/��f?9R�}�"�(چ������D^��?����;
6��f#{�zr���ͽ�����u�.�1��N�8�U��QH.���n���:bF�N����lͩ���k�!s1�W��*oA�neSԱ{�ֆ-h���+j�-t�%f�W3aS�,����ʵ����{��j���赢�ԯ����y�3>����I���K�W֯��:��>XĳC�4���IG�%{��U,�O��ʞ��<6��4ʩ��i�#���)�_��8(�j�~c�ھ��S�M�G2���]�-.���K�,���V�Vz�.�Q�U2-z����5��D�䔹j9`���ꆇ��>�J�x�o����߯��ܗ�U2�IJ !��<��_�!=\o�H�����������K���T!���"/�B�#�� tfD���rbĨ���V�f��	]:�`�`���ݍb
���?�p3�``ѩ�U�%͈-�PΞ�1~��o��;9�\s�1��# ��t����M�#���p��,�P,�_|E����Ȋ��3���{7ψW�K&w)F��%�QQZ�ܷJ�H r�7U�t�$�Kq���U�[�v�<l�ybg���9(y���������r���c�DQ�gK��S�Y���%��~������=�<��{������V�}�8c�;�l�	{_��-Q�����|6�1ç?��·�W�(��˟�y�Ʌ��:bȒ�`>��sɓ�;�8�M͑� ����/�4��=g��P��c�;��ҽ���5Ui`}�   ����H_ʣ�O1�ӯ6^a!����E���~7<(E(4�K�7�%�Ms�;]�Nw��͟�T)��(}��B5�L�M���)�"�i%jw�����sA�%��J/�����tv4�)��������\�w�
搗��0N{[�~2�F�!��Bܤ��t����'PS[--�~AC��YL|��u�:�l��!j���^f�u�ʐ�Nq k��F������/W\�FLOΞ$H�?�T�PC��#��\��W�u�3.�]y*&�g�3Z�)����ʥ|��x��ҟ`���-_1�ٌx�!�Z
ph���*��F���Dq&H����o�4��W�!���a�e"p��[QX,�D]	n���lߏ�W�*x
Ѹ[�#%%$�ԥ��n�"����d�ߘ��bbS��^��c>������2pX��K�:!"��=�V�E��	دV�l�z�?O#�D��7:9�{�L�)xs-��O����� z�	|n��Jr��U�������W���Ρ�* ���B)>D��K��p$<'B���3"@O���E�1~TQ��Ee[-Z�O��ȓ�T�7K��tH�TuG����/�%��,C�ϕ�/^1F�0I��zj�n���l���яi�ſ��P�VҊQ��=q\�vh��Y<�ssXDu&�����
�-��e�S���Oiy��h���~A%��e����/���n�s3��H�H=�X+�!-�D �e�N1���zQ���H2�.�� @8���u7j�	�vQ�	9����?��}��f�Zr�M�K�1�d'Co/+]#����@�;�误M�Ja�<>o�U����b��[7IՔr:=�i7��D����4:-�@�f1�)�UoWZ�pYD"���>пs6�#f#�[G-�W�x�]��5�\@<�)�+�[��<�M��u�����cD����>	"8��㭁��zz����c|��~�"si�rV�"��rI., ��<Zn��.�8�^|�����O=Z��,��� �� z��=�0�qX�����پN��^b�.��g�����5{}����eÏC��K��2,
���<wT(jƙ���Y��L'�pZ��<��Ɛ��\����]�bJ���������ys�o�U (�JQ�h1^0�Kjǝ�&Bބ� ���L��zⅢuF�*wƨ~���E��jz숓pl��Gi�}؏ (7��-�1/Q�2�����
n���mM5�QKvb]A��g];�,���.�,�58*�įO�f��%���;z/���~��F��V���_w4�&���m�l�8��7�^��<��>�E)k�JI�#�\4/���[J'�{i�-� �IW�`�!%�<n��Fn
�"�ů\�;�����ok~�q�.谒�}xJ ���TD��M;�oצu���&F�Np�u��tԈ�E�s�@��m$�+<��Y���䴅cMբ�����"���<f��(j�ll�](�s��%��"˧��K^��~N�O���8�_j��(�9�Pl�bP�`��W16=@0�__B̂��}�#[D֡d�:E����C�9F��������buK�4�0[�8�Ւ9��n��Hj����Үw.M�������S��	4�	N(VX�S�R�J7tH�R>p��۸�
��%�+Sދ�qLV6��-��)+�o��CV�|1;��-Q��^b�`%�W�|��d��Z[C��ݲ�O���֗/%�Ó
o!h���E,�g�Tjw�zݦ5jU�d�[�xA�27Q9%�<-?��Vr6����smb��iW+��a7�<PfCxO��ϗYtj��k��ޱ�8-m�u�rCz4$��v�O"���%$<5�M�N�L�P��V���! ��ff��cehYM���`y,��)���	�D��`�EjoPB�^�V������6h�� �	D���{�$Ɠ\h���8J{�!
�'d7���w9;֤��*�3��9�ܿ�BK���e��쎬H��#Oя��dC��-��$Fa����yę��Þ��2���Q�|��$\�ǭ^Gc>^wD0�:\��e��x�^S ��x2�'?d@�sGq��oz۹���͐xk�ecN�x��Ϟ~�����]:��:A-?�U1�^�nLsą��ơ4ļ�ऍ&ς��x!����N	b��E��|k�`�ATv<���^wRl��X��a���*��%/����՟��Wc&����.��S�v(�J^��<ggcԓkQ#?f����c��QW8�PI��GaGZ
_�,����Y�c���Qt+�w�=U��l=*�W߂���mK��`t	��1�\:�o3iZ�tE0�4G&�P:���].�<ڎ��c��X�I�Q�~3+�l:!h{x�(s�c���v��[!X���s$"=�����x�Vq�F�H2:/�\h��y�4����S�C�\3�(��Ʌ/�o�/�����r�!�h���������$uwۼ��ub:�����J�%[ߦx$h˾QG����dS�fj�_��)磫@N�P?�� d��h�*��$f[��e�r>{��M�fZ*Ub�[�4��^�)�������GB.�0#�6�c
���mF� ��99�g�u��=��X��^6ʘ�J8�*؈��VbY}c6#kT�Έ���Q���
�%���rM�6�O��}P���[6�]������v[�L5����w˱���HW|v��K {C�)P�a��6���9N�^#���+
cY�EF���Kި�I ����	�9���䨦�d�}�.T�hm�C� Ѕ����4���ml����(���Q]d�Sj�)��|]�̽�����|�'�ÜfSK��o-��){���*�#.;����~V��j�¹���^�ar]"��[�Oy�U�T[Ho�iJ9� �{SA���k�{����p�[�(�m �}
�d0f^��ƥ��H!��eR�/��ğf7�Ek���3�r볋0(��k�g\aSQ�
u�/����2 ��#u̯3�}~A�k��0:�T��ɒ(�mC�s���OZ���$�~�L�G���N�M�J���O��2!�T�A�4�d��乯�΃����z�?Ŋʖhw�ʇ6����������;�5�.��%�_��k�����I+�& �Z��h��*�Q���S�a��86������d�pQ��wdn�֬���Q�!U4Gb	��ϯz��`���=�G����+�����t��-Y�$����'�~x��6��OD�R��Ϣ�;#vH�E��#Kjj�h��u[��ǈ��6^�w���W���e�N±��<P9[����rѱ�K�KsI&�'n}�q�Ve�3�(
>5ɛ���Vs|O��!��@J��W�Fؗ:�m��o<��n�e#�v/��0<��}`�`�C���
yT�f_8�n�0Ç�|�����������e�����ƕ��(9[����ֈ��ɡ�Vq��!#'i�D>ud=ؒL]����O���@3	3��x�t�ݬ�|�i"���kZ��(O�	���q��w�5X5}���PϠIl�ѐR5�KM���nT�2����t
���Z�67GT�{�=O)g�O6��0��#�ҁ�[���б.@;(扤��f �K�ci�5���������}<�"��� �uc妫����5��ɮ��&l&6tܟ`H�\c|�	gv茁�	s>�f��
�P�G�4���Σ3�-6NG���y�D���0�FL�$H���U��0������c�ҟ��/��ا$��JB�{���&B�����|y�H�J+Q�+s�2;�0���@��j��lZ��t�*�ˑ�F�C�}���O�	6Ø|P�G肛��؏A�)�z��V\|�.�R-43[�D>��?^�.&N���b�1����,2�Ż�D�F�ߤ�Bu���l<�,��.jSX�
X�%!�Bi��������(:�|�[
�oId
7�t���`cf�}�\��RnW�bK\]��^����7Bk�L�k��W��U���W>�#:�z�[��e)W���T�k�K�7p\)��&�PΧ��j(����a�8�nS&,����j*'$h���4A����\���-U�̙�P���G���/bzJ����sHq�4��<���4�/dS��	�"��ف���;����#��b�wpX�Jؾ�H|Qzs�4cB��:#�jC���q�x�\]����4�y�#ZI�Fc���ֺ\����K����-�tQ	�u�������ZFv�<`ש3L��k��G��?sI���#�:�S���X��jv��b(�r�a�sb����)��k;Q�pk5$q(U���&�x��4cenC/)�-���������i�/���Y+�C1��A�"|����p|�y��O�$]��,�R����k��/w);_U��]�+o�N(��������'Y=h�6c�A`�[>W�����M���V����Q$�"� %�11��}Y]0���4#)�;���AÊ�.N�'zF�f$Z�ɖЄV�NnJp<HX�yg>�v�qK�y����+?ҹ�����ߗ�*U�u��5&'�������==���t|��0/�3Kt���-�%{�-�\�:�u���c&I�:+�
�&9��y��63��j؝ja�.�d)v+ܵG9%�P������-�p�f��<`�.2bX4�*�r��t[a�O�!�Qn������I~ 8Ǚ0�����-�y8^��X���8I=Z.@���T�\�t�� �������=��������h�I��ռ���G].�t��.29�"�}Pn^��R�L�@Ru���~�O�"�J�}v��D��w'(;��GѠ�wa[W�t��m]T�����5����� ΢X�~��v�ѥ�� �"�P��0�"��֚ݲ��!�
��Q00u��#��̐s�e ��6�V5�곥�2��Q82��WR����"�� ���6G>a��8����{!I��!R�֯�('`}��⾿�1��8������h�J�
�����ߋ"�uo[��`!�CR�	,�&Y�X�m�_��9q��`d�zM1��)%��.�[��4T؍Hg\�[�UR�h3������4̞g|U��\<˗���}s?�[Q*
T8����$��Fov;h��#0���������D+��ƹzX�W��d�Γ�QE���h2�Z���B�u3�?�솳��e~M��x��4w��c�nd_cN�VFK.�;�`�V_d��m�Z��!,����baAAҾ�aQϢK��ҽ48�Rf��)���d)2[�M��O�\��/�PU-��|� +vG�7����i ��;l(3�O�E��\-�J�#��Fhx�
*�7���2r��)ڀo;��?���#^��F�5(H*9���٫2Y3��zt�e��c�����fm%U�M��#W��ё�M�%�����㟏=��=��;�x�x�Rs��'b)��K�@.x�42����\k�؈��=AJ\۠�lsJa$��y��P4̠_�
��ƚ�č�xi&~���	�0(�.�����T1�ǎ�nݥ�8��5`	���� �.7��wɓh�	��1�oE� o	Ot����k�|����v�P!h
�A��03�?�ۭ,��1���C�x*2��T�E�.2
P6@WvV�u���`�J�V[
�lcD�B�i�QW=�"9-����cL;����cR B:�S�c]�GD�Ʌ�$�v� ŁH1*�^N⑵��EbHRf�4n�B�)ǁ�?쿢��� �g�q�GM)��/��,�+��hxoFr�k4?����i������o�t�����\l��b�ix�xH;"���� ���ٙ��%�ۥ���#�{L��oo�G�ޛ\�T0��#����D�%u%x-��/�b��&�N	���'�U�t_�_֘�d%�y�����ͺ�<��ȶENR��ⲔCl5�ʛ��Z��]0�5*(-z�(�d8�Z2������B��<�����0�Dq���cS�ŻK�;����Q��\�2��u���~ESy'��<JW���5��E��Ռ�Ir��rw�9EI)�ZC��p���B�P#T��Bun��ލ�rԔ��oXΎE.?
�|����۽�4u�4�"�V-��������Jk<�6�rq|EQ�Y���1�~��av��HN�C�~!��B�7�<��mD]�厜�Q-5�j�Q���rB4�5��4A@�ڜzt�m+;���r�	tï�z^l�C����ґ�-|�h	u���rہR�1Α�[	1�IT�*�8$k0�����z�KJ���}�< ����/�V"9�.�� Q�-z�Y�ol�s��������U=q�m�^�ʊ���@R߯� �7B�F	���?zC��v��*����[r9�{�DFk�H�����u��{��n���i^%a�-��,QQ��f�b'�[/3�����Fw�ہx~��֔b��|<�E����a|�Q����g?ŽC����;r���a`�wΞ��
�pR� ]�nǥB��[ϒG,���ud�gU�:&���޶��y3ǣ�Q��ԊEO?g�[Ma��Qx"�O��xJ%w�2�d�Q�'��m�m����ܐ�=3�G�A�	����u�YBŜJ2G޸�`*s�f��ԕ�#�|n���j>�9����t}\]�y�k�F'Ho�˕W���K�,%M��9�pf4'�4�
ݫ����F,o])��wl�����G��N��h�}�%aNz"ħ"�k�?Q]�_u1屜\�)b�N�Vc�����.��2�GY��>��"&�D�W������J��j�f�8������ׁ8E��U����\`ѝ��&a��ty�a3F,�� Եp����Q���34�[i��G�����#��(1�R�����7<���z����4N�/�k,��(����0��B��K�_
��*�nz�"�l������d�Ca��J��n��8��9\v�7��V�K��ģ�W�0�B�(���_9���g����j/S�@h_~�J���T?D���t
��W���ӵQ��!�Q��v|Y]������N�o�U���0' =v,}����9�	7�ܫ�S��vW���v.8n[��Wnr��%�TH�� �k8Y@��w~�`YÁ-?�B�?�D�}h�6FH��δgg��8UKR����W�$�NLd��e�N�h���	�f�N:d�)S�O�6b��%�l�w#D&O�_�-�S�>�׌~�Fra�C�&���.3.>w�gl�5�j61�fޔ���H�Խ�+D@��0�g�/����=�Bx!��~WM�)�Wi�P=�7^��`ȂQg��PLHG��%BRL�,{x�(u�:�l}��&t��4cN{~�(釉 <�oJ���J�6jH�F�o��d�@�E��8=k�
�ҍ�Y57��/��s��'��<�'��e��ǈ���Gd�"U3쓙��|��c��* ��ْ}��*bZh+�K�^v��/�v��0�P�=B5'�.+M�ZN�H0L��/����5�2Q6��n3�Dw7��^�J�P��7���CKBT�z��dOU]�'<���,�j�����maJ+o��[� H@A���C��P\����tK�W̐ǹ9&�F�Ā�0N���4�w�꒒�-��We���Q�b��`�'@������x\�+�p�����@@~��7/�ʄ!�@��=���m�Da;������āy��)��Gǋ��7�� �]=Wd��.B�Ա���8��i���P:n���m�<ɮy�j: }�Iqڌ�.+�s��{C��[�ti8��>	�o��I;�wI����a�
.�p��Þ�L�o�P��&<N�؟�&9i�-�!�{/9�	�3/��zaU��Ձ�2���s�Z-H��!�X���r�:@�/�)�m/bo�N_��bc���L��N'��mh��\[��9�B�-B����"��bI��uɍ|%2�)��֕�$���Е�o���O�gg���!���F�Q����v�v�]�N�ػ��j-����YL��7�� 3T:�E�4����Ѓ	d��
1�o>�.��ɿ,q�\�	2@��,�EV��Lb�Q�ur]8���8�򧘩p�|��NR��k�9�i�Q�6�K���ߤ�̚�4���gau�:�K�>��W��-�8>�+w����F��� �Z���X���\�齍t�C�x<c�|�0�&���
�Fr\X�"�"����w1�OC�%g?,|MLi��� ���Όu�~���ⶮh�����֧AdQ���E�� ���P̹1�,^l�u�x��}�dt�ܣzx�)�Bn��/���4|����{�S�L��S��i�Md�HTD3l�H�tW�������fX����l�����.��s���y�{,-#q���hfI��ʧ�ݝ�/����.b�83�N���
q�-M/�S����{�@-@ҐW=yUM��W���Ƕ�k�|P����@46��m�Xwe����Ŕ��u��:a� |'_�{Z�e�-�U�.����w�яt��N]h�7L.�9)�T3u�j���������VG��&�|��9��B#��9��Ǩ%��L@��H)��R8 ��0�SwP�vP�):��ey�����k*is*��o��rJ�j�����=lUės �Od��c����y~�O�OTm]��\ݠ�<GЍ�F���-����'!�O�~TPj���ih�߽4Ηϑ��ئa�c�Ey�^�	\ܘ����o����o����C��E��xSХ�)��2�-'�D�q0�1`,�|M��4If{!D�%+Gg����	^>��0+�\DP��m֭����R���:�ݦ�ڡҏ?_r�l<ZV<ݻ��+M)�< 2n>�i�Ŏc�$0Gꈋ����T�	�Q_�r�����A�|'����DƤ��f�0F�iQRf"��3����[�|.ۘkDmx���Q�;$^U�l^z�e�W����_�50��X؛�l��nZ����w����(�'�\z�>��0F��_���l�c��#�h��N��6_QV[guJA.q��J�bhF���&�g[��M>���f�J�e�A�=�֡�6�.��lQ<������>�ۢQ������T!�.\Z��Y�+ *a��X�h�Q����C��3.�!1�¼�08>�B�u��A���!�I�@����vI&�먽�[l4<j��I�.S����~�(��/�E�F�
wq��U،Ҹ9<P��ˆ!B�`�A��u�D�y�QF�K=_GXt��J-oḕ/��߆
��>~�Z�q��*��p�
P1U������T)�z���&��Ɠ��N\L(����? ��Ą�&yf����,�]Ъ˧6	<Z���r;	)���e�a�|���y��_8p���J� ���"6���M@�[�{���a�5������h��.�p�S�oa�Os�T�L��C�c����G�L���~:@�,8O��ڶ�[��_�=?��2��[�F��K{�0��2, �۝B�1��@�r������36U�lr��.���D�p��e�Z�o�;'���i_.���-�6�2q45���Ox���!�UC���*~K���N��yO��D��S���M{��/�Ȯ�x��q	Izpe��dM��nl�EB�)���z}ͦ�R9�b@hC&�Bʿ�X-h,�ˏw�Ř�Q��z�(��;�U���u+v��BO�Na����ȓ]���愒Zd�,��=B������?��\���2�Yˌ�ֶ��N�4��fP��[M�����=�Y<�nUٸ��q�8y�t��� ك�b��̓��T�q�����If5�O/����Z��Ȅ����6ѣ����+��vD�5�Ǿ�}���S�8�U^���[��W�/lM'�y��U���/e��q/��5�l����^�{��K���s��TO�5�=Q㋟��PLLdI���\���pq>�gU"'���4X��9��P��ӑ�/�p�ϵ�m$���?d#�lK��G�~��H���)@�zx7��6��]�j������M���ʍ����$�WE;�s��N������w�8�o�_]��z�N����nx�%7I���3˳�w��A.mp�!=0�';1�D�?5�C>��:q�/$}�qŮ5*�J	C�1\�w�Ҕ�g!Oa#���V?̨�#�8�0aׁ��q���Qr�����ECy�@f�s�B��}[����ADP�9��18Oy%���{���wT��mv�7��I��6�][tW��}*V���R�E�u ��u�w�D�G=�ԋ�����eP��K��T��@�2���Y����_%����)G�$7�d�xJ���!�i*����lK� �c�`(�߭����W�	��9eMc%�-�/��b��(�g;�O%3S\*�;�n��2ք,뽑8!Gk��aD��
� ��H��3�*t+��)��S")�QTrGVT�;��{��k��Ќ����DC1���1Y��\蕪@�r�r����O��c�Ӽ��+�d%E�	:ͻr��}u�mO@%g� 9���މ�X���1�$�+H �x�<q5�sb��cr��7?8#+En� N�y�q����Vxq"�j�;�(�l�.<�w��N�rJrX)N���,��BM߼cF�Gc:�E�]�f��͚O8[u���Kw����v�7��.�`��� ��ADg�I����(��cDw/�IM.���4�����v����������j$�IOC�������M@"y�v^��6p�����ێ΀��oֹ%al�؋��r�	��l�p�$hw���M:rƿi�rQ�\x/x&�YC�-��2��;*�ǩ�,kSXu�t�t��צ��I�vԔȲ���^R��5�JE���)���x�+�^"���ܲX�l������D�_v��`,���h��r3HJ��v���Y�h#�	E��Ԅ�S2v���`=�PA�����ր�4�l���W��F�����R���(:��(�aX���l��D�7��ٶ�����8؇|�ISk�v:�ր�.1@;//rN��P9p�3%��5Ya�6�'�d�L�h�7��bBW�RC�}�'2�r}I��u�V�s1,��k���K0<:�}j:z���2G����>��w1�'��+��
�ۢ�G��Y� �P�ZOU=�o.�,|"y��>pӁ�������G���f���.q��Ь������'�V�Q�k���m,�@��R �yw�v�����Y�EhH���US���.�xh#��a.��R�����(�~�zQNV&�N���x�]g�mD����}�ѵ��M\iM:�"��, ���C��l���\�����-n�E�_qD�t�.�B��e��f�1_R�hI�[ɻ9�m�\�U��^����h��^'HĂ�8�m�_{� ���	�ׄ�)�bT�_0K�ju~о�"�Cg	�)O���nLx����侸�&��q���J�QO��â'Q�g�)����>�O6���Tt��H$oi|�h
d����k��'��*ٍ��Be!���R�c1c
%��S���� �	��]|30��|45&��O/2(�{�m9[�DT��uX�Y�{�*\(b��vI���j�'���9��0��}ak"��A3>}�Rq�ߑ����;ym�B&��<+C��c�?�xQmm��q�w�ڇ;̗���1U9�ko�l���x��K�[S��.���\>�?�N���3�"R�����7pN��-�6�.���F����̍/�����(w]��i�T���� t�M��)�G��L�P���������m�Sm�܄����� �&OP�}Jb�~�O$F\��jO@[��y�}Ys����\O3��V�}�U���z�@�x��>��k�e��^XK�HKO>�k�G5���T�_1|����m�g���W��#z��mv���SC��vn(�Q !�&� &�)��'ŤT�B���E�R��=&�WfgmwW$����N%� $�C)��XUMqh�7gfPS�K���� �c�$���D��qDI�9�N`�0!_$i��he=2]!��F����E�W����q�Y`�O�D��;�ο������� v�Hɓ�d?�v	�-��r��D�O��1=-:Q�����w��^�� X �A O�[�
�Pl~$�|�x݁J]w�g+���YZ+M�Q���z'�t���%d���O�B�Ing9 ����5�:�6F��זS�-�y8�yj���@����L���37M@�Vw��D�7훺,���-�<��^A�#���7�fz%DLD���,��7��^k���Hre���d7E�t	��s6����:���VukGW����ޮ^
���js	(�����!+p!�m��?
W�4��n�8��G���3���$	�R1�s�
Z��{����o�G��F(�y��G/�~dp����Qd?�%���s�݊G\N��v�'������v�����P�$��SC���H�1�DS��19q�?�������� ҹ"� ^��GGY3W�OѼj�� �"oT-I:kS��0c^����ס���>�/,�Zքٜ_$��E�_��U7�B�*����,3d�E�~�˖~ޛ��M˪3���̚�<�|	����"g����@96�x����!�#0 C4T�/��U�7�Dw����=�����mS�]�s�9��z�EA6tByz��F��W'��AמaS�����?N��l&�/�|���&�Z����J4�<��9_l�nNǪ%��W�O�~>WJ��n������NHe�<:̵�W����zP9���˲��޲�!��-ib���d_r�t96|k��8i���ÂE����IA�q.���v `t/��*խ�8���ν�I��u�����:��X1�y8G��F�E�Ne/M C�Cc��M@M�EMa:\�m��)�TC���Gp�:����+|6�=�ޯ�,HC���kפ+�]m��'��4�}���z��ʽS�A�gq�
�1�}ΖZs&NC��E2�N�m�.YB��].EaG_ףn�Ry���ϥ�/儮��~�Պ=t��đ|a�U����y4�Us˺�����p����'	�:������m1 K$w>W ��i������JX�K\bQ;���'�ֳ�Xb��<h���
N.*�����Ҧ�����~	�b8e�[]�"6�St�iפ`UD}c�����69ץ�4�Yby�\�x�����ٳ-ø��Yn`l���B�b��&S��e���tX����*x=V���P{���۰픇��}�9A���e���
���;)��XU$Re�9�x���t�
���)��O2/�w\f�#] �3x��_��MT�"�δ@��y���0r
X5������`x#Xa|�Ġ���	�e�I�?�*s)"�X�ԛj{s��9�B,��23�s��7K���Rs����'�4mq�s�/_�2��D�=Y�-7�Y�)� &/�8� /�hp���{�OP 
��f�<�́lD`���v�$άaf[�bJr[�ױ@(��T��V���2��l�%+N��8&��'������xi�]i�,P^v88L ���$]���eϐ�i�J��p�P赧 l���kѹ(�r�.mQ!	�ϧ�Oz@��Gq�U� �pו��ވ�,u��ܞBش@�����s� K
F�@���S�d��W��<cz���1؛D���V7��͵|#������x�0a���+ 2�* �8A�hz�u�-�_���Q�C�Jq�w15�]�mxfp"ju�B�ҭ5��f�2H��W��'X�d8��|w�i�r�E2�i�'��,S6�P���c���Y� ��lŌz2�����_U�f�>SX3�EǞ�j
�Z�?g�Cf�N��d[R�eV n�P�ZV?����ݹ��c0���Ki!�kb!b�h�բ�]!�t�t��[���,Gvz�0��r/�R�B>]�}�Sܪ�s%8��N��Te���`��"�yMq����i�6b?��4�#�d���y=i\yۯ�g�?�[p��'ƥ9i|A�Byi�0�{�ߕ�s`w�O��j�u���Sw5��U�Pyp@��q�~�\jG�{����Om��sY{�+��j\��C�,���/K�:� � [�pv� r
P�<�N�1�v���)ϗA��[NV�,hO4�"���p�����8O���6��F���m�YΗ�&���2?����,��!�!�!i� e�l�)�-�ܜ�d�K]I1{��02��ɿV̖=�iS�^�i�О��f�E�G���1j�}�ᛖ��*ȍÕ�H+�L}��/|?6
�pY�u�E�f�P�,8���Uo�皶)��q�H�^Z)ߙOU�G};���nۆ�U�w���[40�o�d���Z6��"��ݽq� �V�{G�N�ϡ��=r�71vСN���+�;�`�����m)$�#�hn��yJn�d:-J@-�e6Z��yptM�:vP>�D�dr�}���C�M�`�G"Z��Ȏk�M���S���^�>כ7�0�\[�hl����t����}ٌfz���L�'�ß���ǱW���H�06y�����*Z^�c��k���?"��TRt����İvl��^4k��e�
�~��tMC�a��.�Z[��i�c�U-�D[yvPg"xOgC�j��j�ϕÕ]EW��n�#T�#,�[^=������l�;���z�o��w�6����iuY��>[��R0sS�wĠ1[0~Y6�V�&֢�7Kq�mbu�7�ڇ�,x!4t� ��˘x2v�f�,
�~��"�������,�ﹴ���1��]���Hl��Nz���Ǯ�C7�Ŀ��T$�CƗ�w�F�����֣�K��@*�K�1�[Z�Q�-��z�n��1��36�3*�(���.K?0`�lve�B�4O���)탮[fT��[���w�B�[�T�D�q�]f�܄؈�IQq�]�'0����{]�H]d�:�g�XV�֞��P_õ<Q�{)o����x�3n��TJ�r�Q�i�D�fA&^zq���β�g�/q��HXl����nC"����G��y?F���h#)d��I����z�$��|)��~u��l���Wp_<�ēQ�G��n�Q1�%1��A�D0��z CPpl��&6�`�e}:��)��:�C[�� �|!-^��_Z�e��6]�����p�̃'� _�d��HE�!*��gR�����bӢY�Ϡ�NS�(��c*�C��i����䎬�r�+��IH羼�
@���
ν .i~�� T:�`#��Y�N��W��
�e���E9��O�5�-��T�v������N^+/*n+d�K��8;X��"�ޏ{��!V5�~�f>�M~��mo���~��e�Cdػ�vצƎ�iū!�3"�\8��J�@�$Zvwr�K�&D����yP`�n��1ݑ�8��.�+�zR������ס|����@��^K�G�#2���@U�����,���`��dm�A����ޠ�rʅ��MK�1����P����?����$��<�ɫt��!7c�1�����!>c��D�Z�D{���V�"&S?'��I��X[��/'�ی����iQ �e��.ml��p6�q= ��(��G�$��4��Z��Sgz��%�d���r7��>�(�{>��,Ԧ�PC�K޽�(Tr�.���!6��A�f�V��|C�W���9u)���P��v=������
�_�К��^˰���$����)|�R����q����#$/J�q%��㨽ze��}lXU��0��Ts[�پ�#�7u�f����x��w�BwLB7����7��^�>3��/ݯo��%�V� ��* �T���r��x;C՘}9�-Ҷ�0o͏sJ�<5�!���p[�k�Į�
�%����{:�n�:&����4�҄Kwe�܊r���i��C&�&���ޖ1s0�t2��1�(�,%n#g{Iqߥ����5��&�K8D7ncXV�ެ�y�eG�Qq(��}�jZ�-U���L�~E�+��y;.]T��S�H}�lE:�s#�рW�TZ���]�wo�y����:�[��!�
��M�-=6��v&Ft���3����!J^9����æw!�9�%���UE���zc�#T��P ����n��\J��YfE��"�6Xܢ�!�1Aɭ7�և�<:"ڟ�q�9�jB"]Т����b���P�V�	�୭��%4��c[�����v�-B�ZvW�L	1�~rd�V��7� h�W�$���:����'�јYi���G�Q"tE>���v�`��F�)�I�����n�mb��
C�3��S��˩�{C�>�Y�d#|YRPg���=���	�l��O)�G2@����!��-T�]nґ���4�~��l*����w$�.�@d,i�[�|�4�4ԃ$�g�h$=��!ʙ�6P�aQ9ϡ�]j���0�F����U�-�����q��?����>T���.6h!n+�u���@_%GQ�A�3�9�ko?��D�q��˪B�Ҟ,Z��j��UǇO@�]����Ǳ�sy�*���O�����nH!�7X��sVx�H���
��fT�U�S9Vl���}�@�të�ݨ@u)�lչP��!p`pY� ۈ��c��(�j���\MX(��9�ay�yJ	M=�����\�D�
���rq��x�c��q i�:z�{L��r]�,�I|~Rm�BCzl�-#]���A� ��O��<��ׄ0R���ȩe�#� �447�l`�	�t5v��*�OxqhгE������G�c�r� ��s����"��di��I�/Z�P"&$ϲ4"80ѱ��)�V�Go�;� 4�M|Q��G��4@O�x-�el�� �w%L%E7�t|+��yH6׀�e�9�^'�	�fO"g��aHG,U��CIw�V���^�[8�`�@��	�e���j*�1\Od���h��Ҁ�C��� 롿��>}���çO:�N�>�/>�D�K��񃲕����ی�M?$��"<�i�Y�Ի��	�$0vcL�9���S*�����E�Kr���0.bgNJ�H2���a��Y�ɺ>O5�'OI|�e��ktA����P)|� .�!��Z�Bt�w�}Q�߻	�b����I�����C7��`fk��G���Z �7B+h��4{�����9Е%9V̘1�Q�W85�V-���'9�q�dn�j[sN��	�R�R���
G!{���K&VS�֝m��xi�ܤ}`y.���p�}�A��s(4L�su����̚��Vm�mx��ж��Hb�����0�;�a4 �e�"j]��:
�4����¡1�_��[+���*�Ɔ���(D�r9��fF~!9�8ɪ����ʌi�
�0�sLMIe�%��>5\0�H�	kS�W�رƄ��m���?�(�<������\U\���l#���b��#�/�����^�iΖψǑ�ܴ��9ނt�0¾��aՂq��ؒ��1K~�-�0��j��ֶd_�3����3�@F���(ᇈF��`���� ���:��P���2��\*S��tM+���^���Y�m��K�DJ_G0���|�����M`��幂�̺�;܎NV�eh���hp]�I��$f4�9�(�u@�Q����k��w@��4���l{K���mP
�[Dpo���H�o�b��gpc��mX(؏C����W���Yl�:,�5�"�x1�o�A)�c�s��%�0b.*�+��I�I��k��ݚy�s���I�C�m;��ʆ���hј����m��7�]�Y\*��#�-������w�l%W6z��;΀�zj<:��Q�W}eQ�b>��Xg��D�h*k�6��e�o��i!ܭ�{�/�80>c�p�MQU=A��0�28fъ5��Zn^��yL��N;�(Ċ�o�{V|��X'����wb����9qӻ���W#���S�e�b�A��`JYm�������� �Z~�M�P���4���}��c�y���g�|��n���0��G�.68	�C�د-`��	� �<�B���a�P4�7;b�����.�kCY�$P�$�=%~{B��7�P�-�0����c�^�-T0)H(��J�[�7 �xv��,�����p�ͥ�Z�P��-����3��8��p���Y��g��N��d�[��	xIBjb�n��4Q{.i�+VH��]O��9 N0�3Uj�s*��.�:P)�	Z��zw�ق������h]�G�yֵ�fl���ߦc'8&7`����W�z��@8���8��(q2����/x�O�8^	V�w�2^����y����E��iP�;BRb
D���_�1���q*�	�T�����az$e3&İ@$bA7�?&p7Dkŀt�@��x����2g�Ƹ�U�JC�i-��Z�hs�v䷮��t�����_�����L:��tf�6���3�+�>W�ryJ�桮V�%�`��OMB�DHCA�s�1�����
M�"x��@�G>��z2��G{1�$�H����((�ĂE�JZ�se5�p%r�8�S㴇g�=�D@C��59�r�ꚣ��~�#��n&W���+$���K�k�5�|�e�S�uC��#�l�[��-���;Z��d�s�q��!?��ބ,�s�8\�|��9���|���n������{��7��y�1�][2
ǵ�����=�F9Uv���Q&�>�U���N���Q�mfH���mq�����j��[]�?r��!�!�W�֓�@�G3��j]k�?4�;�ڜ<�� _��L*WM>��KL�dϹ����7���K�B����[�
u3��E��5z�Ճ���f?zp*���|˄�L:~��6 @[9�l��š�M�2>S���:k�/�$���5B,����)����3�M(ƪ�w&.h��+E#��Mx9�m�F�j~�S����ʯ���H��Ǭ{2�E�R�4ڸS�!����-�ꦞo�t��CS�;k�7��|�V98�����Q��m��~_/���h�աsPAd~g�9��U�(P���U�G�ƙ�D��|���[u�
��|���ǅ�u˾y�LJ�(I:|	#�b`�7�Q�\��/&Ҍi��驃���J9E�-���^�S���Wm�qړ[��r��c�\��9�R>�<&!�vd�@�P����>���y��붣�T�=�-6���J|�8��4�E���Ad)��<?���ICymB	BMRe�F��H}4Y���	�K��t���'�D�=㩊&S�4�M�3��8l��Fo+��q�&X]Z��VJϳP�H���¬"߃xi?3��Ȉ aY���Zj���tsR���/Y�j���EW'��ӭ;��<��	u�k�s�u|ެ&X()3fk��bq6b��}��X+?R�a����1&�e��*�x���N=ӹe�,k"�b��)����eە���,Vbn��c��dD)����Ҡ����I?Z�Q����-Yz�Y�~��� e�I]c�),N!w�S�&��J*1�;�e�u/�V�¨iI+�Z\c�a�bc�n(J���38�Jt� <$AC���M��f�F�D��~���N'"{��he~fdN�l�)��&`��ot~I�Y�6��J�d�9�L�� �Jŕ���lΈ���M
�Vq&Sp�ʗ/n�׭�*�9�fx)k�~̂��:,�ތ0��y�hO�Y�� ZP����}��cq�x���A�j�rd/-3��C�H���_~���퉯fr�i٪h�Ć��`��!g��xv�M1Lg92����� ��k�5s����D�$kN<�T�zq*�`�z�,t�7oi>���#a�UƊgE]{��Gu@���f'`N��ƻ��j�w�7�Q U��"zx���v3]H�h2�u0����%M��?q�{DD�N^���k7S��].;UhT�MkZڎ���y���o�{���k{�ʏ) ��6�3M�	��ܚ��^���l�v#j��9V��0I^PC2-�PwO���( C�Dv�m�����WK��X��V�4���b;՝�C�����	`�x��=[�7`O��me>�YM��_W����㔁���Hhr�5ә.dm7.¶��TB�ѕ�ȎD7e�M�����#�<�P�B�2�z�Xy�v��P`My�[�-��e��hPjL�����&��B��X9��"w�ɍߙ�������ӅI�>SH�?YS�n���"Td�zY_��u�)�Or/6/��y�k��fF�*���wO��{$Jဃ��M@NC:�ĖT%׸Јz�~���yg��֜S��u��{�}A�'A2C�~:h�Y+f����G�+��88��C"��I�خ�_tk��`�bR�,� 1R�O@�c�}�[�}ZjDt�8��@���h��`F}�Il�^W��>o�qf��9Ȇs�����V�P��\��s��Q�_SF����_Q�8��I�>:�׾
x����}
��E_vP���Λ�B��湱�Ba-$�3-��WN�]��������n�Sy��8����*~?�s�"o25����%��~H��G��>�QTE�w�c���4��m�M���"_��I�"�[��Q0�'���0����O�)Ea��,`����ZP�c]G�Q'��-sd^y	J��[ȧ���'�������?/�r�\�m3I�;��ˀ���u�_#\�8'{����26E�TOl�E�?������I6f_]}�3��R��^F��ʻ���z����W5��ۦ�;3�.�7r��r��pUe� �|��z��s}�^A#��$�J�ۭ����=����v�[G�5����9-e��x�A2IP֤
GAt�[6}+f��=Wfl�'�N[��=~�͆�U?�k�Jvt
�5"�i�#��=�Ȍ�k�א�O�|k?���B��b���[�7�(��n����+�V��m�~BV��\����ʗ3Eu��;#��O��a��D}����,�����%����ѯM2PT�k�tCmCx����Q����+�kn��E冐/;��K���ϼ~	��"jn�X �M��p��P��	�	Q�oC�A�lA��_>6�A^P���%Z{�x5K�
�br���4l�D)H��r������Q2����T��@^H#��Auҵ�VV�d�i\�gg(o�ې,�}Wwk��2>�����
��F�zQ�$)�jgpR��x��O����W����9mg��v���U�?u���t��9��/-�w�x��s�;Jd�o��b��_ޭ_/�U�����ʅƙb;ǋӰ��7�ůg�>\�g�1�����<��Hœoa��,�Żm�p�ٷ��&C���:;��`6G�z���ك���s�N)N�n�B��TnL�W>-&�E}p��Gh�YҟƯ�D�3�X�ꇏ
���
��ȸx[��F4��R��FJ$@���O8���Ֆ�Xt�ea��5��c+��d��`�Z?Z_��s���8
������.��پ�'M���8��u�s%@��]���h�Q��,/���H�y��K��D�W�B������ ���OՖj{��m�.�ꂶR�R��0(dlzNu�K�b�=�M��`-%(\����.p���²cLU�S��/؉�m0���R:y/?'f2���
�����!��i��-�aRWdj�,����R+��ָ�|�K�2�I�G	Zc�Ls��S����;�q��M�n�}�\K®�� 9�ڳ���s��ƍ?��x�7O�t���{�H�f��9�=�eAS�� 
M�-2KM�oYZ��� G�YV'YQ�M@���OxytS�W����@�����,;s \0�n�7�fo�㴭���:��N�X��#�U��1YS��WG�|wy~%��4��d�ަM�u����C�%��F����HP_�DK���]��$4�ė�79X��^2�&�Y쇚Qp�~Tt`B��/�U��xaj Wtuh��5<a�
�
"Ҝ&� ��^0�o������f��(�'���h$O0��V �D�� ��φρ|�}���l�E��n��R�m�nӑS��O���k����<�S����0/H���~ϒ}�M�qQ��{HW�"y�VX��\�d��:�����_�ju��ħ�H}35��Z/�##�\3����p)�7r��y;�/D�<S����y��1=��O^���W�*�	ʋ�z���L��u��U��"�&�ZGU�@�_܀Ш9�����9�9?h<��*Uܟ���&�WXB��n2"�m��@IE��=G�����EF�C杇}���\Y5Yg�p����*��:tg�ٴ��,�q�a��k�Kf���<S��(��cGݑ��/�p�G	l��β%���XZ����2��g��w%Q��XR6V_�W�IE�ٱi<m��{β�M�J��ל#�%!��h��/9?z�O\�JIt~bkl��f����K�i�l�X�����%����C�k
��u2X��-��޸<�r8���t����f쩗�*|���Z��žFg;!��W^�ċ{k=9;Т�4���p�?�/iF�'Y&HO�.κ`{���Lٲ\���;S	CI�!�&���"^���X�exoE�f|�d�۷�,��HI8�C��ç�z�Z��i� W�(�G)��u�-Զ�A.z��T���&���y����r�p��֥⿯�/�#Bg�̾),�L�'E�L���0��|��`�~�KK�ö^C9�VD����4)e�H=6ng5x"�.bb�!�(��^\g�c	�:)�)��W��i"Q�n4��w-qƒ�������H�lE��c8#��KRL�9�6Q�K ��DH��PF�q{\��k��� �ʀ��!~�V���*�4��|[�oe5��=���&G���~���;���@h�M����5�[b՚�c	>Vl�1jR*~�۫\�ɣ&��W���AJf�Ov�r�β��x��j��([`� ���iί�y0�@�[
�f��j��6X)�����_���A8�'{{�����'�V�p1��F-����C)_����!ޔ#���M�Ŷ��XX(�5BPp�-��lyb<��ܕ�GvjT�)�?��v`�~!�"�C*�_�:��䊗J`�:��чC�l"�Jsӹ$�u�p6*��M�{�P}���x���w��"�����JzmL��H��C�$�ð��̨�v^|��:k���K�5��J�c�oL*��5��(_��$��n��&���B�q�%��v6��v��� "k�E�\�4T4��Pk_���1��-\�EJ&45s�UA��՝�7 8s�]��ft}n���&誶� fڡ%��7��M��0�`�t�t�am���'�M��]��Y�O�,Cm������Z������ ֚$�c�긬m>�!��0g�&n
��B_�Q{���Rˡ���YCc�0��f8=p�CՇrQ�P?���=u��T�)��uG�|�C*s��:M�a1��EO�F�ZC�p�+�7Q-P����(&�}FyϢG�0������{�e����m%�z�Yl�%��qO �}��w�b���X1�(�œWM�%E�ۖPJ,�c�)�j!�~; �?�+����t���s�O��Iܢ�{m�����%��Q�E`6�ƙ���ʦU�n+���,K+˻�[�$��:�K�w(��]�oW��㙚L;5���ˮ������t�r>�+u���w�RSbn�Vn����l�b�C�x�WH�
�d��B�TO�K����H�q����J-vV�g�"X�j�]X���x@��1f�4�q	3�-�SUŏ�%Ǜ���X�w�q�g ���P�8~6Hm�7�^��Y�/��cK�(�hR�M�=�V�d��'I��p�r��.��*�����5�	e�O/�P�d���6P��Y�Ȟ�'����ohQ�z��	��/:9D
�ar��o���E�&,�TR���C�����j-XL�X3e�#�[��6�,�j�YA�G��}V�L���0,�O�cW�P�J�<u�9�'z�Qn��[N����N�84�^������O*kB`�ykv�C��6|��yt���!ͭ��4u����BA���
v�̒Y�Pd�3*���`\�;l�B/�������~)RA��n���y$��:�QI\5R�R+Q;��l�ch:rR����t�p���L�~�n�k{�����mJ�"�XLG�V���`���� %����iI���qS@���v�kHǒ�Ħ�q��n�E}&���
��w2r��Xc^2��M�ۡ*�H��X>d��dlwƴ�kɛmRVdx�W=���(��.,d"y���>?݆qQZq���� Ǳ����LW^��$BM#{�%'���W�v�vO��M8�3�U��?�=㖆�u����J�KOB���T�钵���������w1���&����a.�r�oQ"ނh&lQ��qE����r�'���`on����[����YV�֙�d>|!"�������O3.{u�gG��0��P(�*�MF{ �\��sjݺ�.��m�A���\�_DX�����Uz�Q=}<W�K���n	܀�#v7-��P��yhn�ՏNf�7�X���z4X�~�#׀c2&i��2�T���]��*~Yw�c�ͱ&"�����\7�3�PJ �=YmV�u~s��R��4S�R�KYz�j�Ƨ�</��pR�HS{�M�@�vWF���=��ͼAYu�|��Dg��_I�mI�����K�SZy2�I��+�dX�o	��W(�"~�qb�n���蕄!�"�4z�Ye�̐4�-0K/M^zj�+���+��N@�Eg��Q�#y�S;jc����!���2�M��NC��g	P�c�%R 4vE.�i3�Z��q�W�9��R����n�h,T
�k%��:5�}��cB�W��6���|�#�]��/���S������̓MKX]����]v�c�?;|�b/�/��oO�qHyH_P�ܗ�7q��E�H���=$b�4%�[Q�#��u�����6���|��:܆֨z�!��1��q\������ıd'�b�64@c�Np*:�c15q�qC���g �oѱ4������mM�\��ʨ��cH�٪OK�l��z++����R9�JG��y4L�L�����-#B
�>x�-�G/��HX�}��(u(`�Ź���L7f(5|zZB��J�Q:/2�zkJ9��#e��if$!��5�b�?PX����h�D�Z�õ�v�����FDz��a�ͺl�\U�_�	��n@���%��	�z��C��h_�"��3Ն�`�8^��B�y���	���6jm�X)u[�TUJd���زR�f,�Es!c�)ө��yN/^��]�`GY��!4�:SzJ���1�]-���-���q�ym3O�ӥQ��jS���{nv��8��폺��>FVu^��Y�B(�3���S!��C�d�~a�	_�W15����g߹�-���ַ ��^�h�:H|c3#yKm�N�e)h.21�����mi��xh�S|V��4�:�S�֚|rA"���*���)"Tm.5y�M>�M�����>W҆�����4�Xz.��z���o�k����.�,|6D6z}7pK�瀩]�
�C!�a�a�tt ���&�쇸B8���xli�\�F�l���Ms��?0F���2�?*��V�wM����l߂"�QX϶�=
F�7!2���.IX'$�ڛR���"}He�&�} �����vJ:��\�à�	�g̺��PaG9������e���P�/��u�\��!�(����m#�|~�L� 'K\�����:�kĴ���A������pY6W_�?L�d�:��X�&p��B(���ʂ��)�Nr����_˩�7��&�	��f���O4�����>"���`�.�4�ֲ��5�o�!0�����#;�J$|h�Mt�~IY�+�/��m��0��7�0y8�^��Q12lX["�	ަA��z�w�u6�ŏGv�}��t������d�����g9��ڷ�v�nd�е��{��|́��'K��>6��Z�U�D���Z�?�[\О���Kr}�k�M��Vn�x����Y��XX�rJ�<�|(&-�/!ڛ�54N�Bl�`�W~8���v�8��~�M�~9���C�[Z;���6O���e#����
�PV]�cN5s�[�Y�	Q�4!|���=�[�<�0� -�i%�^e�R�*�p���ֽ�k�58�#�0�.����ң�9���J`B{g�4r��iw�7��CE�(�N��v\����� �����r��e�ֻ�	4�%1���^�m�奄��۷uN���U�����p��M3��ș1P�GJ�`���-�mv���a�I���7��<ǂ65�'�Sd�V���Ѻ7�5�9++�O��hvfGž53�z�� q��=�Ru�ɴ����{�E�b�:���0�T$�:ֵ͈�!&v�Im��7�dEv�s�D�mf����BR\0���ɇ=���rZJ	C\I��Ŗ�A�9�ֵZ������Ǚ-��͗���_-#�uC^Ӧ���I��'�7J�.�Q�N'�Kv(3V_bCI�19���{K��*�4��`��a��;�xA��V�#sM���3ߟ��r��C�b��Z�G*ѯ����@�<y~CS�Zyt-������b{_�=��Uz��ڨ�o�%|�S��=@��}n��)K���(q'�z�B�)l�|���~������{<���g�B�=*:���哕.]7V��MlO�ʪ���A���0��T�ݽ$^,�IN\^�wN�ʠ��?l�L¬C(��^X�p�>�	7���'L�e��ﵘ˂k��\� ��8qAp��4#Q{2W�t�i��g��i��2j�p�����E%39����xdQ�U�ą�ŊR	]z�(G6f�Shu�`�W|@������E��+��Ἷ�S�0�����F_���J�����̏�I��ꌻd��z�7�e�攏� q���1D��y;-�;�/���	���Ѳ�`	$J��T��DDR ����s������]���N^s�{�b��\Q{b��iݨ���+� �v
�((ϡ2�t.o��௄Oẘ�~�F��<٬�#<"o�-��������U�6�(��B�^�V�%wi��&��|����e�h���D7��jr<y+�O^V�_4��s�ZD�m����x�JH�K�6��l��"�O��|�����I����5	�����ڕ\Wc!�ϼ'�^F:�<�J�l�����yaR!odL�>�i��[�vb�_f Q*��nt5�m����O�E2��RIxZpI��h��� �N-P���J4˔A���o~��~��8E���k�
-�3�$on*�Km+�+`�t4�o͝�6���%��5��T�"w`"���}�����c����o1�0�HP���W���>V���V��P?�]�����ɹMS~2�";#1�QB����YHJ�z�1�� 3#S�#��-Q�����n�$/����Y��3���;^I6��!n&cp��G��}8Ֆ��!)i�V��"Zȼ��23�Ywf���ܖN�t��Ɩ�ް9V�#�=���(���G����<���Ap��aW�p�%xPE�ҫ֨�.Į7 ��@F>,Iߡ�~��.YFIl�]�P������#�^��U��m��8
��<��5��$�*�co.5H,�L&��Q���-	[" ��eȡ�K�@�!�	�T��3���9dh8L�۱��iH8��0Ϸ�)C�����hNսFeG��.\x�h�t�Op	��x����~5�f�ޙ�wl���6���y?yaDdzM��QH��Ⱥh�ߪgc�K�1V��|2�W��̸ �}œL�,���+�ON]=�XA��`�˗Ry̇,���^XM;ܣ�D~���ԢP�Nw��J�DFn��s�^[�N}ؕ>��r�4�9:��]�`��E=Tr���׺ҟ�'n�54՜�
2�i"x�LC�ae��5B�#� �E.���#��Ŝ����w������Lq��}�y� �z3��]�Ix���|����u�U�/p?sE��i糳��t6�B��0W~��
a�e�
C��_����D��&�M#Ը�]l~_aஔ��77��I��vL&z�U�s����I�����jP�E_X27T�*1��o�M���og=�P�)�)�o�Nv10��|)fCZ,g�H3�������9a��}G�wG2<z��i��ۻe�b�]%�w�ד������u�|� s���WfИB鯿R�����eMqu���@� �Z�h�yy^;�%;r$�l���[N~�d��yO{ۮX��.��{�2I�<�F8��Ck/�d���/q&��F����&�_�<ӹ�s�޺<Z1�����0��)fbWd�?��*��8?��VѬ<���=�h��M}���q����:-�8K���DZ��Q��X�ם�ߐFo{SU��!�l�X�_�G�z���3�/�Zd3����C1w	G���h�u��A��;�� &�*U�G ��]Y&�xd�6Q�X���o�a�w+,�L�*�ѣ��B�ɹ�V�b𽻘�L���[�۟Mb�j	؝��w8n\�p�*,#��%,�"��Eq��WR9���{�᠅ћ�Ns�2���aI����MV�b@�U����R&�>m}���LEPT�,P̐;� ���3F�i��B��ZF�j��܌Ҥ�C���gh�+���d����M����Ni���A� �
w<�;�N�n�b�26!�\V����pHPB����ﾏ\��|;��cԎ��g�������D�&FfVf
�(GN��[ڠ��/{��J.�_	iZ�Os�Ð��5|�]��!s��ʓ�=,VOH�;0���u��݆:L��&P��Fv��_^a��V9zr"�f�^n��&�ҩ��"G[o�~2�}��������R�����]\'L��KN��/��9��
Yc+�T�,�~gO?����R4���e��F����*��������f1�$�^ۣ��V�3(�	�c���\o�R�7?r� O�L�D>^d�8����Wq�sp� ��K*-
O�:�qs'�C�D��mLe��H��Ⱥ0~��O�����̑)I�����r��v����+ ?}}��m���/�BO����Pp��]W{W"�K�a��갮z����|Չ2̴z��1{��-?�Q��vբ���1Ix�E��]��ɿ��G�R6J�۱�d�9�%t,��aO	[���qUeN��OT�=!g� cye�,��3
ѳ��ߦODGS<H��l?.�֘c.���ZjL[����0��T1p��i9idK��
���$����\8�WU�G�}�Hl�:����~%�=qc[��#-�Ϙ,����c'� qȟX������Y����V
p+�H�$ː�U��wv�.PW=�#/:��vm�?�aN�W�!ђ �������)+�eW����y�bE�^ �>�o�#�^:����z����I᭙�:��U��C��?ǔ�����<1Ƙ�7�!lu��4��s����JWmӑ�;ĕ{Y؎%V|�R��n/�s��q@-�kd:��7)�S�v��[�� �x;	8�}�4�r��В;�\���aX���[����FL�Bђ�o�邶�x����&�!����U�xiμ��&�fn�g]/$g
(�thZ�{�lE�j|���Lߍ�.,y] "�H�ŉ�D5)^��U'ܷ����� �����1�c��9^,�C�n��l2)��V94Z�-�t�)i��+�u������ظ^t�(U����n)ˢ���~�16��:h��.&FԒ{����j�}�|�N�Փ�X4�=�T�]מ6�R�{�ID�.V褥��vxM!�z:\1��e#1���{Ý�JB%Kq"O�1���H��,'¬��Pb�V˞�~<O������e=����R��d,?��7,{���
{��������72S^���3m�A��������Y '�z1`�)�bI��u��1_y�w'�ΐ�Ž!��z���֏�4@S����<��#�p;��P��ݪ�f��m���.o�����DP�`
�,��(7ĸ	5����ģI�Αo]>/9,5��2�ӂg[�֖j���$��UZGJ2��7�x�0�H��J�� �����y�3o�1S ��gC�{�7���P��K*\����y�կ��H�h1�����>�U{Ykx�o�n����%i6/��i���*`r�8Mx,4އ��mP�q`�ϩ�f��n��q�����8z�g�(�=�"#���L�N�;ŅL!h�����9��N�/!�]LU�t�c�I��!�ύ�U��sZ��#
���?��LA��Uf6�C�u�z��O��&�-��Z��bs~]�}:C�N�N�*����"S��nfb̐8(��d�ˋ��Cz��sƿ�#߷U�n:<nG�"��(�<U��� �*�/C�����Y�M�Ⱦ�%�g��}��d������p`����X#���wW�&�v�u�gv��v�-G[r����!�
q�z����r�<���H���f�+�7F'�-S�9"�n��ԧ�葋%.쿵���6ĭFp
��Ɍ8Ay�Hi ������z��\m�cO����rk��?��q?ipª3�h��h���4�j �W ;��kA� �vo�7��ywm���'ᅈD�a�A��1�&��	W�����cΧ���RuJ!^R)lM[�Jd���p��^�upr)ïN�e)����2H�	Jn�;�?��V��:S���&6�Q�СzՄ�['fH���@:���5���Z9�N˝v�@�7�F����7�4jr':��[��Zj��\���L�Z	u'�)9���N�%>�:�R7ų���	�3u"��6ݖ��y�ӢHD�땆��[���!Ւ�Ŵ�ވ\/ƻZ�i�r��SM�\|ݻ\�Q1�*:��	���.r��<�-�g�!9aI�GE${1j]�Jl%��m§E�Z�p�]~��T������ɛ�x����/mk�s�?e$���i��� �Y]�OHZI-,K�Q�ci*gS �(�\<��.�',��m3b��X�P_�jb+�-��>����C@|U��l����4
@��KjI���揂cL�� ���2�o�igT/*�N���3����"a�c"�5����Il�/���d�Y��pS
��}��[���a�k�=g�.�N=�����v �f#��nL���������9Ez�An@�X���g)7���i�ãݗG�D����r��U�z<P��=r��S�`>ȱv��}��0�9��+�?�L�#���=�x�T���E�x�nO��#/$d��Ӕ��g�������{��}~�|>â���S�(z��J�;yȓ]C�&B�D�P։��B��!�y���<oYا�6�u�lJ�18mq8ߪ0�y<�%��an��Xjwڗd�zQ9�ƱY�'6 ��A��N�ܷ-,2O�{�P��[+#��Bm��䉠�����$��������&���{��Y)Z�&p�lCA-A�!��V�%r��0���ce.$iB�3:'t��I� E�a�d��lܨ3���=N�	9 C���{τ�!#\����PA=\�	��z���	������[z��{6wz%��C�������}߉��Y��kD	����[r��(��slxv~�ATD�"Y���P�:��r�Ȥɇ�9�:�˥mY��",�:���/�$[�\N�s�g�T+I���u�+2��do�R�o���H����2�|����L��6�B��O<��g�8�����]O�������:5G�~X�Gw"Vw{e!�XbK�^R�x-72CpjVBV�o�,a0	���"|��G���b�z}&�{q= 
6�[��I$�gs�𢚜L QJ�Ea�)#�J$m`�����L���P&��eV�e�<2i��7�i��h�u�cF�Rr�Iü�<�����R�	C+���"�_I�	��)Ǩ�8��Qۚ�ף�!�C����Q��������3sm)�&>�oz8����!�9`�Vy"΀J�������C54?C����݀�}��{�Yl%zf�� �.���ӆ�5γ�Ok,'*L�nGsM�Z��y�k�<��%�2R�����ĥ�vIq0�n%ȭl3I*pjLL19e>,g��i�G�H�G	쪜ZՎޫ�.� T�N!��N��T&���G8-�-_޾��9i��`�2��ل��\��>Ez���t���4�l��5��2#�m� �X�v�	g�	9 ��o��G�Z���+���4+�V
J��5MRK�ٺ�~�.Cۀ7��2q���W`I@݈�]@���jě\����j�h�t��U��h�Ş���&b�j󩓒�]�N����(����a�q&蒺�-�ĭ�W!tq�J\�^݄(�m��m�{�.��@�#�/�NW����+Ov%j��\Y�%�ɯ���<��wX�S��2T(4>��X�d(b��++[�5e���JXu*�wTɩ��cJ�P������޳٫Җ�j��!�j/p����I��w����Q�Vs���k/7؋DrI�e�soC�����2�O�N��xOg��o�X����א_��@���/0�X��e	�y�����@Y^4c���@�>��us��G��{:��v'�����w@ɀ6�h�.~�ܘw0���0G��������Z�|,�!c�ޣL�Â�-��bq�5e�z�EE'�j��)S{��T�&kB�z4Y��[�{\H$ɣzN�r\�^�#�^ؿ>��C2k�c�Y��ؑt[���1�^h�Nu�s����][g���q}_�v���@���=���CFf�b�P������[��������]x!�c�������F��oXzd|���#o����yl���Y�ָ����`�tLԹ�ip.(q�Z7��������e|1�0�7���,\�̱>O����m�ΎX�.���.��G���~��Fn����;O�֥^k�Zee�"��:@���+�����a�eH�u����^�Y��ۯ4�5����,~�;EL� ;�c�a4e+�6�p�Y���/���Ḁ1�}{k�6����;�TW����!9,��$��'�'RUb���P����`n@�Ú�	�1�50�R��PЁ%�8�p�"�1ڮVv^�UF��W�6b��n
�>���ـ8k��l_���-����OK��P�_��������s�"�ڣ`�O��Y�?&7�m�J�_Bl2Ύ�C�C���M��w&<C����p�F�9V��/���v���c�x��_��,`ֶ��i_�fO[���~���_��Tuith*DXW�.o�J�+Y��
�L�S��l �=&��etwX�����T�o4�1b�]ZHnW�?��̏m�m�(�L�#[�q���2���|Km�~I�n� gD��r#S�6���V�;��aNC1�}]x��A��h�c5�ο����5�1��fL�-��J��ن�x��Y�7�����e���o�e���S���Ux;����D�5��,��`��]�V��׺�!���q���V���P�7�����"��7Wy�t}O�����18��i��EZ@��)��#.7�V*u7u�YѢX�QI�ϑ���Ҽі��2��1z��W�,z�v�H��c�J��]UW��٥�ܑq3î2��'���Y���3Y��c\�?���/���\+;�|�h�n�m}�=����U�Ɂ_�)�7b[C\�BQL!�?#C94�I��&�����	y첞:N,f���m���.(+.� 'e��'��Z�tLb����5��2DDF� r?�P��'Y5�\��n�BI�Ph;�mM�@^�����
�j+T�r�QR7�����l�wXPK������{�.�a�|\z�YE�,���M��.ǁp~9ز8�q��i�U�U 'S�ihy�7��2��}j��f��7� #�u�<�k��U�8*��&;_{������R=�*�
k"�=���҉�_�k���Cp��j9"{����z�|{��}�:FMS �r*�,7�.��uQuߺ�ȑU�)C)���V��Y��y��7�u�u7���QZ]{��`��� ��!T�e'5(`]���#� ��&f�L�͓��v���'�Y�5+���D��� ��;rc��]s3��9Pī.��gI�� ���ߔ~�9��g��ן�L�h�����]L@�E�{�k�+�b�Ꚑ���OD�X%?a��n�d���� ��w�����jB�8u�^����,��b�7/y��kc�/���u�P�d�3ԽÃGd]�����E+������8~��f�v�o��R=�'B��x��/��7�A��!��`�(^������ N�K�J_�T��d��� h����OIAv2']h�����h
�|��|o���"U�\t]��fZǱ
\t��$���L5Q ̋�o�Y���R��H�跺��h�1�@|&5��8Rp�k��{����:&q-o��wK?������"�i�1A�︆��}8W�'��'W��ʶe�#}� �|��E�v�,*�b�_!G��AN�1�7!HB{�uB�5Vn��:��1	4��@��S*2J�d����3��65�̊��R�GC��{��q@�e���]��V#���aw�_�0����C�j�U��W��M�����'�#'����Q�p�.!j��X5�������q��ԛ�yS��U�!�4 �!>Gm��F�<|��t8�dҺ}8K>g��|/� ~�nM3y^��D�o:8�����?|����H���7Ӊq�Ӝ��=p��[_W�:�#��Y���$v����\�.�w���#0pk��%�a$�j���j)��{(IPV����Qا���_��8;��˲���|<���@�o�۸0�9�����Ґ����&*���B���6�4Z���b��^�x����f����NG�;i�, �HqM�qб_��f�k|)N�	��&*g����v��8a w��<�f��Wp��� �;aŦ�s#m��Ԑ�b��͠Q���p~y�oJy�ԩ��<�g��+^���!��ܒSR>��oIPɫ]�e��۹��%��?�5�D6�����Gi?��*���\���b��<.�@�%�����!Q[*mIr�����`���}��L(E�d�,��^R@K%4q�՟��7�Ef���� V�(G���_]�P�ڌNsn�8?(Cr��|Ĥ��G�pj�nf|�^��J�������͋�:���%lj�-��f��b��
M���Ix��e �����,ͅJkP����:L�(l�xk���;R���,��z�։G�#�D'�j��#@��b"�@�����Z/y�3['@,!Fo����pP0��)X�`��L� �p�R1��Ggυn-��"V��R�4��m�%'Ŧ�����S����Ѳr���(ȬC�Cbp'M��M�
���B5n^{Ǎ���N��k�+�,	�5�Ц4��:{��P���Ls�K��ǅҰ�T��k�
g�g'�X�B������Q���V .�OY�w�5�\=\�>3c!�����0�b5�0� ́���N����V�5��}�� {��kz�� at���8�i/PԸ.�.����ch�(����\��:����)�O�Sr�DE?��'����U�'��	��"b��:9U԰����#|���],�=����.���R���#����nE�)HQ�Y(�@L���|��z=�o���Wv����y/Z�~<l=p�Ff�J�g j5�ԍD�t�TQ(1�:)B�����t���������jH��E�>q{O!:ڳ��Y��s���V��E�u׽��(���-��w�q��:
��1�/�l5�7ҫ�`��͗!�y|"�z��c����|�E8`v%� ��´��^Ie���e<�yF8	�|v�ʃ�,���[�u��Uc�$9."�<���/� �<e3�*.Jp��ȸ:�C�G�HS_�ybkk5F�u�u/�/�J��w�h�~Kr2FC�4��L"7��Π��텢�!�r�����n�Ā��J����u�jy���/�5��zg)ԥ\a����x!��_��8p��V��z�6h�g��Y�.IT��hA��[��2�S7��x�+wt����N��mY�Z��^H�����R�ޏzd`-�a���r2�Đ&4�EFD���<'�7P/��B�M�BZS�P*�	1�}��O�%��2��/r�S�בDV���8#['�n��y�4$�m�0����õ^B�.�O�	��&���)׆i��u��|jg�^"�R#P�q�����1ܐh��O_���k���!)���s\��1�
7Ԭ8 N8F���Z+ˆ�YS�k�[�vOD~t%��ܟ�m�N>/"i�Rr���F��r��X��S���<��A�Ĵ21�$����T���St�+1E����gZ_v���J�Kg�|��}��[�_<�´���@j�\��AtEYr�8�壘��wPN���?k ��k�"��T��3�y��(x"Zփ6'G�J�|Sɘ������H�,�j�b'������1w~�j��������qs�؜|��������� �1)u�Y��P�3=�do#r��!p��@C3�W�~�P�}�
;`�3,C��FS%2]�<���&�����L�q�&;�=���4N��Q+�tY�0�9���Y1��k;7�o�7�ڿ�Uu��xi��`���&�5嵅�E������*j7w<}�cO����7D������-�7K��+=&�<�~⪄�巢����0� .�g��
l��{����cF�W}R%�#�� ��ж�Op�M.�T\�pL�R�&��׵�(R�.�7���@�Q��1��Y�^�Y���?�&u_��毑�[b�N�/�8:���^��.�sa��N�*�.��e"��@�S,�#I�RncuD1Q�0�rȮ��D�r�t0Y�Y�?spm����9YyV/3~k�et�#�rb� �G������΋?a	�~�1�-&�\��h�U%������ti1nw��C=ĺ@
i��<4$�e��ݯ��^hӽ�Ȧ�cc�a)�>Y;���U
���pBC,�Yz����G��2��4���H���?s��t�o5f
�+ {;�G�|���A%w�s�.��-�s�n��b6]RӨ�"q�����!s?��C)0�2�*�L:��J���
ͱr���o�������E7�(bp3G���⚞�Q4�4�����4j@���� �����C����U��8v�TJ�4�5˥���!�E��{nDg}�3��A&�O�]��L.H<����DtN�[H�27O����EU��\<����ǉy���T�-����M�4��AyE3�XD��t�-f@�G�_�(���������4�C}������s"0ױ����.�;�Ǵ����e��R�Y.��T� 3����a�)���ɌE0H+�|W������ۃ���C��[�4���@���j��	Ix(\�Z_(���o��UЦ)@�LCkRKA<�N��7�$���w�)�l�D���:���	1��*ygfzԒ���SV_�D܅��(���>&!�Qދ+F�zQ��x�4�0��'�?ń�`����ilkƘB�8'���"�`�՞.6�֬�����Ri�,�)Z8��1�An����4�8�f���\y`�	����_I��¹ܚ�kN�M�A0��f
�e�XfJ�k`x$�P>f܊����0���Ц�{M�?!&���&��=#y���e>���&�m�(]($���:6
�4@z�OL���.�����D��nV�ٰn�*�7(�M`^���C�!�{1��vU�*�����A*�y��K�
�я3��i�u.�p����6�c'�q3��Y��K�ݽ���k��ZwE�3��'�T4i�{��]�8��;�	����~��拑�{$�����C<�p,�\o�ᩒs-#���q�I�ҝYN���S8,w{X��v�+����>�׽�XE$�:�;�A����W���ؤ�?S�7WG[QR��.w3(�N�G����E蘸��M�sH�,�A+ppM'0���yKC�k�9:�	~���{_�]����!̂2��Ԃ��ؘ.�7+oi����>���단�|θ��v���1�EghC����5�l�nn�[xf��	�&�v���8�eF�[���/�c�ʄB��=2$�D����8�@%m��.:�O;�����O��.�8M���+vED�WXT���:���r݅�Cpf��^-���a.��0�(m`��M;�*�<G{M6[�� �^^?Y(0�.$ab���D<79��b����TD7P�;Ee�o���o����s�&f����!}��F�BL ģ�-{u�Oi�ᠳ�ۭcYP��86ׁJ���G'��:�Yq$/E]�O��i�pz�j�ֈ+>ĺ�f�.l�Y<��C5�^���S��Q���B�j'�E���l�xLWZ�"�@ ��T�����3�ϡ�
p�&���k���{!��fɖ�>g�>P6�SK>x*��Qؓ땺_�l�\Oڧ�?����KA~�#4�������\J�q�@
1�#>�7d�(���b����ն'`8�{L����㩋i��j�yN�O��R����Mm��}U��q�_�Pײ��A',���ܵ��J}<�r�[�K� B
��f6~]|T[�G�/����~��tF�q�#�ӽ�TU�|���X���+��A$��;���G}yY�:u�
�VH��e�$�]V\����Q������d�]�dn%-t��ܑ��W��	�L�3}��+֐�ހ�-����ɎM$m�g�P?��T��������?�1PB�(�3m�3�o3�#�.y5{<�Gb�!�n@����9ݍ��x��co�1���/FQ�8��5�c�s�<�W�=�E��,7]��-;�v^XHd�Z|����hcM��h��:__��{)+I'��� m}J3��9d'��E9�q�T�/�+�����x��G���]��H�y�b��������/�gEҼ�,�3p��=YS�7�i��R8 E�ڶ� �z�O�z�JU�z-'mVw�,��C������B,��Eq#������_>#�t�MȽ-�Hʯ���tj�[� ;��]��x������z��%b�ƀQ���������~��&��[��҄&�k4���D�'�p�<~�C��9���?�8�%$���$�zNP��^�0;��T	LT,D��O����}��AѼ[�톞�x�T�P&�Q�j>w+?2ZE��}�bM�/������_J��Mτׇļ3U��F�/ʼs�U�XR� :qW�����ʞ�`�H�>���Qea����Vc��� �<ʝ����B�D��H��NZ;�Ѽq���(�aY�#������H\�;s~��8��}�*�z'f]��tڵ|<50�D�R����i���A�õP_��-�ШAԶ̎�?'�j���VCA朡?����"l� ���7�+�N����E�}��_�'D��\���cbx8|}B:�h.X�׵�E�H��a�Tm��չ
�Z~aό_�ǎ���}PQ�L-���~�`<�a�2	w3Z��O&��[���+q���f��r�6r3���(=�`?x���˂��f��2���7��
��L�7�P�g|8�Ta�ky�)�ZG�l4+�*�"�  jekf@ߚ{8���T�,T>��.�'�.�,��WMA�I�gTSv-'��͸3���x�~�e�zb�P��P��������i2�?�^W��"���g���|����P�_���ԥ�O���U2���e�CDN4�\�Q!�]�> �*'�~͖��{f�o���0�3r$:������d�P��+Aq.���[�k���}�Z�����g;#�WGF�����+b�!dz�8�N�`�a�,�ŉ�"�+�A��KJ�W���Id�L<6;T�<��΍(	���dj���e��J��=f��p5��%��8��D�
|�N�9	S�-!�f��n���*�%5G���E��9	�T�p<���Me	�.*�}��w��T���y��ʌ�=^Pl�h�.�Pg��̀D��ߴ Wgp^%^j�+e��Fɏ��څ��]4"�m��o�b�����~�TLC����
�a��w����Gr��Ģ��Y|�m�.k�dB݆V��*ͣPD�@F!{p���B{̇�<�r��n�B.nMQ ��&.t�!��j����)�U��*u�@z���g�L�N���w+Qt��^0�Ę�L[���p�����ͪ�	�/�Z�����'�|tA���U9��x| ��f��>,�WZ��bR��Ռ]���Y�W�$M;���2`�At�G��� 4}���d�j��q40o�I,��헗;�W�U���B��p״���b�gT��v%�C �}�&qyȜ�5��?�;5��R(v<���]�:
��7_��6�jP���*`��^y�<z�@2������L�P�e���Hp�SZ�v�2ע�Lf���KwQw���^�]l�MVR��#����{x?��$
�v�}}��G���/�]�4h��WT
s�a�P�0hg�����.X�C���Y�W/�z����6�Pq3N��Y��O��h!~�4K�Ȫ�����������&��ELE�x�)`�����"��҆���z�}AL��}O	8�Mis�"�	8w.<�����#��	C;g��u�E��;�e9})�Α!�`���5�t�"B�lԈ_��o��T���0r�5��Y#&(E��Y �/] u�P��O	z���S��϶A;d�n���S�Ń���ݛ�uh�F�?p�������7z��U��1t�s�ֿ������u�19��#O�[��ux�����G}ɰ��:P ����L�ũ��?ghn<�Q���ER�K)�n�k�.�����@��O>݇G���E;�kP���m�H#���v��1,�Ӧ���~�]Ggi�	hGQ}��i�ZV��B1����Y����˞Cʦ�lE�	�;���j�T7��I{U�iw9���6�|:\#���̅ '�G4�'A4Sc����5��p�Y{��C��D�<�b�*H���_R��ς4L����U�[��9w"�8^��r��w����K�h�^�s�VM?-���L7~i�P�-���ߨSs[iY����>&O�G/p� �5rzӿ��i�J�[؋��b?���C����������ϩ��<���2Ԋo�%�&��'�0%f����Yq�D�{�g�?�_i �7
B�!~ocoe����(�3H�%�ύy�)�,�4⬄�V��(\���5Xݞ�狗$9�7D�&с�� �]5,u�%�O�p�p�ׅ����*���٭���=Z\���L�������.�j9��"(,�X4:p��2&ϫ9G�;=��Ԧ��z0�9�9�ʮ�<3=� 9�;��صK���D~+�hz>bK�u"�!@�;8O �	V�D�b�T��3�%�x�*����/RK����sQC1&:[��=j)�lr����M��G��LcQ���,�����[��Bl$�����u�B���,c����o���Q5�	)%����{�%�&���"@��������ڜHb~���5̈X��Sv��1�����=~ �Q�se�׺�wF��4�3��eR��o�k�����Ok;;A�gc��V�����ޤ���ެ�˖?��JQ`%��V�G�z0�D��{L��h�8FU�>�_�����i����������[�od��8J�V��d�u�_.��Gt�9C��d�ar����X_lGI4C�� �ƹ)�����vF7�0B�W���sWV�l��Ԛ؝�n�y�=xk3�Oz����ۊk6����������˱	�ఘ�N���e!a��yE��<-�-?�g��D��8��-���A���oeG�����ꎽ�t���{�ĜA"9d�C4��8�D��S�͕�"j�-nUewz�*���D�@=K��t�޸�Z۰�arm\eg��t�e��p�_�,?P\K~?�	�s y�S5����)\]�-O�B>h��Vh ���t0Hn^�*A��+{������-�rv�ߵp8F�dR����[O�'���O:���*F��8+gK~Q>B82*M�0�b�U�Lg��ݳ���%�6Ѭ�/�-����\���!���L]9���>�S�m@ɳ��":�m<; ͹ГRb}2���PW@����a<6.n� q=�-A ��_�|,���bqK�xؔHl·�a��Ƭ�/zt��B���E����%�U.g�)5�yM5K���i��1lmB��}��������S����_!��a��K�z�>I<B}�j't&����v�C�ج�l��f%F���+^C��t뙗��՝�T 3E'
�}�b�9{�>�����e��׽�?�RN�}]�H[�CV.~C׬V�T��uWΜbl���x/l����$��-Zh��.6G�y��D����O)����D�l?�_a�|�H󞄽b��W�=�D*aM���=�M�_��!�q'�L��iWSd�{��#��8�!��L5���v���Yl�9����9�[T��Q�A����P��pORh��o�T�KO\d�G��(Z��y�Gq9\�%"$��5�0�G<�GL���6ԂA}kΙ`[���׼Bo��%���[��5D���L*�L�aӔ����gχ!�l�gx1���l졋Ӑ�dL��$}1���!�G��m����nJ�W�P�gTd���0z��;�n��m*F�蘧�9b�,ǹ�9�*�#5��d��1�Y+��#�\�?q��Su�ٻ���n��o�ws�����/�m�O�@���xu�T։����;���l���F�u�C1�Scv|W�r�Q�!C<�Ɠr!άD���K�Q�: �*Y�L@��~��69����9����6ĝ�?m��e��)�W%�&�V��4�~d��BP����$�1�¢���}U�tp��\~�ogB������=mv����m��La� �{����ir�%O���ǃ^�':{��#ƢU�=(��5ݳYZ4��b�܁�q�O��h��=�S���h^S�'^�K�n)�|����Y��l̸K��߯s�Iu��^bd���-s�Sl1�m�X�Ad'�Δ�S9ȾԳV���	"�-Z Ha���������ļ�>k��ƧC���L�
�&�JPsF�:�fM�8��T[�ĤQ�<��߱�?�=�l�~�|��}�~��\�z�{�-���}��9���c,ٟ,��Sm�R�,����H �J��|\�q[���j�؛����K�F�'�]����&��@��q6#%r?<�$w@~3Q�yY rZ�GVb��b�Ɵ�=}Ջ�>N.���w7r9�l�~n��}خ>g~���-��(�'g��{ԧ�[.r����V#p�xDnNl�`�*[�ZWR3K�Q����;���TB�LI&�-��yn�*A�yy�����N���0���$�<�N`\�d+�e	 ���\~IbA�D�r���ӭeF����w��^ec]�3@��R�A�#E�[AL�U�C9�N�Z���b�ud��M<��9�D�n�o��9�Ku4o��	B�e+���}lPݤ�4����=Y8�g��*ff���j��VÌk� 
q�7��[�j	������[��P�lȸ��'#_���y�p���Нv��d`f"�6hTC��Y.'q�D���ć��^%v.��z>ҵ�AVk�A\��Jf�&g�d?x���Jj)9��\�����Y�'Z�Bx/�Y�xZusD�T�j�潩�C��n���S�\��c��ۋ�ph(�`Ѓ��ac�,�3S�"^�{w�I����WX?h<Vl{���n,�./2qn��9�t��
�e#�G��{j��

�*P��o�G�+��:��d�ꑫ��9QxgLod�g�,�)1�U�� �LWr:�_ɝ�c�#�rD�0 `���S��j����&q'�;�l���V�ρ썬c�!s[[iG���]t,�:�9��K
K��h�辑���Bꌒ�c�Ӛ�5�Q��Ü^��o��kMς����̔Tۘ+�3�v��^��M8|Q($?a�©�	}�}z�<���?FY� ����Ԁ.#��j���<�U1�o�N��g���D-bT���oV?��
��w�����;���a����̥�LM9%̢q�x�n�V�N7 ���UӨI;�fX����ip����!� F��|ك��5
%qt��xӂ5�:Su��}�dU.wOE����5�1F#_�$���Kk�7
�ڒ{�ȉ�L��U~E� �:��9J�q_��|�1��߁E���]��	�X���7�}����%�����;��4C��~:?X��5&R/iM7�R�m�Z; j-3V�����Mm��k���^����b
�F���9���й��qfZ������uг];I���ԲJ�:������,�J\�#E˞t���(D��{������Nk�IdryY�멉��p=��Q�T��#"JSX���$��y5Ө��{&M���7;^�m���T(��k��v�����U7Ρj��c�`�����gئsW1����(���;Y1�� `޺@���*�۬H:����sq��^�ɱ������4��3F��H�OFٗ&�M����ؚ���cC�M4�f	-$�򉿒�z������-����yw���d��E��N�5�S'JC�[��z�x6�w1�j������֕eބ�^#���Hj�����B>��4��j݈~��,�����|���Ȏ.��K� ,^�M�^ȫ�C��ΧDܷ��Wȸė!�ě���j�rqerD��ُ�Q=��
�ܘj�@T�B�Lml�0�������G��͸sV�MR� lMe3�{�r������a=6Ǥ_�!�E�'oF��^;�Q+~�?���r.��t�����'������a�'������s̕��-�Ŕ��y�DXHz[��OZT�i?ku_XP��:���{2t��u�k�[��k��W�n���ي�����^O���L�]�'EߙZ�U��7Mh�Y Îv=/��ӓM��Xv��Z��҂U��Z[�nU�q��eC��e;�E��1��G�_�i�|��S ���<�����G��X^3� ڛ
�z��k���	���eL][Vd�����^��_�����(lj�?���oɿ��y�퇦��D0+��#e2�J��ʻup���� ��q	����$��t\0>k���%�$�"r�5U�n��׺o����z���y�s�s�O�F�cd	(�i$q9�Gd������/z����8�����i��1�*2 ��A	F4n�_+l@�?[T;@/zT��Yc�y\��r9��d%\v�����᎗l��s�+e6�h��!�P|��Խc�����'�G�R�_}�4�d�@{���V���z�#��([kҸ�Կ�U��g8�c���ԍ?�5A���c���u��W��㤨m����i�U�[��W�G*Vdu%��8Smߺ�*!�gg���b�k��VJ�@"]�cRT*�ٿٳ���'�3�/���<�j��g!+���њ�`Ȼ�EQ�_�j"�<Ђ\(���v�o�����R��n�G*𑞻�V.���>s�R/l6����5:��Z��''U�~�¶ώ8 ���:s�F?3�F�=��
�B&f���S�5\���r��A1v�� (ÅfA�H�utp�Wp���\���D� ��i��L��S��tS���N���"a8��b��y�Y�/J�S}'���Mq������H�8�.1?�m�}��<!���p���΍;�vJ��� 1��{���"�I�q:��h�<S��g)�a�������1�� �I/R}s[Ww�Fd�cc".T6'Ɵ7��s$ 5S
�N��I��w���ZF�f�>�
2�=��M�_�Z�ڎ(�w�a��(�2K:�H��lq%��U 6*Y�Kز,����L�C=h�M��#}�!�pJ~�W��s�AQ�;�;A����Cd=h��y��WW0؉^,���x��V�'�b\]V�	�!�������[�%����p�3�M<?i�z5Aa�ç)��3thP�Z��B���R���:��Ѣ�o�r��[�Y|�\'l������!����$�֐��]t������d!��S�־��#8\�L�-n[�ecx�����Y�j��߾k6,O�~��ד�(5�1��d!?�^�`Μ��B��!'��pͱ����I�2I�)�>�l^�R�8;�v�8?��:0N�W�j1[D��ІWk1$"[V=�h����J�A7�<g;_>�������#ߋ�r���x�}���[��ݺy��53�	rf�sk��7�pm,?g�����c�N?K��Ǫ�uD�ݕ�!�T3R��$Dk�G]��l1�x��>#\�r������{�(���{Gp˳�/M���R�0B�{ȡ*3�/�Ԑ@��_+c�0���Pƭy��8^ZΓ��L2)�ϊ��a��ɛ��]"�$l�ʋI2ј���H�)�>��:�Ph�l�N������~@�?Zn��)Dv�:bp+>�8ִ���|D)����q{m����q�!Ρ�i���L0��B�hJ UBVE]��!FE��I����4k���׏)EH�\���`�2j}�u��>���e0R>b�~��y�F���/G�aS.:�-V;�]��G��fC+/��f�ܤ�gS����40�;�/�c�u�%����K�����+��������]sں
����Є�]u!Jg|=�����3���9�QB!��a��Sv�=��P�>��S�y���$�[�������=3dp$��3��y-^Qh��v�BB(EaR���a�>*�	��\�(�M�s ���+��;��=��+umN�{m=-�<�&�a%�����P5�.I��=;�(���j�ԛz��0`�E�%�&nI�����䦨9)G�(���ͬ��h����j�� ��'�O6�;�[����C_f_�i�\�3�P%
\�|�p���=jw�\C�0�,��QZ�>sW+����O�	�p�$p�L�ማ���Ul&��]}>D����l��Y"u�ɞ�k�iH�=�Y�!�Y�U0r�x�P��Ɛ���>������C��`�3��8[ me��t��d�O%J�������S'�#c-�����r)�t�-�b��9��Yd��ӄ�qj����XZ}�9Dpb��)NoB�����ݟ!W�rn���6/�A!�)�Ơ:����	�G��B�zi���Nz�\��{�/�wފ�v?6�h[��0	��`����v^�{�n�E�'�eU/�*w�[�)5�^'�'����쯡���w�r`�ެ�K��-林��m="���g���1/�׆�Z<Z$~U��FH ��`��%0�)���ʑ����L��	W��	�]��'�X��b��Z���`��[���M�֬x�T�����������j0l������d��=Y�Q��B���6�X�#U}��wb@>�#�c]�[��Ç�<��>O����F,mO�AS���?c�)���3�ҭĂ���4��P��(��~"�C�&���QX~�3m5�p�ժ*��i�XTz����ñ���#:�n�#/1�m}��y5���t�X��qN2��Y%�`��4���5�_fI��#5��lÙ�L(�v�ec0 2A����H�!$1U�;Z���3\� E��a�v�T�<X�.���Ji����hˋ(���	�m�1~��[�|��4��R��,�g>�q�Y���oo3��_�\0*O��]�%� ��=���_ќ�=�N"�� ���^��3�D {�`�����XYA�|ᖾ�̴y*�*����Sz?��N�|��%ȟ���tÐb?L8!ӗ\O:h1�7��Ǥ�`�Y䢶,vj6�쇬a��H�+�@_e6�WД�Kv��
T�h�J��~9s��,ŝi[z��R"(��3m����������I�`mo��r�	�����#eFZx�x��m�� ���<B7��x5�/��H:�A�k�ӖS�KK�Os��ӨC�Iϻ9~B�{7.�&�<x��h�r�'�pLb?�����џ�=�z�2��4-?@"�IJ�� u�"�!�6�,䉗���z4_��y<|�lޒ�yM!��ց�GD���$���+�j9�c�x�.�l�ּ������|Qbǟ1��,3�O�ps��{vf:���a��!���>���J{�;��� db��z���.d���j֫/ӠW�a�ݯ����\,��B�1�$�?Dc�`��h�/�nY��&B)�4����Q���Ne��94T�=�~�ZGx4��~>�������!�TE�ąNcJ�j�C*b�v��Y/����e�� ����Ѽ|��8�N���h±��n�pp�X��N2�";&�e��\�B�K���8��Tv)�x�X���^߄�X �L����M��NS��!#_�jZN�c�K^ cd��W�V_cc�yޔ�=R�6�4$�*�p��s�u`щ^�I������d�۾֛zE�B�C@�1�q?��mr�V�J�q��X<Y����;apx�.3깵���c,K�q��s�N����?s*ѫa����^c�&lQ�ң�����M��U��Ci(� BT�ƙH�st��I?{q9�i�����<� �Ξb&�xx�=N��$����ԃ[S�+��ʆ6���DK)*G@�����Mq��p`�,�7�n�]%Y0�3�#�<J�1�Ǔ�\0��@��Lւݺyx,hp ң'��n�K��7��ʓ�P�/��������M�V?!ٿy���݈>�K�:��7��t㚬2	ˏ*������L��Vk���l~��H��q�x�5 9%v�o�l���]��~�@,���������+�muf�'�*UQ�iL�l��XZ�rG����=\�d�Wb<=J�G;z_r�P��z=�� �u�B�ګ��n��_ԙ%��lI�H+F��RZ�>;���R8x��+S�l[*�|(���`�E]ڦI��v��2�m�V�:�P��v��/uv�� }�6��d�1�M�&B�L�$�^��Y�nw�;M5�LTG�X�Ohz������ �j�4ArnT���k���$��fĔl��G|�P���Yy�pw�f��D�_��0����Ξ:uS8����U=��\���~��*t�Cc�F�l��+�s��%c}*�!)rɪ8�|�֐�����|U�?�����o�����y1>��~�"�4��P����4�L;��6�����B/8����-�n��<PK�dV
RaB���c���(g��A�ѫ��Jޟv�U�Y6�-7+������#�m����^����"+6��N�˶��R�� ���{WK@\�&�ނ��3#N��j~(zd�K�d�$��t�)��(P;�ۤ�-��Z�)pYxʒ�rC�R5s_�TQ�Ѐ��.x��	+x��]p1��0��F����`
kJ���`�V�4��b�
G���OlZ������n��n�����0� ſ�=_�Z�A��c؛�0I;-;,C�I[;�����S�
�$��5i��y5Q�����g�'�����;6E�$�X�#3^��%�T��e�i���'D��1%�:�J�s!ѫ���[.����U�Ě��4N�������Hp3���a���q��fm%�P�&�\��B���t��	���K�pW�c"�k�簡��������g��h��8�#�	41��I�rB�5���=�b�e>t���D9�a�wB�B��F�'�L㊣G���otw��m��hX�׭��$�6�Ө^zZ�e�wS��3.y� �<�tެ��v��G^��v�:L�a�lȅY�L���ݍW�u�cͣ�X�NWס��B�s{@ۀw�j��7^��Z�wq)Đ��t�Z������7!q�c�x�;��.���Z��޹�����Uz�"@I��� �Q�ޣr&t���
� �3$w��Ӊ�H3� ��*�<��jʤ���Š�TmĬ)x>s�8���[JܩJ� ūv@4�e�Zg,\ԣ���x��ou��d�r���JX��3��Ώt2�$��E��� t���zx�S�`��N��p�Ր!��[�B=��v�L�%�����{�f>p�ow ��Զjd��8oQF���,��e6o!�%6����7`�ih���"�'8��r�7FP���;
]Ԝ��hz�_?��M�2©�r;�/��^���/Pj��w\�(���b�����v]�����*��mcg�(��QI�{BA�pNCѰ�r�H\%F)�=���C'�HhC���q��M��/�O� ��WR���4^K�|��vlgX���t�>>�6�o�F$2Z��3
����Vq�&C�U��3W��Ӑ�����^�mx�WDLI��n+dL+WBN���k���lD�Sh�@�S�@��H�h�Gj���Q�"��ˋ��.O� �-R<c�x�7w�_���.��u1�X/���R����Iq�9�@��a�[>cK5ل��x'-�Ԙp�ٰRp�y�Or��rh{��W\�l � NnA�b!W�=���b�6`ب��U�&��������h��I���
#�yOpP��c:��k��ÿ�.��$q��D;ɚ�;��/-��+j�71M5�M��ߖgL��w7���cuo�}f,C[v�4P ����B��ڞv�����Ҩ/=t �9R�|}�g�����
�W�`Pӏ^5�wU�����;h	��R�\��Ive����D�����>j�_�Q��V�N�"Ju(�(�6'�s+�1@�5�k�o-/����p��:F�P(-�t	�c��J���qu���0�t$���o��r�* 1f�3dU��'��Ȣ��2�V;��(ų:W��X���C��tuO�t�/�lo�7�z��̱�(����[kMx)�S����e�~C�+�*9gt��6���qAƶ̟jU,�=�u.xz�W���ZӞO�A�K0��^#vMM3̵����k��B-�8�E�9�&~앍�c��'L"]AvN�ۛ�p-��/����d&!9@�.s�V\^D�cI����`h%Y�$�"����!��]��(��#�i(+2��?e��32:�H6��>�p(�?�d�d!G���xfl&(=��\I�=w	Te����Vrxơ�c��b5�T�V}��cM����6���o��a��О�o��(���0�F2��E����ꀍ����5|*�7{1�;�i��� 0A���^9D��TW���m��;P7�H�f�$�֋Γ.�@�)c2�s1���PRX�+�������!\.�V��?�Y ��k���Ͳ�w^O= � �N�������� 
Z� ��D|��?��V�|H�gq4�U$Gݍ%>5�r��T���`�	�"O�HeW���Bj�R-�FTD�փO�+�z&S?L��^��TJc��@I��C���6��5,]Γ(A��d!�#-�i4$Q���>/��Gv��C*����<&n��$izJX���RypxE	��[���"����{ X'��պ1Ե�a4�<B�F!/5��P.?\�7��}'--�?�ݨ/�"s�U�`U��75��ǃ���l�o�
W}P���2��!"��=�NSb1���P�i��}��9���� ��$G�.ђ����c	 ���֛�{����U�uy��bxЌ��[��Ա��(�p_MP��1}2\J@a�QT򁉧�.i���`Kt*������,A��4�k��<g��\���g�L�k��E	ob����t-��Z�i�qX�%T�nq��	���Y�$��>x&����B"��Y����P�46����i_��!����ʎ`Dk�ߗ��ɛ~�:h�m�xk2˦�s*�%|$|9+x�ܗq6�j�yJݮ/ �`/���f�%����_�7�y������ ��u ��A[׵���
��Ld��[��O0h��`o�A�a�d=�~�H"AajiL~��T?A4������P)@���jޜ�F���R%^0-�Lo$����_1s� nNbg�Gy��d`(a�nd0�(]M7ݹ?�]���2�O��M��֔F1�hc�I6: ���Y�:���fA1��(��2��r��z����<���w���vW?�H�K��V�f�u)o˴Yj�� ���j��1�`���`#rֿx�OE���2���r�$�x��z�jԵM�_%J�`Lݱ����1(g�e�-�6Ia���K$r���}��Kv�.�� ��9�$U�`w�g��01}��3ꏞ����h�f`$�Fl'K*��Y��2XdS1��Q�QŘtȷC����N�{�n�����b��	/;}AԤ�Jg�F��8�G�9�+U�y?UgK�&���"�R�w�����x�� �Gf�"������jŗ�<���j� �T�H0��d%Ry��� w�JF�p�p��� �Ǔٚ�~�wr� P�)`�9�d��9�q�{?���:@����hoZ��&& M��3#j׋�PPf� ��w��eo	��{�q�ٶl��)O$�&�~�,'�74��f���Ta���%fi�3-L�8�Xi�OF=[��hb�{��(%���i!ߧ�d ��k�� ��t -=ƮE-r�������{ ��ߚ9�;�wޢ���#���g�|d�x��ocS�;����z���[ �����fTQ��r�c�t������N �|CwDl��h
 :wRN��N:�i���g���R�x�2%[Q�O���6��t��z~K��a���%�f z�yY�|�s�ؚ�[�����hjm)U_F%U���ONa��A"^�Af�~kd�?DpiA��>�u+��]c�>�$N���k�c��RZ	�� �v�@I��[�{�w���|�\���L�33�%a���)��]�]�z{I��R@ԅ^�#�}��WV�虔��]ݮ#|��@�'f��:�A�~�N/9���=�JK�iF7�����5:`���=�C����}�3:|�����H#M�<ĸ��)�`����@�"�,aT<fб�2���3�_a� @w���,1��k�;l���H��L�yF�9��A�ɧЯ������\�㥢��ǭTڐ��W��EF�d�����T�~}��
�܍s�hA�҆0�*�;ك�N���Cƫ�~g��v�����O^)c���e$�Z"���s�(�[�u�Kd��;�-��r ����͕�+H��h(]�����}wM>�ѐ%P:$������U!�F�]!�m����Ԇ�%���q�%1�[�P�yTD7o��=���2�3��e����Q|�1��	#�/Y��~�n�<���v��rI�3�@�#�.�s`uT��}5jEW;;�]���z�-��֫w�ZG�����v�ۗU�]ߣȠ��+)q^c;�o]I��t��m�^���w p�������av4�@�>��W����&I�.8���K�y
q&�'�(Kcu`K|���k�Q���5�.S8�<V��`�i��\�e?�"��t��A/>��4O
T$� �<\N9��E>ۻ�:��4ַ��mm�-�݇C��q?mZ����/�MJ�dv�X�+ҥO�Ф2��J�u%X��y>�mӆ"`��}"��@�!Zc��]�eI6�q�U>^�:o ��j�Z�4l����	������o�7�Z��ѽ-�9L���/U�$]����k�Rê�W�浚o	?�+p��g~`'������('���j�j��ϺF�(�j��]��U�uD��'T����7���^?YD�aR-�r�gS1�;�(�NZI�Zr�W� V
�M>����{�P� l�{�T�}��ϑ'����[�����y_��yȪ��K�$�+7`ǒ%��'GQ��Ȋ��;��X���O��e^`c�R�>��T�[*u�Q�� � j��
�s�G�p�3)�J����;#[<J�~3��&����O�s�.O��k�.Р�/nk���M�}��_���o�#�y�nȍ���P���&(ؕ.���΃�Ur\��|�ٯ`<ނ��e��u{�����-`CH.y��t:IKWہy	0}�#gf�$d��ֹ#����"be�::6Y�c	ꇓ����F
�Z^`t�T]�)T�2%�ۧe�X�.M�%5=�Cf�[�M��3�Ԗ0�K09�Q{����:�*�cʀ���� �rP��H��':4�@TSᓱP�jK�F��Z.����2@l_��v�Z��:��i���n����#t�9�Ӆr%CQ�����isѷ�S�7gw�2���}�Ʈ���T��mj�a��I��3�5P����=��7�}�T	wip"��yŒ��$#��{��,��R��R�����������BD�Z�OdS�(?&�-�G �S��`BU��2���o�
!�.�j��G';��l�G�od�/�)���P�!o����u����W�=��F[-�j2IU�BT㇟.�%5�lb�5if�縓"�S_� ���)����&�
�vl�:֋(�*��䘶���q�h{�m�|��4C`o,���"@�qt��M`jĬ�c�M6�dl�p;{�|��NX�I>-B���U	̩݋<�a���M��=�H<r��\��xb�S�e��q�u��k����;��JW��Wg�%r��`���b�Q<���)�ONH��8�9�M8ĲM���e���Y�m����-S��^n
�	�/��ct���9FfC�[j��:H�p�'�.Ϧ���̫G<����l�|���N�NI�D��JIr�/�yڹ=�d꫉@sJ�[P ��y؏��#��}�"���{�X����+�� d�K�޾���/'�p�0��^v�XA2��Vvw� ݶ���Lv����>�3œ���+u��Xf6�Â'C#so4^�����"���K�4�Л�C_}U�N"\����P�\�eL�3Cz��S�w61�{�%������H_�͟ov�y�d*Ib^!����O�����n��8�4����1z��f��)u|ڋ���5Eh���{�i�YۇW^��8���T��]H�ONvd@���*0���C�&
p("�Ƽ�q�t�MZ>���{'n�K��]+��-Z)-&�y;���IrM.�u�P�����G)�A�� }kA^<i4��CbT�i=�3ʋ���^0;(��߃Sp�7��(ڬ��6ԋω�}ή�����`�$ȫ��;~Oe_#�8ژ�P(�ǳ.�Q�;�i��w]@?|icʹ�9��m��I�?@:�\�#��҇��g��ǟ:�0Wx8��gE��x�x���4.jо���W���0W��s�E5~h'*�0��C�J9��}��B�P�o�k���ƥCW�48�
T���4ӏ ���fl�w���i
�K�ot9�u�[��a77���l�e�QԞ�30��Т�<%D�iI$X	Z�?�"^Do�S+6�\s���` ������L,���� �k�}O�K0�_�bJ����Xg���ÿ�x�J]����p�.�j����*���i�Q��Rs��*�B��`�b.���K���><D�tf��lO/v[����m\�	��Rd��u�LU����}����6���*�#�.޲��;�󮥻�j�3x@���2���s1:rR¦E=�'C�@}���&�2M���QSvr��p=�S�K^*0��E+���;�O����@�M��jB�mE�L�uT}�uEqSow�~�儷1b̑=Mc�Lv�f7&����&���v�7���S%螱�Ɨ�w��q�)��UyNI����4��Z`hH�Z�(���䘂�:�6�}�ġ[>1]_��Лd`=䩹O�M�|#�=p�[�e�@`�a�S��ģ�A��T�@@�.��O/%��};��:O��WS�hj�������h���؏w�Ht�#;(uD�������4�#��aC�q�J?�����x���?31GIrs}E���i���`�ʨ\�,�r+���_��>���T�M�~�a2ufFyE��N<m*m/��փ�Eh���MAP�A�L�����M4*H,� �f%�ˎ�H6�}��DC��Oy�|�3+�f6)`óP*2�C�Y�W-�G�ڼ_k�����n�#g6��E����%�6q�3(�u�DK�;��4EPp�}0�'���6�j�"/�$('y�p�L����ڂ��kQ��A��w �6��ϣ�s�Vuf\4�I::��x� �	�(��&��?[��'2���4���$�s�u����7I,\�hGIsY|h���O+�� 1�N��ՐVfG��Ê�(���m�gZ౭s�'e�f�u��$��=��9��`�*u�<>Ku�3�
��]�_�d�Yr���3��:����޸n�J�"9/�~��k�K������Z樼�I]F]�C�qY=%�i?��1e7c��PP�l�A�|��v[fXgur��F�M\^/}��;y�T�c��[���O� �l��Q�2��Ĵ-��4��N�����Co�8tKpv	�1.��a��FobǪ+ix�,7b�h3��#��F��=�V�3����;m�8�A@,#о�V����;{߀�"϶nю���6-+�ؾ_��ش����<P?�+ʹb� �0��>(�hΏM�F\on=QlY]P��m��� ����7MGV]��C�l>���e����~W@&;d��WDU�V�<�\�.Hf��8���uџ�Ac�����j����7��'�_k�������;��,����2��*�z��ے�q���<EȀ��Ҁ�/���_�ld�@:��m���(6a��J��$-_�ͦ��v���y��Ǩo�<����R�!��:��u8�ϵ蝖����;�=Yas����U�.&ƿ)&'eY
�=؄U��m�z���.�SL1�](�,�c�6g��Ϻ�{d�c�L��7$7KV���s?��CQ	/����p�p��6�c9��mK�Bj��+���p��E��1�no�j�Ԕ�e֛M���5�l�N6���h0�A- �J,H����KJ��zqJ��MHcj訙\�ʨ����`��P�Q	��̾cޑ��an��"Dp~���x7�����iR��IV�@�aH\�F[�!++*ؓ���Lb���q�C{U�2QW��%Qr(�K��1Ӡ)��^"C.|ٴ��¶e�m�:��0QY��C�{-&�|��c)o���Ɓe��j�o�w=1R�����V�m|��22S���5�Y��Z9@��6(��}-?Zi�Qdc�)����'l�5�/�?�`iL��e4�.�-ht���-��Tv;�O�����|��_��
��Fa��k�(�G�#<P��i��YlO�@������:�!����k�а��5m�M������Ϙ2 /<&�Ug�R+aܝ���1V�@*����u�ѳ$*]0R�����r�6�,���k~��5o�0߃���D{Rܛ�3��Y������M�^@9�P,���Ij����Џϝ,�Yxk�F�=������w����\�u|��y`��kӦ��;b}|�{+G4Cǐ�­��2˰A�=����~	%��\�X�e����(�Z��[�Ot/5\����uBrkdX�C�1�)T����y�"�W�i� ƿ�/����d���N�,AZ����9?���E�e&�8�'c�ȿu���}ɫA�T������鰓(������C"�'���Y�GW�֎�O���s�T;�ϫ��0��OTi�ow�%�������in�|���7�i`W�,��Y���V���'��{�D�a2�{q�ϙ�^űq�*��=����N>�(L t�č��]rZ�+.�D�	z�'�k;����ޑZ�#<Eq���{��R�Hvck���~E2/ C���JYn$�����������NL�-Tl�<�[����q��
2���{;��m0d�\^U!u"�s��b	�ٵ��K�t�;�XT�V�~�`'�T+�ҡ���-��Ӭ�)��&��B������`�Hv{f��e�� N-'��?�I P���$��R�~-�`=���6�U�D��B�p��5&jg��kpX����@{7b�h�r&5X�{I��|��7��hU[�����2{�u��VD
�7&3!��v�y��ZT�*Lc!|�̄�1��)��"���ü��U��kV���>h���o(��Q��d9�pQH�xBn�Ʉ�揽v��$�9\���Z|��9�Y.]�a=���`�)�ucj��O�����&���1�0���X�?ͣ�c�3�O��%��'e^�5AzYd����B�]�#uz �@O�#y<��r���K�#n	(I�9��i�q�,p��4w͈A��zL��d e����Ӳ�v�Ζ"I�9xR�Xejŵ�~���q�l��j��J��<�V��h��/?Nj'ߞ���o��[mA�a^��[�tٿ�S6Ѱ;���P�����B4�dT��`,�G�ck��`�E'��y�$�C�F��&��������eKG�q����,�R�e�^Ve;���a�Ҧbf�{��7����>� �!^��e�FAC����?�UR�Q+��kV�y�#ڄV�@��o��>�7Z
4+�q����^(H��0�l�<��A/�K��b�
�x4Kr��^�aO�"$�����'�u���1�ub����ٽ>�ĽZ<���HS]�Žde�I"�ux���l֫k��P*��Mʊ�Aʦ6T2��Xm��#��#�%f8l�Nls�6r�ݤ �"�uF��SJ-8:�����z�7 � }[�T��D�˹,4j+oY��R�����e�[Wȍ��R�:�����P��"3�ȯj��25��]1YN�{'�m�ܽ1yC�B��������\��ԙN�D����Y:��$	�C�	v�_���<�?/p�Y
��W����;&��~H.�¸H����'T�<���}�\���������{�w�������4}�����Ù��^t:o�wՂ�}��`m�(&�W�Qw�C�8�`��m��]B�ZG$���)����<�7��y�^�/}�{��z�=��wԩ۔E)jvGy�,R�����&����+���-Ah7��P�7��H[��3��L3��`u}��Y�hS�o}��OU�����HhV�4�a��=�$h$���*^�ՉL�d�_��
�'�('� .��Y6h
��r�ۺnʿ��/�fq�/�uJ��g��&)Py�s��I����J���-i?���Td�%�*���v���n������+�v5�0"��j&7�J�h��`Z<�B'q�b�ߢ>�(��a�T�S�����U8��P�7�����"�q��]$#��J2��`�|q"SNڢfU�.�Z$;Ecr�?=6}�êc_n3Z���V,p�_⇖xABq�aZ'jSi`��WȤ�}�[r�e�`�# A�u�0����,g�_JO|�;�"K�PS��>��#���3�6,On��e+�"ʂY��N�g^��D�I�p�'�K�1S����ښ����ա��e�Cn�`ri��L��OIZ��ZV��,T��u-��@'��ٟ�.T�zy�Dv��M�Io�h���$�=������������?1<�	o����ѣ�x���&3W��['��,:�`\���R��5E�#�&�3�@�t٪����k���Or=�#f_+��'%�'�0�KKS�>��Z���,�Q�5M�C]��b�}�G�H@u,��7�������f�o�q"�On����y1VL�����r��)ȿ&r�V�_��hȲ����yE�K��)��U��0��#\�#d:�\��-U��'PP�g�9�l/��J�ɻ�e�LL�f�Pы�h�k����؇����#s�j��V�ޭ慣g�O�6:���7��%�5���u5����td��xv��	����ְoЈ��4�q�4p��۵���Q�\�&�1>�pd&�?��qH+�rЦ�E�������❻dIq���a]%��p�|����(gA�dGjٮY�A�a�^K��NM�J۾/�؉�۝�
��5�@�!�)�r��<����]��%��&_�Q��9H������{s���� B��qG.h� ��?J>��7���;�O�F��~��$�@=^�W��v5�����`�A'�Vk�g ��U��Q]�{�sk5�O5'��IH�f�3D�X�)}�P�`��B���I���o[�L�_�� �CB������4��CQ�H]��_5�R�O�O�,�UD"s��"l��"a6�X=[�.�)&')�͇�6�l������+T����8N�=����w���ev���$v��%#�9��aD>	���ٿ�'"N�:p�n���L�$Ђ�k�,�r�6��M����#l�&k�}�Q���;|i�AxY�w����^y�}-�*db��p4�� ���("�@��1�_�l���J ��J!����g`,W�����䠥��#��A�jq 1���j�-W���}J�~5!'��ו���zE_��i���;G��W�0�ȥ���6�U�t���}��U^B��B;�yq.V_dF�� ����:���B��^˨׷�,Z�켽�Nv�cwݫ���CM����t&=gg�?e����45_s�Н|�[��|�^��&�ЗV��ƽ/5��kA�l�`��!��?��1��掵��>���&��1��,�v�s�Y�ŷ2�~�1��O�3{��3���x6E%�jS��#���smh3���pf����'�t|:"J��#�D�%(E��Æ#��1uv����l"��v-I�s5L�ڕN���/��f�m�b�+�֦'�IwIo�I��1�|B��acܽN#���Hȋ��%�F������������	�j��1d��ya���1ԯ��Sl�i��^,�wg(��%��&���?��k�*�"2���9�6Q�V{"���7���fV�\�ڧ��#=�f)٩.�[ֽf�,+͓���S�RPX��_LVc%M鐈�ѝT��'r���|�q�lu!t�rP����[)��v���A��
T8R��d����A¦����ڹ7�G�1T����=fZ�c�`�>smV�|��A�f�O��� �V�ĹbU�������n���b�ثN�[ya��l/f��!���ͻjz�{S�v�iƻN��〧�G�%�b�����N�x�(�,/�9+��n:ױ�`��гS(����$"�> �/��3c؇��06��xG���$D$�����Ym�I�y3��Y�7mp�b�W�5�PR���!ąv���U�/����
{VD��v���3E���vP�C0&EcF:ohM�G��!C3��cVbV��z��z�&��.Y��/`�C��_�Ќ���!hB��Ѕp�M���0���	�"\��Z���l�v��L��a�"�`O�^�Z�<�5�<�����b��O�p�Л��&����87�2�%�7��|UpbcZp�f���۾��9f��a_�偸���l�Gdao2;$��h��|�tZdd��Ůw��찭}[�H^ �1x�	��){�LthY��<�/6��W���J�uњBӯ������]�s���x[�f/��cV�����SC�@P!"Cx/�t�ϛzޒ�[����~>���k�`���5Jh4��pm��Ӕ���6z�Q�yϮɧ����}��ޅD)��Mȏ�{+iS,*�LyՂ��X���;Eb�%WZ��:��xsewi��̝���5� (�Dls�g���*T��\f�G�չ�]�����(��s|'��ܥo�UYL>y����L���>��4e�h�Ⱥ9�oʛq8������%m��UD�l����iǼ�d7�X/�f�h*[�d_���Z��-�������z^c�Ҥ9�/�%(�7F�'z�Z6o)���-��U"�c�{I���R}��L��l�B�J����M��W�"�gs���g�/'�7���;b<�}#�O�6MY����ڲ8�X�U؍�O9�w����F����Rs@��آ?�yU��9,"�_���Nm1]	�R~�GJב0�?��VL���1��aw�W�����Dx��v�}m�	�Yp{)0�P޴���"Đ$>�xx!�Pr+i���{&(��KF�D��kW,�l�ہ~Bu��hd��������pd�)�(����븜Z�e�t�j�8��zwH� .*z�+�Ud�l:�F�Y�؍�����&/9R�T�G�f������G�0����e���f�=J5jF<QY���΄��~_l���ba��N{�8�w�|h���V٠,������'ڛ��5�iW�:�_u�3�(�\)&K���ڻ WW�k�����b�7~n���Y��9�h�R�A,�e�wi�t����yy�^��%�f�w�u�K�-��)�����'I�� �<�'�R�ٓ��F���(������2���}��L�TR,�$!�2����E�d"!�W�O������u�f���Q�v	T����s,�D8�@j�i��D`��%���	���ȿ)��8�F�e�Gu(g=�ia�\�d7�I?1�5~�p��c�ڈ���	qLc�@���	gqF���+ìW_�S��KkK	��NDN�RR�j�@��� �,:�"1z�L|9|Z�fŬ=r�B���rג�9I]_��ec>��+�W���#s]0�iLR�ϛɟ\U0F�b�P��"Z@�'��O�#��dX��e���8[�Z�Y,A?��ܜ"@� )�Y
�X�5U��ׇ=��0EO����mN!��`�d�hy�� ���s��^SM}�����g���"��z�gseT�p���۳�o�͎V����g�˧ը7f��;dZg�T��꧶�.�T��k����5P��<�]5�2�]3��gdq3ܵ:�u �Ѯy�m4��uѦ69�V i���jH�)�C9���-�������Fn\Zwdt���b/����rZD��Zpo�`�^�(��|7w��YԷr
��p{A��Ո9w�
�]���(j��5R�y�R~ɦr9o����]c�I����zT)��y�ᮒJc�p]��@67, 4p���ӊ����Ű�F���G����.����\� �Kؽ��Xk��"T��]!>[�����O���u'߹AS\֣V2&���d"ܬ��O����|��/ &ޡ�Y������n>]��b��/���!�nY��&"$Y�-���`�y ��ɯD�[�$zj��';�^���R7\�wT7���b�Tsv i0"Dd�����7�^�WJt��T:OM�y���+�t��Ƹs�~�q6j�A)�
���=1tg9n:< a5Y� Z����G3�����SЖbs~GA�M>���յz3��δ��?H��&)��y�#��
Rr���{Eos�R����5��5N��y����&��;�"'���~���?�c����=�٥�m����9�;�1Û=�#p�eg������V2;X<���e؜f�c`�5���hb�Pf�Ȅ�/Wz2�<Ҡ����Pch�*H�#y����T����W\d�����As]V�c9��F�Mn����&g�}G`�J4��r��W�-]t�JoTn�����t���}:g�tU��8v-���	��1F��h��b�N&qv�ɧ��y;�xm����l1?E��z tnL����aU����}ts�;g?i	Ӆ�ԩ%uf�2!�SG3���pi�hf0�7��0�&֊6�3n� lΓ�GI�����!���$H���xWB�~dD%���t�ҏQ�7g3��CىZ�$Qy��+��iI6���2&VИ��XnǕ��av��ri@V�����~���a�{�Ͱ�瓰�[�n�kyZTuc��I�?�y��6�at�/P��j��JT���n���ch5 � 1,h��^�[�-�Xl�0�(�dS���C�R��_}�/ی�N���a��Z�7���9�=$��M�p�g�7w��y;k<i��+qY��AT��s^�¹'$�S�b�$�)����������}b�\�a+����!ΰ�V�J#��>F/���cm0������I����� .�f�����=�T?���盜�/}T�sD.�[%�WC���O�R�(�{a��ao��k����
�N�h;0T^�c�YmZ��E|}LNX9�u��O���� �aHXITl��m�F�/O� 7mH���^������ =9�:8U����
���ܽ�2�¶_y�|7��I+^(��s/�k�n�����̈́�S!c}8p>�4Z�K�s���jC2�3�]��j�JJn�^�Օc枷�^z?�X�Qy��7+g�N����@��NK3�g�H�*�� ���e�-�#�Z*@Xh��h���o��M��iF1�����V-����7q��"�v�[�� v'x���+��E�����F��߬�� ���7>	i΋�_�t$��|3ִ~Ih\C�_k�"�+�ASfy@���K�O�����8ӧ�S?����l��a��<x�e�	C�Qf&�N�)��0K&�y��$�����%8�`�s�n���K]�38\����ۤ;�:���Z�,��EjCҾɃm���K<���C̄�E�{	�ńI�o9HZ4�UZB��Z�ԕ��O����^����_ÊǛ-�5��%�\��W�0[a �\yNP�/�T��Մ��;~���qLd��/F��1�ea��T����5���ɻi&'�����Z^�țD�����D?%<s&=9|���eT�?Gk�-7ͤ/R	Ue�N��&#�+m[��4��t���(7]��p��RP;��C]����/5_H# ���:��?7�\�y2�=\��2�	�cl�\Y{�$�zJ���(*�T)��>�rx�R��;R��	b����� ��@Ld������ޜ�Ƞ)��.����.Ɗ�qk����^�!�>>Z�s��+Bf�&�����b[�F�B�xMXۿ7���k�`e��ҭW��?+[���2	žk"�fϴ���r*d����"~�|��:���q����X��@���gN�̉�w�w!��1��,������ܹ;��"�^+*�!�R���f�~o4����K����a�;�ƛ;ю�)�%r��V�'?��/��Pᴵ�L,9��̶�0ge�i���a^���YaV�M$0l�>x�� ��-�*j����w��[ �_1�3����D��;��]Ƹ-��0Ys������Y�kK9���Q��բ]]Lő$q%�K�P �K/�u�,RS��� '->Z"��h�u?\��l��R��J\�0mtP�^����!��+]�F�_[�o�(�c�	�+��Ι���Kl4��u�����iǡ�I��7�R��2��x��v���ﺵߎ9;x��k��e4�:��SK��`�n���Jvu.�Q��{���?�ȏ+����2��k��K�r������1��;���CŖ"�N���}�r�2�)gv~���XJ��K�7��-����$I���i��^��
W(�k^����ȼ=����n6����hp�7^A�L�����`�!������9p�'.	=U1G�pzOex�+�R��i]���ݍ3����s�qk�^��q��1q��g�����F����2.��4���D_��p�#����<�9��gTu�i7��B0���$��R.�&��qrB�ՍӜ�Q6k��H��sDD�;t���޷�S�N�����\6�����M�m���U}r�����u2V�7L*�qf�C8Ŕ��&��9�8�i�/t��a��9�� �b}���fݴ��������x4|"4p�-[�����1�T@�$"��h�����F��4�ߢHm�4��{5��BC��?(�D���ja�՘���Da�(5èARLF�t�Q���K���R�QB	��rk�
�[�.�GQAFJ�Qd�j�3�j.���0&h�hg�c�I4fޒ�����9��|'x����~��)z�ն��Z�I
�NK|6G�?��D�B�ޠ�-+�`V�
��Jc ,��H�[�Po&�막�i_mX)H%^ԓr=�%~����[$����e�Z�Lԫ�\P�u?ܼ���$�}G�ť�{�kJ`:�U^}������Q4>9�~cHN7xq�CD}V�p�2�as	�S�h���������� ���
�y��% e�xh���@n��Y������@V�w����v؊�}���Q�U,�®o�a��e�k�C/����r�����(�i���jeQxĳ�_�α�P&Z-��Zo5�%��4���Me��
�`D�4�:^�m�qi�W��z��#y�M9x&,ls��� T5�B7i��:v�G!/Mr���ɼIM���B�/M�Y<���\�ĵ.��ڤk���
�YUU<� m<~V�IF2�#�`.n[0�߀�A]���@/����c�{E�Ìv;L�9`-��Ȼ�$�<��P�J4�*A���J�l������4�u�$�}DE�ь��!Ԝ��xRhi�, ��K��"�c"��"�n�1����\�N�����7n�@���k��?���g�1��ɹ�5Y�|r�&�]U��VN
کH��ɁΌ\�V.��"�m��4PL�I�>C��ϳ��8��H�$��*3/��b ��'�%ὧiN�&^�q�#"�\�]8ݚ����qŅ�㭠U��_��>亡�8����yB-��)݌��W��*09�<N ����-e>����hSس/����f��'��:��a膁'+D:'�r�.
{ ø��6n��ԫ>h&��>�_��S�w�cm�֔>�\�WiiX.��� ���S�#�z��A�	��V&R�lM��ʨgG�tȎ$��	ҒMF�$hjQ�lڂ�
+47'�X}���r��3�U�0����-� �[(Q�ag���:��%̿U
��rK��{�I�Xz��;}N����� q����X0��� *nS(O4s>���2P��|\���gV�����6�N�J��Vq��<xFW�2��6�_gδ0���K��!��qi㣠�e����Yb���������~��
�gʮ��܆G�㩻$%�5����5��Ï��Jx7ofa���8/kx3�߈[�Y��w8{�h��#2w���'�e��2
�������J�'O,3�����/������*U,E73 ��T5��mҎ�M�;�EJ�ܝ���#����[߻��o��Nuw'v�X�Vp˦Se����l�B��<��s��S	��@��'��5;��{���/o]�_�j�Y����HN��v�t��d�������Lħ��0��>�?v`�U�'�yz����}@��&]�H(5�6�0�5�g�iǸ� 7a��1TO1�<��ܥP�S�S�M�?�.h�(�"�%��a�����"�H,�L��w������]ȥ����S�D�̹�q�ނ��˲7od� ��h��pc��K�䖞�$	��JQ��B^%��ѭ�z�1��8���uʰk̞�P��@�"�����K1O��]���w3�}�ȍ��|���X�#�L�����w������{��&�u'�645Ut>�^�7hM��Tw�|�o�c�����5(yx��B��9t �.71;}��~�XC�ڏs�I0iG&� �AL�� �U`>�Z��Ѡ*�����x�h.)B�}f���K�upR*�߸I��.Xy���Z��B��=��ʊ(���t+�tx�����{f�]�}�&�}%@��[=�]C�`tC�$ͅ\ή܁�������(�k�oA,R��L9Ђ�J�A��v�gh:ԆX�d��%��*�e��b�� ��ܜ*��R0�;�����V[:Qօ�okI���b|B��:��z��%N���ޝ�`< ���DB8��
I�31A�A��0���=m���jg�b}6YU�(l�T���yc4��~��D�v|4�w���������Y�![?�#���r��+FwW[�]G�8��r��|�'!l�7��W��	i�v����삝tN,�>αJ�)j��Nj��{��(�D���!L�󛃝*���`�6�֠'j�;,̾���#�� ~�U��tq����zćˇ%���!�Xˇ�Ξ�g�3Ojw�CU��"/&g��l'rF���1�{��x�h_[�'s���81Ʒπ�T`�&f�%VRH���l�jtlI���.��4�/���\�O��w�
��S�-�$'���i����|2��Mk��&��-��L��V�����v;�kԵƃ.q��'ڑ�xj �ʰ�E�"�A;E�J��W�U�!Yt:����;U��/�oA��	�c��:���aĖ�J36$b��8?�P;�)��dI�C�62Is�4X��@�S�9�v'�H~�	C�ӔyR�&>�^	`�Wy	��lzB��>�V�e���k<�:#��)q����En �#��7c�t��U��^�E��;(\y�Z�I�O'A%�t"�V��	3ȥtqX�>�:Fv� �R�n�F���,���|}�K��=�ݎ�/�E"���������^�a����}{�P���������!�qSx���D��<�j��gύ�&�o)������CI�3"���o��4H���''#��|��%���G���i��iv�Xdr<Lޔ�s���gl��Ђb[΋�W^[K��wIg�z��.����'�*���<�T� ��e)рE	��Z��J��t]��d�C㩢���a\�����䂲���]���5��!��Վr���3;a�S��n�}�ܷ�h�
��V6U؆�O�6J�U���VP���`�gUa�X%m�'~5��ܯZw��'Ճ���y+������<8�cu�����Ə��|��Ԫx%VD
�j�D��[��p��f��c������XD��xV�g���1nS����B��yƦ}o3��p`�}'�P7_zˎ�F�z�a,��F��Ư:��@��d)�Í�i��Vf��e�+4_�F�%0��#�L-f�i��r�xI�ԙ�y��ؙZT:�	��Y�c�Tk)��V7��� G,�]�>��C�#qYrl�ϱV:��[0�xX_�KXW���	�|�]�b�rF�e�,#G����Ze���Օ*i�?A���"�֒7жAm���|/;	{�F��]b���T�5a�K(Ub��9Whb<��XD7��=Q���Tt�b6����n�<��R!��>:Ci���Y:	�K"�`�ܼ)0�l��������i�FaQ~̑��K��>t��S�b�%�p���LS�+ܝk�fa[O��,f�K��2.<�8_S�'�v�Ī��@�Nd������̓����_K��򸌘ա�_�w%0�����j����挶p�LO�&�jL�J1;f�̬��k�HU �Z֮M����k���h{��}g���(�o�����'�3cOf���(��l�BrI��-���lA��9q�Vn ��-bb�hF~�+��C	�2���n4D��!ݤ!���MQ���$j�"缿�ɭ�s���W�t��R�7J<�LCS��� �iFbÀ.�ñ�@�i5 ��Ո�a�.(��\�:)XcɆ�r��/�W�P&w��1K[�Q�&��Y�M������`�����2ѱ+��~�t1eA��F�@��Lk]E�9�2�=4�j�>d������Y����e�I��T����;XfOm���C�ʥ����|c}��VՖFdd�� �����s_�ﾃs�����0Y0vĂ�Q��-�����!�U lH�Q�̏�sɞh��ROq����X�	�W�P`���mGou+�U/����<�U޲��򉴘,5k�r9�������:����kT�0H{.[ԽO�	'c���&>h�M�w�ő�X��u����Oŉ��+.R�&l���|�0��$LԒ�բ੹oa`����R���G�$v>ICP���^�uEW��4CIR�'`����{˭���w�5%�cI$���{ֿc��D�3����H�3v�1_��7m��fe���ZT�/��z��Ρ��x&�ȎZ��U�����y�0��C�˙�)�C~��!��J^.}a[��P�OI��*���ົ&Rcl�TK~r�l����Bы��;91����GJs׺�\�3T���̻��܂�X+ҫ�������zf:ȱ����.����[��<Qp��R�`L����^%��$'��=�(���x�l=�o6`i8=O�$K] � N��U�1�%C�"���tx@�t/ԏZp*�������d=u�J�/�����bV�����/��I}'ٰ��~�T� p.05Ͻ�󪷁�ᯊ��>B�	���J���;�8(n�C���x\�jI�3ee�B�iĸ���,�o���8��Pۭ�x�*	���A�V(�
��mk�yo�6ІlEJ?�mg,�C3�d�bY�:� ��a�M⭆��31_H��Mg��1��DmxR7�ƋDծ2l�C���� ��U��MA|K�0�G�ދ�tw0���C7!��������`d1�<%
�_�� 8PA�C:m���}�Ĳ� ��׃�,��_�̽O�k�.��_��K�a	���-���4d���z#-�c�c�MxNR��[N�MOak]���`ɁH��/���GvT��6ݫ�R�	�らxǩq!�y^&4,B�������$uq38�+��'��Ot�޴�� Ё�c�r��	�L��[�4[ʪ���#)YJ��Ȭ�����,����ѥ>Boȥ�����\P�]�����1�<i��d���k�ܭ�.X�9[�b��s"�;��@��T��{@��Q����|�(C�B ��G$?3��U.
 ����F����z�&Vʻ:��1��a똲Ϣ���+�'.�(<Ճk���4
Z��9�ܛ�0�
���"�'�?�c�J8�� nK���j����6��Ӽ(l�C�ԱLZ7��L8�V�Tы��Ix���`:�f����7��.�Ł���5��œ�����se���+�rY!��o�1ա3o�VG�|,�P��Ҥ
�0�蔠��=�����_�Nmi���fjI���|��+K&k /@�o�ԁi#;��0��6�����ӈ��8��Y�{8ww�d�>	���N���w�M߷e����?Z>%��姅��L|�R\�,���1[����/ҭ�}��ýH&�u��j��#L��q�s�!W����G��5�t�a�����GC�ha�Z+�'�tv)?v@�-��5H�A���b���
`�`��
��"yy�˫�ơM.�P���ɞ�W��H���bS���������m:���I=��f�C9����2����7��m���Iǣ�һ��E]���(kƹ]�A��v}rJ�-��	���������	��C�m����:e�Q��,D}�E��L,M���J�]��Vh-�y����Ol���k5�7�yv`T����GMw��)��j�?p,��跐.�=#�V���J��D�5����%\>�ݡ�p�	Ƹ������+�%!୍.�qC{��c [t�/���,C;	A!V�n�7a#C���[�Vb�����̚VJ�߸߼b�\�����L�J�kĬ��J9���B$�%:u!���EsS��#�6�/c��7���
�γ���v�^��6uoƹA&��A�||W�Thf���+%r�?��Ѹ[���&C0ڲ�}*¡�D=��i�<�9�/��w�	�mE�&$�4ш?Q?��J���Ή�N��C,�e�}BU{�:R�����h&,��I`��>���Dt�������,B^â���cS�0Yp-� 2�4:�K��?��,�0��IW��(��տE�H���Gݳm������(1��%�mr��Iݐ��M�����nKyX��&�6mB��̉��mR��r�7*�/���؜��2|}�_?݄Pր���]"���}�����Eb%5��6|�n�<�7�Q�Z��LGv�͖����o��,���Q������.w��LT���.����	�(��5�z݌��݀�3�m���E���/^zHq/��� ��@��R���[>�y����S��,R*���v�'��8�w�J��ѣ)��Q�p��"|Prf���A�͋G_�t�P�[Ӻ�M�_�	��Ŧ�t�'|
�7�}�t�&P?w�%�w�h���b��Z��ЉM
}��9�������&���˪��m��]�b}I9�Ei�J�}�ˍ�/�ݓ��}�C,b ��$yo���W��諠)[��1
%OGfq	`��'K�7<pO���NP�f_���?��2A9?�~�9�@�-e?������>���WǩVA�B���&�x�G��=b�1rT��0/��|��!r�["cd���,:��Z��~۩���s���ScՑ�p0l���2.t��R�q�t��;�,k	��6J"d�Їғ�q�ߨ�v`�Ž���CGU��O5`x_RR(�ꅰ~�Ԛ3�2!�H�����.�%i�d7�>�Cl�9_+(h�����L��S���x��1��"��M�?Di�k�_Mb�Z�v!��{F��RZ�J �1�;Xڊ"�Xi��� â�h�y�%�
�A�|삨b�p��G�ؽ,zY-�EEE4:���o����R�@�p�NNO��n���
{�,
�'-�F�B4�^{��?�L���E��=xV���U��tO����/�K��i]eu ��fC e3����Y�CT����0��$���8�|h�������p¼�B�k1����Xr�ٸ��T
�C,o�����*�-.3�Δ݉r�
�I�
���S0iRB�\.b�vHjV�u��3Tߘ7Tr�o�lZq����
u�J���.iU{��"M�qZ�j�[%����pG0�i\jJ�������F:F���f�ؒ�6�S�vW��Ů�uIt��	6V��+f�T�7m�{�f�G�[�(���vo�6r^eyz�	7�i��+W��%�4�7Mз�O~�(n����%��8�y�+*o�WE�T���^��Ԟx����%M�(�pV!a2�O�#H����0�����Hf�A�������zI�;�ƾ��&��(���-e�)ه�@W�_㨠|�G�0Q�ky��U���C�d7�\�m(΍�YDJ/p�2���d*��"�\��#�*�_�Kd��ޏc�QZ�� g�b>���j�	B9l��|�Nu]r�*nK/f��� t棕t��އ���ލvBPunz����G���V���b�7�6��q�eY�#>(��pW���y~�k�ʹ���	�~>�}�$���m��^f�ۊŭ���V��3uF/�e�ذ��G��낉v�=�d��a�1Є�ͨ.�Fe}`�	�x�5��>��Rq���N�ED���Pu!���J�����Q-���^�f��\�~�t�K�a�S1@W�J��0Щd_��aS�'{��c-zɮ['=���#���WM�sR'����~�R�[���b.}y
�S�~�JZ{[�18�����g�	(��^d��h�����X��(	8PN��EKxz*�X��qM���@�ne�:�& �Hf@�M}�R���Ɉ{�����zo,���[9���MT=�;U��
���vǢ���������Sl�@�kk�(L��T��Z+E�b� ��~o������u=.����hv����Ք|6+4�J��Y]�0�'�~#jc��u0�ɢ�������ʞ���+�.���	�J�.�C1��ר����Pr��4�
�x�n#>�nV��=:�I/Y1�e������%�F��G�ۍ�G<�_�c��#r�����ָ7'|��/�]�(�|��P�O�5i��i���	��2���|L|�N�aς��(�8O1�5BD7���Kl*����v]�@X�����h�E�o�k��Ο󟏥���aE�>�a��b��"��ʪ7Y�kO��4���aA�z̀�6��>����N���%
�E/�Q!�`�`P�Ð�g�����DI�u��D�֨`��z���RuZ�ԀPO�>�����
�6D��:��>_΅�T]�mߥ��Qf�f���[D�� ��j߉�%\�Dr�����Ui/#s�M,�S� r�@>�/!�K���n�
��K/P���j�$��aLm��ނ��R��c��Aq�?{�s2�74�C+7�ZP��L�O�e�_a���2�bh�����>&����R�qQI�}�F�Pd+�����L�������w���.kW/l8�n�Rܓ�L��Q�H.��U�@�����9��wU�}�)��뚋�l�o��|��G��ģ�νjS�I���S�"D=Y�
�����ב���"���D�\�"��9�>g�w����W����%3߷�&�;�t@��@��}��b�	�\�N���e9��XS�$"��C�<=���ҥ� O�4q�e�h�I��S�U}��R����U��s)�4��������-'\q��N�tՠO鴲(�
�oF/'�;�y�5��c&��5�0C�P�Tdw۱�8D7b�F�̴���Z?+�	z�E-B5���/�՛�Yb��>K%�7�=Y?.�l&DdЛ%�i�c�Ƿ�nb���䯄��<5��0f�UXhI��l�9�1��YH^8�^���Z�0z�����<Q����a:d5g�h'3�'�]������E�ckK4���������,�(�ں��&ŇҭA�Ȩ�7�q*q��f�>��ޓI�d-�'(��(�{n*�3���[���i�!4�g�1mtq��KN�x3�ڧML�|�oqR{{iV���¡�Q��9Uj3V�fҠC��2t������؊�d�u�#G��k�;�.����Cm���&��ǵd��o�J�i�>�,ˈ+�Q���x���>�Q'$�n� ����o��Ь�Ầ�
	��.s�������|�p�!IT���+���3�d�(Bc�Q�+Ԧͭ_�aD9���jMP���Ju �,����d�����D[��gh64�)e��@; 
�%�D��mLdd��a�C�C��"�i�@�ȋ�`�����Y;�̷�H�E����n���Ή���K�
���M4��.�L��X�X(c%7�::���cR�m�P���"��C�e�=��,t�eym�,�WD�.�:�ס��70$qD���s��Yzþ������ ��2Po����Y./J��|ՙ�hn$QnNך�s�4>��:�G�r�I�6nZ��=̈́F�FR��$������,5�F7��ܢ�����%���\�n�*8��`�Y�D@���b�a�xtr��"���z��R�V��b+e=���!��A*��O��~��[��&�ֈ���s�51
���'o������d�H��a�2�j��a�Ā8�v(ڝY3��+-}��-���M6X�r���q�c���*���u!.�5���HY�=���H�z/���f�g�����r�����0F=��ǒ&��澧����!�b<�\��[L��4q]�C��ږ�������{Ζ��#�ъ�>����6��D�;�p��;0.��hmI&�!�7����j���y��������.�'}`e�RNr����{��S��.�oz�ЈS㭼 �o#�W�y�"F](��L���26�/�:�Y�����$ ta-#<Z_���e���Æ��[x��c"f7e��?Sz��M9�T�[;�T��S�`�{�=^77���LYJ�(/OG/F>���3�K�1ɾ��}x��]�,��$CH��lI��� �]2���NH1�_���m����*Q?�����f�w:���Ȏ���,�I��K+n*�r=U�}8�P�M����'sx�y{�#cQ#�h���;�(Wn��̥��)	��s�,�)�g{{� �<&�x��։a���vF/�!�C�2����}���|�:9��@��Pw�n�*��B=ΨD���U�����8"^�s�/�t&UE�j²;5/��$;���h����y���?J��F|��L�mc�J^�˗4x֯�^-��ŏ\�۪�nCjRs֜.�'�3��vn����,�Z�X���D�����8Y	�p�E�
븰U�
�8<���t���v��8���E舥�:��"�}~�oIq8��S�O��o�~�V<i���!uE�$���&:�Ub�dG���PP#�>�f: ��d�Q�Q�v�/R0�#��,��q0ц�U��b�����2��0a�$!@�N�9��أ��m����aE���f��@6�dх4��L�m��${�ﷸ�D~[�RI���3���Y>2��S��oi��_�
����}��Ճ2�le�Zc;J۸���F���2@'a�lZ('����T��J0e�ҹ��@�M���%W��J\��Ts���f�.:�`D�U`� ��
��ȟ\���T[��X�B�%����\$K�ѯ�/��:#��Rά4}�Te*I>+��R����xGC�P��}Α��Cd���qoO����k=��p*@�;�PmK@0� D%\w�X���C���ʞv��A�n8 �@��v�ф�E�	y6+��vKl���ס%)*ox6iZ�{�&#oX���v��>����j�d����pE���a��"z��]�L;�O�ME=�b�(=���\��q��C��N"�Qo'�U6������H?�v�J��%�����U���0,�NYK�?��y|���8}u�T��g����^ <��s|��O�b����$4C��01:�����yzH��T�HF�J6J��-�H�7ͬ�t�
~1�`���� ��H��y�J�ʏ��ˠ^Z�i/�/��>BL{3��f ��h2,�qg�J Z(^*����A�\p�Y-�������)�A0d�E�"��q\��P���wߓ!r�#���N��Jc��8#���$ r�o�6��~�W� �.�����N�7������3j�&wT���A���v3��a�Zx�7�|���tO��94aڕҖOʪ�}����_?
�;8l�%5#���y�����AΥ��b��ͺ;V�xO�>˫tW}p���tm�<�iJ9+	c�S�0F{��I0���[�#M?�ƙ�< y�­�E)�D��J��Ε��H�Y�pn�J3��;� &`�R`\�Ԓ*�!}��HdLlhV�@�wT�H��H]��H�������l���Ƥ�l_P��8^�vf�B.V'4���uQ�����LF7Z���8���S�,>W�kS��	"��W9l
��� A;W +~�ǗW��!���r2�yW�eņe��>��Fz�$�8L8ǝh���yB�������@d�}�e&4 	ʇi���D�:k���9!N^�G�`�Ο��v��<��G|��Jc��DOҕ`����Z7�k�87a7�S��^��>�7xu�>t��0T��$�p���K��<�4�=��Kʾ#�o�*�-�=�����&�UGX�1c>^����;�0٧��g�r`�g��v���|Ûf�-���ը��xL��(��FY������ãߨZ��'D3���L��j$��[�CvMP��b�o�o>��:ڷ�0V�/ �b�k�F�v�e�Oڝz��\�n˟�7�S쯩F��r�C��=iN�e��̍������om�=�]َ�K���	�g�KN���ܜ��Ǫ�9�6���=X,C��$�������h݄t���I�wY����Adc�`~�N�c�>��	��tX��|�v����{��F�?w"�D\���a��z�~�(>����]h�_i��	�I�E�눵}���`M�� ˯FXU���53>�م_mNǵ�
�rn�:��~�8�C0'F������+Z�oT�s�T��i�{���j����U6/<��J��^�����_���	��5�qH:�������]��;'
h�bN�L�����'���Wݹ*es#����,��=�ŬF���b�ؘ%4
%0�UC}_�B�u�f5�s����ʘ8�X!�~i��=Iu�~����3Ԇ5@�Ï23{�CqB_$%���#Uؠg�Ks�}%ӀuI'�8�~���l�������>����p%a U�>q�J�C��X�r����`E��m-} �i0�\��mۯfg���I�F2��,JjlZ`��uK·�D�w��.���7'��gC����ش���d��A��A)1&a1Hh<�K|�'}��O�*��д�	�VnmUQ��K���)^�n]������pvHqp�-���d~�B�[x���+��N�|�5�(H����OO6��/�}�i���ǃ��2F�R�X���\���@�u��.vT8t��K`�7���F��z՝�B=��Q�Ǜ�ᲀ�+�r��hJD�ⱅd���,w�<6"�H��f[������{��:�^����H�ͷ%��&��-�_���ݍ�q�z�hj���v��M���{�����?!�
��8��E��w������H����TX��J�6g�?:�6᥀^*΄R��mZ��Q�m���p��jE��z����P��pu�?C��AFd���.����gcZ-��Ҍ�We�}��/���m��7VLP`�<�_m���=��F|RI�0��`K�M	�c��ΨGQG)�y��3����?�y��"-i�k�ô��1`����B2���9i=v���>9���h��PMm����$ 4��+�^���<�j�z[dM*)��J(N�u��Z0��-#$૳+�m�__6(��$2���V:s�V"�b#r��V�|]5���TN��#	�L�"��N�������.}��qZ�pN�f������Raz�G�	��s����JW�ꋉ��l*i��)$�_/� Q��L�m��`��ÿ_be��T����y״�`<��x(�AK���jD��R�Ԝ�z�ҵ�R��ov���++-���g\Q���i�ϑ�f��6AU�4kv<9����f((ZB�߰�i��r�}�?V>5QE�%2��`�9�,���J����3�;�Zy�.!$ ������������6�K�zK�J\v�h>��;�ه���r�A�v��
=����OICQ�6 kz��x��ӤB
Iwk�px8a�(4]F+�
K����~�-�a,�u�v�W�B��0Qh4�2�ñ� �]��@���=�h��Y�X�#�� �#|�*��l��E�Ol���rk�����S�����$���7 ����A_gۼ��J43��̷��y+��-¶|�Z/���2o9�|P���s�x�v��6�[�m*м8��ʔw��pGX�S�T  jrU���g����g&�jP�&34ӆha�y}���Ʈ%���" �,�(�Z��"W�q�_�H���)W���Ʉ΀pP ���L�6���]�^���\��%4�Ý�:���6,|b�^X½�n+�ߑ`�;��M�5���6�3���0>�k��QP�,�xh'k�|9?�W��T_;��M ?B���z���B|��7q_���R�o^��@����F��]Oy���0K��ʨf)c"��j��h���_�\.�a������0
���Հ�LK;��,ߣ�l�px��������l���!
�ϕj7%��i���,��:&��᧘�3{��On����2Ac��L�V��-�JyU1�^��1s���ں�h�A������DK`t)�Ό���
��@$��\!�k�kD������$c�}��a�9�Ҭ7��Q��'�d��k�Cq���]a#с�<�8�(���^1W-��FՐ�+ &��Ǻ���e�H�!-����kO�'KN�(A�I1yS��f-��l�w�k(�";���}�0ރ#�$/(G�J%ݴ�����Mo��1��S�/���Q?-PT��j2v|�.}��96���(�W:��h��+Y7<����^1�*\:�~�P1x
HB��cif�+J�̵&�H�q���x���h 8\ ~G���/+��C��C0�˕\T �W�4@�Q�ˑp�3���wpY_�x��|5����]jk�� W���������P�UB�A.�%�Y��*C=^j�����(R�t��-#�1�Fc��J\�V<����T����j��	{��9�]#EĜ3^K;($�ْ�Z�����+�C>Ɉm��t�f�t�p�m��MԔ�$������eR����<��c���87�(�w#��o�oJ娘���1[�юIRY�M*�����F�0�w8��a��j�G��Y��w^��>���߁s���ȷ~�
�r�}NR"G�^P	8�|�Č��R�����Gڵ<�w�PWZj8<��W�?�X꺧�T�Z3��k8�u��D�kt�DʏS��e�^(��(�p�$4C�4#�h����J|V7����0�˾��^V+��Օ����)��/#�9&�bPg��	J�GaY����pL���]�Cm�qf!2����$X��[��u˖��������k�0L��G\)d4R
�j��fXa��=�\��i�u&R�X���6�\�0�4��&�E��_�b	�="��F �z�v����OءC��]�uws�u,�XϨY��d��Ӱ�����˭�U�~�@8C�T۳[f��y�F9��[6�4�qԳ���><2�`	h���j�C8ན^#4&k����D��#JV�L�ec)r�8D����_��:�Ɨs�_S͸4�!.��=�~�j��@u��=ޏ��DF�1��5��GD��W�>��_��0](������#��sL�����?����I~|EL>���^��[!+Z��a�j�[����e{z!�N�k怫����uWL�t�����2'������v[YY����HQ�z�W++nUEpc`+�#F���~�b �u����8{uPg>�WC�cHC�������ko����ۙd�5M6��w���sh��o��[���{a��J�hX���H���J�b��	D$@�g9�Y[�=u��A�s9=u�q�$��
��0�Tt���L[%��,�%�w�k�7*5֢����9B���iyu�GO�JG�
7���&4��O��u�'��IV;��Մ}�*�|q�xaG�(��9H��!�,��k��H�b�:s��Ηp��3tUC؛�Y��Ku��L�]��.��D����)ܷ�c��!��@_���*?>Z�ȭ,�	^�HW�gW�����(��0"�/�.�,�P�rU�!�W�ծl�ʒr�Y"�Mf*�o�-��Sm�����K�>+L�tϧY��Q��n'�U�$�['b�[LX������_��tJ՗S�Km�L`?��z3�B9�ف�F	�"O�-���6��*)�a��%X�Ĳ���(�-�(yK�\,��/q�6?u7s|sE�:�JY5��cR�(�"RU�y2Σ��
���h�ܭ0�{���JAY�t sI3�?|8� :}����Pu�|�]�>h͇�J&��Q�{�6(W�$|���y��f�Yڪ&�s���	�@�@����9{�qΫ�wԲ���w˱�޼��DY(\S��N�\�����.��Z�В��X�|�Â��{�`�[6Ş x���S[w0�ݙ�"6�(��g���VnAp_8����ß�78G&�gISX��͎6cmְXN�]���u���H�-��w��
�_�y�x-G�ɧ���Y{������ �����a��Z���TM��*~=��M_��'+�6���U� ����S��?��_��Yq�!c�ToF:M>ąc�%�x7�`s>�ώ�~���a1��hkH1ΙN1���V/��R��/0ڈ�	,�*�n���R�jZ�.3�U�.��Ϭ ���!D��1��EO���+�&�OQ�]bh��x� ��pN�T�jq��)��>1�Ȓ;�i�~B0��힘�_P	�̷z/̑��.%)�qH�<&��DT�թE��]�� @ڣ&^/��?v�	�y�%�����̶������+��g8ήjQ���XQPL��K!�M�嫶}R��D�{)?p��NF�6N�z3���B;�c)�3������A�% �!� ,0E�m�F������T�~�M�y��k�候�I(7T/���~�ݚ��R�ދ��M�|{�e�3)~׍˜#�n@����C�<��1�Py�.D�ڱ! ��D*���4��u._�@[����D�����:��{=�lU�=�(ϋ%n����[��է���P|H����zܷC|p[�y�i���'dW3�I��K��F�~=}�	�p��A�	>�����nU^O�� ^(;�0��|HP�o78{�Ю$5�B�X�u!�C[5��v�*ߐe;�bo�^��2�Y�j�;ǻ'@���2X!�=%�����BV�U�4k���s��仗�3�5��3���� v�~����>F�9�D:
�+P�I\�֝��A\�xIp�@�߽���B� m_�pv�? O0 �I��(=X'���쩔��d��i��-��<ł������!6R�]}*sF�-X9��ӭU�/�*>�R�~#�-�h�������6��VHk\��\��/�`�X�O��_"�'��	��'0P�.��А�&�u�^��bj�� h�B���U�V�����&//z�"v5����ؗ�N��8x^k�"@�|�c�M�k<~;�J)L�W���ۂ
6`<`��N�!N�e�m���6�](��{O����y
���j������� ���=�V��q����<Sp,;E�J�tD�Ҕ?P����n�&�4�Y�"P��6��M�༇�|�{$v�OvLB�hJw������G�����p=Z�5��	�rM��+��6����l2} �Jxj^S����yQ^f���ǲ"���3,F�-���ABj���?���Xx��ؿ~�c�i���sR2!K/|Endr�[�L�0�9���b\�3��L�s��ƏZ	����}(�eU�b�K�->��Nq��Q�	���P%J�v���)�N�W�s-z��������%ٴ�V��-K�BI ���Ѹ�t~����(LMr��#�B��ǐ�sd����c*����.A�a��{�KC ���v�U�����%8�����8�A�?�H1-�-Ut�xA���-��GI6�a���y<aˆ�V�=� �"[�[�׺x5�{�$�fk���g�|�7�d�Go��O���{vQ�M����	m��Aq�;��E;o~�:E|t����U�/������:��Gx�p%T���*}��I\��<�3��[7*�?��=(���f�3�����R�l�H��/�[W�t�����4�dF2ʼ����v�ŏ]W��ݟ.�B�7"^��C��謬�����iٔ�g�<�6�G�A��w_}�Z�&u��a�{��.�y�r�`_��vR'�{���Bx�7(@� ��;�hrP��H�Ǯ�Ŷ����	��{?���+0,��v �⛽�Խ��LsW�7�b�R"�l�ܓ*i,����̠��W� �*�Ǳ��Ut���'�o$^��.��+l&��AƎ�'&�atj�v�1w1�5�e�A�P���:��O�������u�#᥉������;S��?��K��ۏ���328��0��
�+W�x�Ym{�a�չ�/���,�Ѭك0�>�
;��[�ghj>�Kr'ǆJb�~9h`zz�?�� C��q{����DF��N���?�[��}	t��f�����Ӓ�<���K���.�_[:���E&���5̌'U�i�vy~A}�<~++x�x��n|��-m�&���kѢ�]!���#�m~U��SF�'����R�[:��y�"�������*(����S�C��ٜ��)`R'�MD��u�z7L«��YCx��I)bSTu�O��-e-l�6�P�28½�o�? z�!�=�k����q�£���xt�I�H@������$�a�g�ƚP���;L"�.�!�yqJX(=��j�tZ*����1���E�0 ��[��G�����_�"�R�- &�����Ѡ(�;Qy����^|������DR���JI�}�ì��,�������1��<���4bk����8e�b[����a)f�#��8�S��p'1�ÓY��	q*�a/+����pЧTh��B�7�� �Y�X�9ڹG'�廰��e�}�8����Ho��R���uJ�,\���nU�������i,x�u�\Io:�C�5'�g��������})��0�9 ����#��:�Kk�z�����y��f;b�����{8��:a=������|�|��&��X���;햜+~�*�������p=��Sǯ"�E���^Y�Ey\��=�	S�K��;ni�?��?��1J�6F�����kS���ւ�}_��#?X*��a��Cd0�����{���D:�/p��Rm��N[����m��5#�3�"��צ���FN�6���`6.�����c����~����4*��(~�cIl���@�g�� 4�R� ��ڧ�>��&k��Z\5���R�����FM`Gz��*Q�J�2�-�����kEe𹮳��K�S�����@  ��v�sr[�VuI�:�$diܼY�U��-�PSR�K�4=e�O^�����/� �5�ԓq�$�*R�$��5H;C�Iѹ|C���܌�@M-�:��uy��|��|�Di�[��9�n��n��p��=~���m���2�Ư��[�Q�`�|7�ˬ#b)���O��d̸�8I��8gy��UzwV.R)d��M�G;~�UP������Tn��dݎ��g�h���٧!M� z�3��d�⓽���!�D2*����Ѳ�l���,�����h�ĺXac �'D]�g��/X�܆똔�z��t)��ͽ��HsRX��\�� ������ �P\; ��]H�PQ9/bp8"aǾXK0��㨀���m��M?��n�P�c���