��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�_���v��	����}���g�GH����U�K��*Ѓ�!N�=�Bb��w�����9���\&u8�gM
���&@z��k�t�Ļ_xaI5�~�z�07��L��z�	T;Y�Q��ڱ�r��>~�}a�A�(��@��W�zW�*إ!UNB��nOY�3k�W�2� ~�0KJ����r��$!OoKg��?�ǃ���Vs_�T�+,����,��>�����M`A7N��;5�#'@�5yj�.�ؗ�pI���%�9�&�G[�������F�k��=Uk�԰���J��~����,��܀Q��a�KoE�	 ��"��.pE��]�M�q]#3���V�թ�/p����<2[�+����),���ԓ7r�̸� <��x�2����f�b!�[,�'�3*�˖u��	�#Ȫ.`�y��t1?-��A`r����+�ɝ2?B]g��3��3���|DkH�~��M�tџ�qR/M7B��'���T]����ﶬ��S�ӧ#�tt��naLY��Zi_h��5�-'F�w9�^����" �|Mڥ=np��}.t�q���N8u�����p��m�Hǋ�D��������ê���+Ţ�Ø(.���������n���r�����:� ���Vg*�1�-����?}ဃ-���AG�!�r��M��IҜb�ǔU�"ڥ�$����h��q�Q��No��;i�[�@x�}��g��z}�ރ��ԋ����"z��b���v����ғ�>'�xGGb&6�;!�>�"?v٬�eз�*�1�b��a�]!TĀ���?%f���:_�^�nKPOغ;�˺�/Ӫ�����6�:�D�A�Sjb�as�빢Q_cy��_j^>�(F����)��N?z$܅�������r�8�Tz�~�Dݳ��sx�Opw哠Ćm������{l��ʉ�9��XA$�Z����͟�l�'����>�3�j�H�pܱ8|�j�!�C���#���e<�i\a=��sr�HK��5r�b�\� ���U\ _"�.�*�>�p��$���? ޏÍZ�(h�1"�1<����g�A,���w�9!F����9/A��6��������V;�yw�֫�$�TԮd,hH"����D��	Ƅ~�g}ձ��sqQ<�}�I�e��{���fW_�WWP�1-�X�,���?�=�M~d�оW��j�����M�y���:c������q��ve֫�1�
8^p0��Հ������3��0Y��=(*����>#��������m��:U���>�hg�'��=F�0�F�I$D�T*��/pQ�������g��E�
��\Х�H�r,�;��n!�d�����%pO�w)�=$����"��+|a	���>�ˠ�U���NR�Ȁ>�ٮ9���1h��#R"?�m: �[��_x�}޳Dk�:{�ن���2�����z˾U�
y��>�B�vc-��
fO���Pj�:��E���:�n�#�x�+�$(����<V�W�PP/�*�����}�/�5��C�w�7��!j4;�h���N&�7�:~�3B3�t#^z���L�qO�kۗ�A�/�s������}�����C��/X��� }6n�E2l�(�&YO��
u�U\td�EG��v�Iy��/�<<œ���`�nŶ�b�+��o=��qe���<G��"VƳH����<A��T�,�V��˂#��*���Nԏ��1�+���[�4.��F�m��~�X|�:� x�Ґ`��ʶ2�}������(�M�ي���m��EcY�(d��:E��F�ZWdmbX$�G��~�]�Oj&��$�{��9���wK�9��q�"Nޜʺ80�@��rM��=�(�%��b�ī;P�w8I3~ʷ�#�[Wk5ٷ>��w6Pbb�ou2��Ob]J����,g�|[ \�?k���L��1NK]�Z�#�h�˸�I��举�N�9�[xZ���l|�m=i�|y���+R(n�J2�y=������^@�j,��3��]Tw���n��%m(K7G0�M)��	7�ڤO���)�w����J���L�������GaDy-Bs�dunA>��l�`�KG����w�V�P#�\ٳ ᒦ�?aI��ګ�-�ǡ�"I4C)ا�qS���(�n��n6���ת�����ӂ����z1�A)���P�=�Tʁ�C"��젘����GW����_�x}!�$5����(��4��-L:�ؒ{�}v	}��p��:�l����$X����C�����a�!�����6�Jܜ�sR#��}��\jƆ�r�8�8Wٖ�I�1�`#��Q�Pظ|�4�������cGb����e���+��Y�L���n���eX��k�Eܶ�/N3��&�vZ�fj��F���s�ǂ�Z���U�]�	�i�v�����0eF����U�PU�jgH�OJ=�=�M�|����,�/P�����w[�Jv��_1�+=_�o��v��D���R��lB�� $<#-3YX��I@�7y<��"�6���9��C�
Oz{���c��ȲoF�O)��jaW�e����a��\j���kM�P�2��$�C�Ml��^�~��b�]�j8��PY��Qާ�j�EZ
w�ǓC����v��(�Yf��K2��D嬧�W:F|�8ŗ��Ki�x���Dy�3�%D�ǕDo-����oU��[K� ��>��y�aP跣�v+ZW��GCph�j��-V�K;��\8ٶ�+v�_|����-V�`��}�A�z������E�%�Ȥ��\T�ؼ� �'�
ub�T�@���-���U��q��;�O������0^��%��M.B��{�9��aʌfu��������4�$����될�W^
&��)6����Y�B%��,c�%$�����\玜�<�O�B������N���^�0%`�}d�j�����&U���H�^&�j��w�̆���ӱ��� H�j	�a��Rj�m7@��^0��&�6%<�U$�-�������V�W�C+B��A�EW�ᷖ!�����|��9a1��W�J}�A�0�����8v[�����?���8�����q��!h�u���8Px��x9�'����Kf�=�3��d�2W��5D����{�N;t�wOq����Y�#;Qu��*�>�bQ �QQ��ȸ�����ns��T�̘�x֣5�k�$f��^�q	V�;듖���ŁyG`2t|.8���ig��}ks��5 �-�̓r�@�R�n�C���{�d��Q�c@�ep�{Z�u�����dW�c����CЏ��R6RD��8�'�JG
�c>��F�Hǫ��%�����sfQr5�^]-��F��Q'�b�Wp���M^ʢ�.[/�k[CgalF|7P���QadZ{� ����*^Y�謞�T���Y5���hjΆ+�����'b�8���je>*��oA/O������d��4ےU#�wc���?O��^{V
��e�[��t?2�� ��Y�|
>'�%��wEj#�Q0kN9���u�0Mt�ɇ� ѷ�Y�$��Y���q#w�Yl	,%_K��T���1N ͱ��u��E�J��F���(i��9axqIۜ�݅����'��7�[��G�����w��a�q��ܪn ����������L�[:>�;�L_�g����3UP��i#��6-��L]���7
/���q��R�k�6?�b p��/t���#��_�ݾN���T#�BR8��$d!1�����2O�d�D n�k�A��iRdͨm�w!v��WO'�#�.Y3Y�=��inӟ�������<��Ŕ�jzj|�ߠ3��62�c>r�Hh��}�������7Wq}�8`��W�o!�Z*�*ĶM*�u'����_��^B�j�?
�ݙD~ez��_�y�f
 G�%�*��hR��vl��!;��ب��^�����;_�yK�}RZ�"����QyƇ	ٵd/]Å��]Oq���m&Pzߧ��+I9�$v>���<�W��m*+�[[�,��wjEu�(<����-lؒ8��`���q�1��:�hr��^n��6�.=0OM�8<�}�
s�1��#��7g�wudQ��nJ�ه6���S����r$�f�'��j�z��F~��2����d\T��?�f�?���(+�#��"�t�g��̓c �+�勺b *��uM=:tS���y�嘬G�~�W1�:
�[���KËG�
%�A6W׼�p�@�@=�+�?�l:�1�����N����/k��&X>��4����EbP �$�bh��ப]�	������{�S��ƴR?"Epy����W� k���!(��7����K��#>�݆��ۣ�T���	���l���ʾ���u�S�p�J��2*�'�Uȱr�W"�A�z_ɓ��64��ؑ�}��2�������Y�3�vG����Wa����&��Q=��*�pޠ<�I�ɥ�����H��C�����atڢ��k�V��m�8��$�ld���]����&��$k�'�XY��Ѵ��n7y���,a���UQ{��@���u��([���g�.��ׄ����14?��#C��W/�@2�k��g�㚜� �}����#�:������>�_R, �������8����ɲƗ�,v�BR�Kx����m�YZ脌%F|_���0<�;���"�K��%d���hv~��,;��_��L��� �lJ�,�&���&e��莝*/��@+�� &�&ݴ�}$�O�7~�Σ6�I���b��3B�O3�̨�!0aE�T���+��6iLli���� Dp���onA��9��H�23�?T)7$z���lj����{����V`���f�+{>@:u%;1,�4�Bԭ�BYx�N��,NC�2�ߛYzҤ���2���Q��(#r�,{��\���<� �@�[���4V�!��}�Em��@̂���J5�I�<һ��| !�r��,�J_�L�8c�euE%�z��w�>זr���Mp�C�YNY��b�c����|q��Dr�Ɲ�k����R,�X�U����yRcn౭?bp� q�F˯�+�3�J�@؎Q6)X�AEx�v�gg5�.��7���p�ֹG�p�ۇ�$N�G�PR9؜��f�C�����w�ɘ�n�\&���Z�����v�L�8��w���No����}bK���t�(}�9�����\*��9y$�����O�|�H�:�<���	q4���|��!-����ř��l���Q����Yܬl=�:�
�_b향�\Y>���`�NF�!'8��O��K��������ڔ��/BkN̈́?�9R����I;�|<�������h�6!�>����n>���ȼTw⢾=!4ZeU���f�Q�89��V-��H�Ei��dG��)Xy\�MƳ����N�^S�(���*p`{|]?�|�o�.!)̓�N�u�A�I�c�M��O�*Pܹl4���c�Y��O��!���5 �U6���wK���%��M;�ZA�EZa���y͙�����A QH��u��HK1��G�Rf���������e�����;�!K��˝�"��B��{��]����(�\�CRR����L���:�@;t�H)D�A��r�	�����ZGGyĆf�&ʦ� GU���u#4���1�Rb��I���Z3���Im��˕\L��Jp�s�̞�H6T��htJ�W��sQuY��[[՚�}ϗR���'ֺ�ݞ�h5Oܣ�=D�k`�(j2.4��_&ꥎg�J�ZG�\�����p�\R�w�n���ǈ^
pAs?pz\��ἡs��N�R�teG~;�5:�"��۽R���,u��+��v�y|�&�d�]2��Xn�c�P`�c�QY���2z��!�:�8H!��W�/��Ƙ��_��WUܕL����x{�]kQ��֋���aV�pt��w��k{�?�wS�%�9_V��SU�[g�7�r�<�f��k�Rsx��ԑ$͚���6�?�i�!ԃE�vE�S
J�G�wy�����ɱ:���o���r�K��yI��bݩ]�����[�󊚁�`�&�ֵ�鄽 Z�כ�-���L�O^�F�nl2�=�H����绱�yU�*]����JϨ��UV��-���XF	=���/Q�G������Q�x^�[����Ԡ�����wM�˽��w� ��*D�7>A�82�6 �$n�x��֮�*)�5��geB�����P6�|�K�o�"Ȕ�V)����+;�Q�b镶��}��7��P%��iHa}X�{o�Ai�Ɍnm�񹘢�\
���PWb%Qנ�5��^�P�3�5��>�N���C>��*��aFW��O:�p�/l'2�o�j�]�[�dB*�n�f�VOX2@����n����9�i�H�Ћ��V��8�%��7q��TL�kQc'����]/���H�3�-*y5���)m���n�]|��{u5�3�H��B��L ܥ�4K{�m�#����?��9P�/������r6�1���z�y��
�By��_�v#�
ה���\�ZŃ�R햃��Ro=y�e�`�n�5�H�@�]�|"R�,��_v��J���dZ�{�44V^h�Z�Ƴ	η�}����*s�?-�'���c�?��8��I)~r�4��|ߗ��2�nD�2Zl�+��]DW����j���cଐ9+)<+��O�)	pȗ v��]ʍH�δ��:	(�
�.�o9A��<VۯF�@q��
��[��[ 	2�s��ը?�6�7�|��w��X[Q��ލ���;:XU3Q�0N��L�-�Y����ם��.P����a1Y��i��chm�RF��d� z�Dsyf�S�R��M�B��9��q�6����}�8,^�����C��o�n3ݟE퉺��"|�dzf8[U��n�Vz��k�'�å�
'��^���.j�֭|P�5E٥�E[pv�#�F"I�G~��
>a1X3��<��<
�!�Y������vϳw<S��wtQi`�.����F!���.��򣤦K0ɻ��ôOr�M ��Љ''m�ơ�BY�c�L�qE	-�	��d�ضh�|��P���X��u�MA>�ω�;��tS�N0��^.�_>:۪�ǵ`!xJI�P��Bi��G:��q9��v}r/�DK&%;T�_��R�	sBx#����X���-#������ �`�~0������|z����2��K�~��ڿvJ�`��g��]��åe��Vl*��;��_�]�?6����"��2��WݥK��н��s
!��� �Y|������ܒ��s��P�^�wH�������RiѾs6�t�t�̀��n|��jb~�M�`B�X6"�X5u�_��~��ִ������ {ޔ^�+�h�ƌ�Zc`���Y($R��)��P�%���v�[���b�4��=�P~�;�����(Y�?\���N���.��%i(S��<<����	X��n^�6��I�A쑑)v��~M����
cmU���[�H��;'}�V����e�G6.���w���T�qv��]zm?�4V�j9�@0�^1�A6䗂�//v��:���S��[��R�~��3d!���&��`�m��.|����,c�Rx�E�3 ��p�ea���ad��>��50�����I���v�r^p'k���=D�X������v�P�a5rtda��M����ĒL1R�j�Z�˽�oVU�6+H�tW=� B�Vx($zd[� ���A���X��W� @��@o�lz���0����B�r�1GKcGa]��S)�lZ����^$�D=/��s�ջ*C�D�4��J�D�ؘ#M�H� ~�@ g1\��X��|9����R?�V�ofgU��c��Z`��-7���~���4k���/��J�%x-P��%�5�fš���
3�=��doS8K�o����lͿD:RbU��֬`���[�\�l�V�0ѱ ��풎����)J6y@`Z��`4�i�$�y������?e��� O��=�V�7Z��'O�+E ��@�BIb&c��#s�7$�Ӆ���'�1/�&{�Y�D�n@ܶT��.���!f����ʁ'���YX�+�%*��9�t��if.@]��������>���P���s��W*eOY��*��YVT8��}��3�E����O! 
�;��p�������(�4kh:���~'��9��+��> �T�˭��C���hS�d2��^�+��? �{����xi̓����^�0��v/9�\)~m�J˖{�>G�,�3X�gF�O&A��.Y%/�i�d�^ ���ɂ�M0�M'�-X� �9��e����@d|9��x٦�^:�y,C��ज़�CN�x`є�;����d�Tz�%!|�*���P ���J���U�V��}y|��UƬ����i���A�#�� )�3gV�ƢE�+$��P2�籦߿��j� "{����}�u���V&���ՏE�y`���O��0��r�G@���g��Ep�cΡQ�ZF���ɋ�[6�O%��"QS%Zԫ�ջ��tR7O�Ei����@�á"tT6
�8�1�|�[�]�0S���|������8�b$���;˶�܇M12�=�$�P�1�p���o�LqX�:��`0�{�P�=��b=��.�]%)Ku¸�6�S G\���F��=1�z2`��xk��0&Q8SSotʹ���Yc�D���
����x$q*,0zL�q���%�v�Pҩ�&"I�VC{1����Ԍ<��Xs3V�Sw'cN	J��/|<����H[�81­��z��c��6���ӽ{f7ٌ`h�ƻ���O{,���J�-$�g�՜i���ܹν�B�2�&��<��~Z�L�^���Α���<���P��R&z��g��;>�ni�CR�s� #?(�L	�6B3CG���ĕ�eMZ���s�S ���RN3ca5�t������U̞����h԰������,l6��%�2Í�	����9_���:L���=r��r�?,s蟩�+@��C(��Q�8�hW�gXL��
KN��o��4!�u��Ĺ40��҆:>�;&������%})f��pTK�M"��^Z���1,�p>��{�ԾމA	B�#��"� ]�����?�/�!�a�'�Me�_�	��#T7Z뒪�W�<R0����m��n���XK���zQ�]�c�mC��e���C߰���;���o���z�E�`c��4<��?#��@Hh��-�w�Բ�Y@�	� �Iɤ�\s,2dnoᄯtW�eI�*w��s�`�8]+HڲL�؜f�H�#�Ί�/�	�V���آ̖�1���ݾ��|;�_�jiyS��N4�t-�N�@i�@������\����H7����@\���4�
�6w �KN/�Ｑ�-4ʜ�����������\�sm��[9����F�r&�#L7�q�*���뎌0T[���$�����IҶ"��Τ�Ҫ�q��\��C�P��&�_�R�Pe2[��_�帲xe��J�'�2��x&�[#s��H_�G��{�r�t�*L�,���T���H;U=���eG�fc��T�⒵��в�o
�9�Y�0maȅ�%����)��7���B+'wE`:>mF����ï�L�󝹰�'=_ۂ?����g�s��	�EWa���q2�"�����ެ�;����P�
���X��AI��X�qR� u�k�uQM!b L7���?�ː�Ũm���AUj���:��Y�b��@�<c�|����J�����2_h�t��R(<M��
2�](�n�E�>��ܐ��F�� %Ɗ��:`��C�wm�U��
GT��1��p�tC�ц����5#:QZ6��d�hWn���x�����7�hj�Ї�2d�G<I �H��
��4q����{���ک.Ľ�J�����$$��F"�׍�b4S���Gr���!�)A�t�9���q\gZ�+��,��1� 
9YA;���P�T �.��7-�'E@)١�-��K��������_�!6-J@����(��S|Ψ��#T�6�kD�o@/t8�ݷ�L�t �H���丹y~��5G�ױк(�
7R��x���R��p@����s2�@H��'������.�7]��DO`h��v}L>mu���djJ�V�;��h�����'e�<.2ks_m��}^�E���|�U6�a�~�E�p����!��%پ\=;���삸��=�p����#����:keF�L�*�_�����"+�v��Y�J�	N',�l'�	�2k������ �t�ƋE�W7�祦@p�aC'1�JWL�����ڏaǨb�B`d��x�ີ�2�j��(fDrKx���m�?~&�G���B}#�Z�Ҕ���c*b�'PB[n�f����@@{�����0l�u����]O}�-i��O�m�#Q��Z.Q�&d�Q��P��6}P�XX�L&æǰ�t
	��	O,��a�\_��l�b��v��t;��sd�c�J�mt�a"�LpX��s?�Mr�U0+���|��+ ��4��L?��4MY	{�`�%+����"���|<�,�S�X�H	S�8��(�ƩECΏ�d;�VD�ځZ�uMZ=��{�8e��}G%p�+Y�ػeT�ٳG���d�ϸ��ZL9�!��s�6��	�h#8%���I�¬�����0p3�.DV�����XO� 
4#��#�����t��~.����pj�|HW|B/�(H�:U���фI�� �ty�M񚍗+-���g�9�����S�.�D$"���#�:�޾��2�;O�&R����L�$�_H�H݅���&���gLh�/�Fn���E��l�j|^"��s�����^�b|j��
MC'�Y2Ř�{�[��:k�a�7�$��A7?�5�DS��پ�*P���u)ta�GSt����j����"����]"�腑ܾ\���0��Z�L�G����uި���6��#��[�#��4z��0S�!����q��K�A !���m�($���]Vz��"?���Gq�;7E����Ugb�ku��u�''z�T�߫@���P�s�uR��o�2�fi$���ם�s��c��:�]7$��m"�8]�S��L��?�0wJ��0��'~��&Q�P�Do;��w�,1��[&�5�޹�8!5ܷ�#?T]��t&k	!�^[T_ݵ�ޥA��CV)7wOOC�PTz$�����˃y�h��/3{�Z��Y7H�K0������Me�p�ѓ��ڜ]f}k_�6E�1��HEPm���6w3�<b�� �h�PaqS�o�NcN'ʽ��k�Ì�"(�41�-�4��( �[�]*��_Q~L���9�a9�P�u��Q�Z�� ;2lUܨ�A>��d�~ wk2M��2ť4��n*�ը~.å�wϒ��Ud݇���FS���2N��������w;�^bj�;vpayana��Q���ͽֽw%24p�m�*g��S�5����gl0H�Cﵒ��
 f�A�=i�4�|S?	%+��>���߬�n4�M����LQ�f�b�9����\`�N��Mc�.�?�­����-���.L��/8�A��v}���\/�@�#q:�OP�k��3_�(��S۽��T��~�eJT~��pJ3f#l�I!���{��}[6t�F쟑4�� %?��ar[M��So��qS鳨N�$�,��C/S���<9pǨ�����$�����Q���qa���ʰ�u�����6A�8%�@��Dk�ȃ�s;՞xeB8^�v�	.�OU�i�N��q1]PvϑM�~��a�o�=|}<����
0�b$
����τ'$M/.�ێ\�։���ސR�<�W�O� �l�^%�Ǫ�M�8I�4[T5���� �ڗ��
7�~�a�*2-g���ԇe:c�~ -W(-d�^�
|�ޚ�ܼA?"�O���I��ˀ�Mt�Y_Ư/���`r8��m��qnͼ��w�Uh#��"6�k7(�z/�����q<�z��6@�uvy�(k�+p7�E��E���[zuiՕ���՟-W�ՠn�j�zc������*N��<�d��¼���I��%̽�Wp\G����f����,�y��cv/���g�pR�:��~R/w�.'���B�f�]�癮#S�o{^�;�����)�N�"F�:T~���ğWj
����2;E��U� �.{@�H��pQ�%���Z�s8���2�s�}��|��'PfIi/2��J�ё�X�}�LY���Mb)��v�)Y�c�G�:(B�Fiš$:�
��#S��*P�U8�6�Z�������(���c/q%���Mگo	� �{R����$��'�?ӿ/aQ��D��ՙ��}M֘%S��C�b �x�����1�~'4�t2p�j�~�Z_ ���e!-�}w���-XmV�xg74�)�5J��#Vnt�s�g��I��`����@����aƃy�"Od�
r�����Q�D�O'�����~#��d��xt����~��񌦻W���U�`S�R�M�]����0������c�1|cpg1f�� sw��&W�� �J5���H����z})60����x��F��ă��ng@_u#!-
b�Ǳ�]}e@~q��Z��~m.�Y�O���ip`���������������Hw$MiǬ@���T��YL8,�V���8M%��Q�^��n:��IZ��l�o�V0ٺ/q�p�J �~ŋ�G��Z�nZ����>�H�kz�?{��>�_��GG���Z�5�B-��ϔ����j;����~�?'[l����"$\	-�8n�G��_=�����r$�E�N)���$��;7�"�4��
qJ��0ٖ 㶻��[���������0>W�����44=M�^��QԘ�0uЏz�y^�:W�'Y|tu�퀉`(��w6�D�R�Pf*�%bʕ�U?V�Ŧ70��g�LX0����V�U6����I�Rq�+�9u��N �$�� OZ��M�<�QT/~,*JV��䥚��v�*X�V��;����0&�m�K�E�y@���V}}z�h�ҕB�|~h\�ݻN�Ʌ@�:z�K�:���x����7�'��!)º�e�֦����r��auP�ԔA�C���c�kǓF�j�vG�cb���7�������ۭ���.�fN
�QGz���sy]�Omi+��{� ��8���kt/%xН@#���%=�Hn����`o�u�,Y�_^%�=X]�oSy8���>�.��b>8M�x�Hg&?x��Ѯy�$��\�W���ԩ��R|Ve'��F�q��Ϯ�T�%�$�/ob=0d�p�S���~�zvѮ"t��|�u�4�K6��\��תI��=�rU�؜5<�aiJ<|���z�6�(���m���7����/���������3�o4P����5D9O��:(��������N4����CL�"���o�~9Os�l桨v�i��7�,�Ɇ�B/�ޕE1U�j��V�L���:>��~���ņoҲW�Eϝo�
yƙYI^���P���"�-]�q�Q;�CQG>s�W��^����W������씉EC|���ھ݁s�.��ju���`�	P���� �|E��AS5�h$y���/cW��r����Y^�g��(R��cr}�t�N�c�8�*0K��;l���r�)m�CO{չF�b��У�!�w��0��/'�6ɜn�T뙐������>7�8�[c���#}��d�sU�#���z`�X��k@�?�[����"A8V�+�"1������='<���Ś����L�aҝ�ʝx��X������^ U�$��#"�����1!&��9��A��==Sr��Lv��u|[�XՊ�T����q�RÝwD��u�
�f?����;����v���J���lX�]���q�2F���>M����"˻/�׽6��tX	����'}�e�/W�ք�C�_�@"�#-x��@�欓�@ޱM��e��\�����H�7�Lu
���#����᤹^]�֜���o���.C��>'ƻ��S��p]A���{�	)�/�4񿴫���T�svo��~z�E23��S�v J?���gl�&����7��ѩ\�ol�Y�j���*�rc)~n$I��	�Q�j�L��㒰���.����wM>��������򧗕�pb����5���S��̃`��mT�!��)�M��=�R��:fP&�����	��W>�U�����fa�P(�m{Z���f�;��$����J����n��:��*�i�P'e���9om�&k�v��(g�_��TJ�O���q�H>�x����Su�M����3����Q����!�B�>�
�4��̲�����d��Z���m���~3Z��M�3��n��b����f��E.\̦%�ec5i��f,��i���?eA�D��Mz�y����<qK�~��-?�>.��,lNg�S���5C���(�4䕐(�ӹ��S�A�p�+�MI�$/Ԃ6�!?�����ŇK��Uz{jy��3�V
ʷ��P���ayɫ� P���%%��'{�����8{��i�z~�|������/UX��޳s��R.�~�?���d�jm���NۛcF��3ol���'����<u�i4�Ԏ;��si,�>��d�	�6º���	J%e0��d����>�;�9aH=�=��PPT	1=���z�i� FT_�3G�0�	0��a��P��@�U�M4�t-g ����na�zL6A�R��"'p�-�v��Y��x�!B%Z�Q�J"LN��a�ѣѱ8b�l"�m�%�D�Z��ZA��p�F��p��2�a�����eĂ���*��ߤ�}�j�>�0��$7�"2�ϙ�����2��{}�R{u�y�0��H��a����[P�i����<����A���A����]������	4S����v�)6&l��M�xN�}Õ���~�����,�?�8��GP4,i� i�p÷��y�����-F�.sq�����u��gC�,Nj��_0R���^&�BB3�D9������-a�U~˼$���D�������9GC"S��u� ����)n=��jUc��m�5���2(��
��wb''Lc"�m(�#�4��^J�c~��mhY5Yfc��q̹�Z#~z&�t��9U�g�/7pԩ�^�WXy��#X�{װ񄗆��.psm=�������.�Ί������?9D�D��@��u"�;1�����_�"_:����>��44X��Ã>���� ��Rɣ�W[F�U�v�D�^&r���F*�z�?ȰNv4%4��[�kQ�e�w�<�v�1��ڔl���W�:Q�(�!�Ɯ)齟3��w#�\�	��Ez<��TL��t��5<�-#��	Nۻs�fݲ��\pTG��.3$����!�a�-
���IL385�bR8��'$�U�QQ��˦�CC���ሑ�C��n�w��r��Vb�kF�r݈����*O��|6��t^p�md�D�s�f5�{�S~~�dRzM��p�NP=T������d�
�M�{}C�1,JQ�u-�*/�u��6k�\�q%k&�ϔӻ�gn�I=���ۆ? a)���ĩ3��lݖQ[�^�}f��ZYTu�#���fz�'S��{�f��Rv�l��#�~�^�h���Ij�5�Y&��C���S�6@r�X�.}(x��������0)v3���:F,3uQ��3�fB��s(�/��)bm�W�~T��D�/��gp�"*��Ɛ�y�yOK�L�%�*W@g�&���or��
�g����X��1���A�J�������Ah�0w(E��B�����w�p5H�+�#���a�5�rV��8�qԣ�;1�KW�������bɃ��'7��߀h!C�7?8��r���q��ƉP���x[�;it�I0�N������x���W$�KQ���(̊f���^[��xd·iKic��B��N	(�r��7%����Ϭ�&\��y0P�-��">R�۪G'!��*�s��:O�;��bW�ά_� �e����x*�*��))�3�T��Vkt���oK@�h��WU&|B�� ��^�p��{B��YH��7�_T�uT{<�V3x�xj�`�{�ˬ�b�4���n�䊑sF��A��	k7|��o;B5���N@����EV���z���o���dNV��w�zK���-�S_�n�J9#chς*IGl���/\�P^L�]�f��K���a�BhC�xF<I�
(PW��7��?Ȫ��n^$�{PO�|@�k�ĉ���c�6�м��=�{I�.st���<?!�,��#�	O�#�����!G��.�=V��4G�>��)4�.Pc-z4(�;b��ϿY��⢤�j�q�V�����	h�~�����)D'���f��]E5?���W/�s:�ԯt��'Y�@�OU�p�|1@ۧ0�1��TѸv��
Eٿ݋�¼#]�t��g����R�;9]���F%�S�z�N�~��=jj���壣���t3������w^W�5f����a��ٯ`��8�+�;��i�w�GHaH��38\���Po#k��/C�})�
��r��ĺMI���)xO?	}��.�d0#�qjjd�DF޸D�+*V�iQ��s�&�����s�?��s���ur�^S�ot�ϯ�H��H���!�x��1Z^y���}���*u�7�fg�*��`.d�t]����[�:�:_��4�Ȋ�Uz�q�dK�諹��e��1!BDP���T���Qp�;j��,A$�;�0�M�K��֚\W2C2M��.��e��Ѓ��}Zg8��m��_o�A�+�/Di��ۼ�������>��م� p��n�tQս.V���������}!�y˪X'x&�}7����ܫ`��F=��N��]<��%?TʙW��	��
?��>*'�;&O�s�	{m��p�H�s+�=�����B�2�
Z֌�/�W/��
s��^����T��a0��Q�*|	*�&(^�Q��-5I����9')�^mÙ�L�MD1�X}��r���L=�vY+ ��#�Vh@�a�F�|���6M�b�I�3֖89�`9��
kN��r��<��se�5�Ȓ}�?$�A_���Ӻeb���;���V�6���T�"BU�
���i��~������v]�fJr�]6C�Ӛ$NTg�^�˵���{b��ޏ_�˿pʕ�Hx�p��e-�y�Z�ྶ��<n�����D&�Tr&.�w��k6��ZFH��>��� �r%#�<�/\�%�v�w,!�L�p��Φh��))M�����ܖVُ�be�X=+h�pm�#�R���Fv���(s�W��?� !U!ik��1l��W'���!�d��?�,�*��K{N?K�`�Rҽ����=�c�kj����t�� SI�cW6q�E4_�u��͗>���^Y^t�݉l����d��ɓ��7%l�۝)w��_���^�T����"��[�N��y���}R���P��U{�����$�sU��R�
fu�|"��q�f��?R�Cb�M;)��޴��������������0v	c�\i�� �%����@��Rr��\|_;�����H@���IêI�U��t�]�8�S)ݘ[��g>�7|\�{��OH�����D�T�Z]�MHS�@��o������O�"K��q����v_����e�&8�s&����r�	=c���6�s|`��j��b0�����%5mO�T��"��9U�:�%��0�`)��2�_�SC�"�P��[�%Z;�2��n5�#�58EIb���kb/��֓uCJ��}�ܠ��1���_m=b����t�s�����=<��7�0��"�"e5!���E��"H:$Ͷ�I>A=_���P�sc
!{!���X�����������hQڂb�eC�<WgU8�2���S��,��l��kDƤuD���Q l��\�".�򎤗�m{���`��eJ�:��2�����y4V%�M��[T����UF��3i�v���e���v��6^��9R@�*��H3N���q�0+{/g��R�*�8�4���,(JFvq�p���k���2D�&j���$R�]S2�c*<_�W��w+�O��Y��'z:k{h&k�B��j�p��>��ǅL�M�q�=oȻ�ۚ�7��tә�
և`�%�)�߂ѿ�MLm&VLQ�4�Jm���G"�!�_�����D���G���p���@�����*sV������G0�[V��௠�#y߆o�X�6���~��������>���bY�!��
�Ydc��j@��]�����������ͪ��=�~db�]����n��-���Ɔ�e�E�&ρu�ړ�����# \�6W��	=�:��P)���h�V�p��8�)�(��'�7���� �,k���؁[�uo;ă���*H����-E��>p�u�ȡ*isÎϕk���P��Mq����h��òҋ�a5��9�O忍��ř5��*�j^��WXHޣjn�S�d^�+���w΀�jU�Uf�8�ƺ��d����O�M	��"����d�Y_��v���$�����Cc�THv`
�tK��0x��,B�2蔵�L�%��jB�/�}�L���O,�כC�"�'��_d�,�d�eR��͚h3N��9s�iR�8�^!ф6���߽#G)�iM`�r�2��m ��p��kJ&T��Yn��Z���\��j���E�e��YR�H! �Aw_1P�{$��_�)[Q�d�����!�����K�e��r~{�,z
p���6l�QB�Ј�"�a�[_j�3��&ET�, �c�B��ʖ�V����:�.f�zWY�wxYfx�iNg��E�%q��]����M�ѣ^�	��[�<w@�
d(������ՁZ���W����U"���"��5#���W���H�S����U��3(��IÙ2L�;��>nn���Q�����H�*q(&N��䫂�A�2�yW3�u�����h
026�P@�eX���L�Gn6/���A���U+�c!��5��Z�q�;d���� ��)��ǒ=d��_��/y���8��[�d��i��Ň��ǘю~@��Ҽ���ܻ�8��XX���IGbg��2��+���!Z^�x��֯���U���k���AƯ��bF	�T���i'O d��@Y���2��߅3E��?��/{�Y�L�_ �]�zM��w�� �>`Jδ�uM�C+��1p��-u�0D���r��BG��Y�#{�=��<�X��n�}����7�G�r��z:����V�_m�v)�ɮ��ܝ�sEo��V�L-�]����3� ����_��R�� }#�<�Ҥ��6��e ��<O�f**0^1� h֪��ft@�$�ȠR��h�*��i���!�����ޏ�pP�^h���vy����#9_�~������z��Z�6;��e���y��d���KF̅�������Jk���\��)">K��4�'�kV��5���-�5 ���N���\��*��deؾ�q���|���0*�@]�\�SI#���b^��+�)��IO)�G�^�:T�W����z�P�L+��9Rō�7��3+�.^���rr%{��ʍ/>��å��Ҿ;�e@������r'*Kߏx1!YT�z1�znڻ�>������d���و��]���!�	)R�k�^E^]*fC�`@P{s�4�H�ktl+T�P�oJ�e�Q�3�,4\��/
�;�3��Wj���A�%�>m�Ae@����y#w�%2/�!���s_j���T(p�m��Wk4	��[P�G�=\��S9��i�=�Y�>����Iפݠ��Iό�M]I-aSY����o�[Ǯ�8*q�|,j�-�s{-&h9l [�eg����"l����������hv:�Ƌ2|��j�5C[���"��m`S���zf���Tn�