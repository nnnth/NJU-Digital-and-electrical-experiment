��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�E3�hoA�zFҿT���8BD���9T�'S ,��|�0KwƱϪ�g�d�FH�^w��#��`�}A�`xӑ����u�;�v ���
>L2��������{���ݕ�O7A)�R&��H�=$#jqZ�;]�稥�a�a؃��{�C�.��J[Q��I�	�b#j&(@��^��F\�Ԓ���H��"�B�n�CZv���[M~��A�ю�Z�ͥ&�������+q%��y�kT&ż|�����K'���I+����&���˯t�p)y��/�j���(��$��Kv�Y�c�4�K���)�"r怒��{E<���q8O}�����"�8���ӝ�az�$��5�B��֨}�ŀ������tb�N܊|4��%�*yҧd��YK��m���?���괋&S���:�˴���7/����	Q��ۀ������(#������!��A�B�h��y�O��ȭ�W�2�S�m�xa}�B߾&�p	���a��Z�=��sAӬkX����Y�Q���K����`w!𝔍č��'4�B&1FN��R��n9��2<����~��t��S�[[�v׺�0�@1���<_-@TȺr+ft�|r�o��:��6
F.T�&2��f�zn�O�#��gڪ�T�=��-�p�^��#S2Y��k��Z�*[4����%j7�ݬzݧ�r����0��+*@$�����%�g��
8�X���7�<�h�W�H߯�T�O��8�i[P�*��q0��N���(Aԋ�8���?#�����~��k�Z���}���q��,Y�Y,���D^��<�_&�C�-��VK���E�h���Ֆ�wXE���&�.��6_7H4�iO�-+��Wb�5��!�۟q��D�]Vh�IYޗ��:�n5L�����������WZ�}t��rt!s�����V��
����J��k�$���97p�Z���铚W�\X���UH;q�'��Qב����vو%�QŤ�z��W�|+�7w̄,�M�{�0����}�`u��-�p�E˘�������٤MUu�݊�n`$$\�����.a�*��~�Һk�j��"�� ;GL�d1C{���I�Ѧe<��zX��3�%hr����+|B��C�86 ������ �:C>U�N=��A�B�dot>7�O�Ҷ��Sk��$
7��Q�s�#ɢ:�5q3G�$�a:u�oَq��	 ����d@|L_l��'�́����ۜw�j�5��xT�,��c�0`vMr� �rA+���f�q���VЗ4V<r��^+�6pm [4��,»!�)�^|�u����Lx �5��2�A��`��}�s���s4����A���h����ChC�,��Qyct���JW9%����FF�p�u��076I���"�+��k�/���[_����:~ႝ��r�JFF!���rk0�꟡����5��"_텚m =��%zHX��o��(w�>�5�;�!�C(~	)@2����!,��=<~�j������h��L�0Ç��u!�(A#Ն3F��1L��m�V�>o�v0G�у1	��Z&�%�o	Nxv�ޛlpwȢ��焾�S�~�u����
o��6�M�[������ӟD$1�i�P�U��+����J;.����t�l��1�;z%7��	������t!K钉X����!
��d�&T�`j`��R �5�;�u�'�SG �W(���Lht��xLD3���q'��+�4��Y3���=g"�O�������F�S��4��v��d�w�p�e��E�w�T�?�������X*P�\Z*I'�*�S6�H%���!h׊Y���J�7uwV¨׉e��Mj�$e�xBDF y�^��*��)��}0�I0D������в6l��1R#�w�g����Ir����AT�CsQ���>Ob=�ϯ�8+,`��؂��'ܼ��l!��c-��Z��$�قDǦ��i&�����ЧXPy���#��-��
b�/���,�a�B��
���p����`_�' �zs>�͚u��j�i� 6������M�G��!gw��{�BwԚ/�],s��ȥN^?.=����5��u�U�zi�Xq1���$ �FV�Ewߦ+�Z�g$M�����l�	��Sh���ҟ�r࢛�c��$�i�\��HG����q���.r���#R1Jf���)+HΖ�-�ޓ&ug�.C��x��cP�����>҆/s��p��@+z�>3^��.����4���~����Nmc�M�IQ��/��{)�6�36{�f�.Mu�{�u�L2d�z��y���]����.B��&��n������f�����4\Յ��6n !Pf�o���_�JCj�)(��������}O�Z��p�˅6���:#�^u�8i�l�e-�;���J��oc;m�s��G���� �iH�}�j�5�/�io{���.j���� |0�Ar|����ȑ�~�ꙧ`2N
B�
4��_)��,��o�t�,;N��T��~�#G�L�r�� �&oi����;�Frq�a|���b���w?H��N��)��7��!�cE$��t��ayB�qS�����Cٿͭ^Q�\:t�[%����>��QX1,�Z��:�E��턾b9a>�`�[]�?[��Z�����p�fJĿB@��f� ��H�J�2����X"�r"��Y��n^��
}1�i����z��˕���$%�X��	�~��?6��6��E�A�&��OیL���[�thA�X��9�Rh�G��6ꌡ��3}���#1?�뱧�wqʸ�w��y�����E�{�Ղ�5����^�A�f��1���w���te�����4�κ��\*%���GQ���M:��&��{r7K�%��jO���&��ۨ쮀��ȫ���>t�G�qX���aJ^&\D3�c�\��3g࿁�@�u�j[�5�ID�3��,���	�3����/�tp��=O��Ȗ�֛�r[�*b��g'��#�f|���@��*�c.��������\�f|z�
\���R{�� L#J������ц��Œ������%'J `��M��1Nb�K@}C�8�bj��𫝯Rc�-�}�% ���cZi�,:<���.#{�h�{N�Rk�\��L'��+��v����B���%��Bܹ[t1>b�"Ȝ;���� ˀk���S����gd���T#a� i+s��q�~���LN7]M>�0�%��}KX���3�		aC��v
�;+�5�s��t�D_3.���T�G�g�'�|��������生8�C�����y�NZ��9&����js��zD��&HZ���Rh�Lkf��9r�?��F�1
�/zg3�s�Z�Z�C�KA�L�M��&_sJ�a��:��A'DyA �Q��i� �{��Uؖ��/����0���� #����b�?~��Sڻ�EAdTM�޺%�����k#f!����4�*w�����'��&kD�9�#�حTP�F����R݂�}�!��3'܈B��Q-1ec�C8j)����O-�n�-ao*O�7����7Cl����+�������'�a80�1N��g�=xS��ٷ�,�{�n �w0�Hu��KM0�Xh�$1-����n��?!��H�X�!`��36ulz�Az��x��V?v=W:�JMև���c]���3.��)ϭKe�Lm�U�L�áG1���w 뚵��w��8<���p�n�������'��o�|w���g ��ۜ����-���PqH�s��JO��=����&w"�#���4ڞV�����@u����ѷ��κd�t#դ���!$<�4�Z�Ǽpcրݾ���O��� �d��/a _��;�7��C(3 ��}A�-��O�,@���p<ɝB�A�N���Qi(��^��`��gՅ9�_��%��HNd�0�lf���Lv
0���`NG}w�؃ �V��={��j�J���,Pz]|"�/Y&�dF�c���w�Dy��S@�|?O��@�J�$m��P&i�ݘ�ѵ�\U@ML���F���g�6��o���Z������Rr�9�}�WsG BK�l���1}c�ʕ����$|p��P�F�$������y,(Q&�z�Y��YGzb��2X�����>b ��y��>�5P��W��K��I�%�ge�=������F�T]��'B27�%�s���5}"c0lIS"W������1�^�Sv�<���
68�6���Պb4�|����m@�A���4_^:}�D�x�o���d��`����}�'��FZ��qN`�qb����pR��݂�:���@蔤|M���4��幤�h�Rn�oGt������b	_��;�ݜ݋~q�ABbs��"�3u��]�lG�;@�QΉ�;!�U�����N��&���{҇�W�?C?��P9���#��@6�yrH�uH�Ξ��\+�jt�4�=���)��=o]��k�/��������eC�����Z��n�V��O�"Hf~��>c.�ҽVq�L� ;�L6�^�+��c��o�1�!�ݱHp�Ғ*�k ��f(�%�*��v16�N���v@ k	U���:�m�@R���������G��v'�n�����>K�Z��a��VsP��C���h.j��F?be%]��"�������ݱ�*&��R_A!節=���S	U5��j���wSo���/��[R��i��
s�H,ˉ��5_���16�W�lO�������:WS�o�q�-Ԡ�|�1���8�x�e���l�P�!b�QW2Ðp�h��J�����1%����~��T�/��'<!*)4\��W�p�	5�[:�᪢u�]����
�a
H@�|g�V$�'r�sn$����p;[9�f�o�j��_�j02b���k8��~�φa�O���*J.�
����03`��0J�m��d�O\�ԣj*�t�:$ѱo���q��_�Mϵ!��0��O>Q[��9mu�°��JxK���2G������@
g�����J'��v��W�_�i�G��T�zP�J��:<f�T����>�4�)o�P�-;��j���5�A���A~z'.�=;�����x�#!a(v����҆��;�d�ܝ�Q��tI$�2@-���D�`���R����i�t���F�}�n���4v��6R=\ʄ�g>�R��ũ���p��n/e�S���z�q�"�4K1ª��J& $ԏ+s-/2 ��rЌN��"㌆p�┚�D�h�F�����d�������L��5��k7���e��腑�{�E	pR���5�=�̿d�s �D� � �`]ҿ�55{˰I����N!�E���V�1��*�Fa'��@����?�9�e�Kn��I��,j�M�k@,��Y}mc�)L���
d|2T���:�>`1�ч����Â}���ד���#������[����8T�\�3����u�K!�r��k�ӷ�`�9M�s�(�Jc�����Ee�l��{��)<�d�4$����T8I5�κ$��1�[ƃ��Ȳjq����<�������_�{� LPޮڿ�gƐ|�����q��~�BB:���	d�
����͂��}����$����h�����q?3�ꞵ;�θ��@��m�*|�Ǧ&«rh�Mr���:Yt�j���ot����ҬV���.5�M@�0FC(]l$��d�r�;8%�NXJ⦚2�)���ql��[ade�c�K��Q;�#�S��\~��Rus��N�h���@���`Bpwg��Ǜk�X)�t��j>���?S_�7�B���%!qu��o��?�վ���ZVG��>�%��W<zv@���s,��5ۣ���S�i��}<�%� b�
,N=/�oo��,G6wI��Sꄪ����6�7
Mu@ݕ���
 ���X��{?%rQh��Bz�h�:Cdp-��t����&��,wr���R�U�J��WKP������^C)�%�N�I$�a VP�En�C�ý�b͹�Ίqû�Z�lf\֎3�~�VР��Ќ��W��/�,O���Ѝ�����ƥ�5�TdRg\��ij����<�jz�+Y�2����L�I�y�ڴJ�:�aV��K.����P2!S�S�	�Äc���x��$���t ��f�~bˇ�W��pV�X Y7��g7� ����^���c1�K���1{C�Kd�G�7}�<��y�m����?B|4a~���Į�$�;� �����	�8j[_'|p&�Թ��9!g�l2�A�~��.�d�Q�\F7��j��xy�-yH���)uS/��R[z��yC4?�u�,�4#k��aM�o�B�!��C�	%�_�<O$��:�V�!q/��R7]6S	�K����AՎ���KKO6c7�$���Ě�嶡�[	���a����d ��Y���'�4ܭ
�W�W���^���s1����%5,�9�q�zJ�8��(p��p��C*e�>��'^C�u�(t���5c�*�drd�-\��>��M�����&�5/���g易�8JL�x��	�G�܌���S@�F�9�V�CxD�JMOճ��1�^�A�Pp<a�����v���"���{ؠ�����	)S`/�;z�w�s��i��(x�P�/�"#T�A�[��Hpޮʆk�qҬ$m��p�H
��L�[�d���E�4��2Ѥ�bj>�(f#&�#_��uW[����4*�!�sB{G\��4��r����+��[�9�/(�b�k�kfg/��?��\u����y�J���j��Ĝoۛ
�F�c(:��G� ��[��"��I��i�7��n`p*�����H�V�^M�����N��%7ր��_�%
m?7��i�m3�A�kY���w�6uՔ2a���.��7�Gn��3��ż����w5�������aj&҈�H3Y	ԀdpXI2�/>Id6s��o*��j̗������s���LLz/��;`�}�(�]��u�h=q�]WYg�ȲY{*�������ET�|�����.�J;�2�_s�g�	Z.�@����p�K�T�VI��P����?	��V�[슶lA�r��Y�唰P��kL���ꁚ���̿�ˁ�t��-f``��CC�ś�Ktnfj�l[1�x\r����i���O�|��T��2A��&��r�0F��$���$p
����S1qC��&G�d�i�����^|A�<���A�Wo�ް�K2�.>�!~������=�	����Iˑo�����c��V����K�&keg���H�]T��i3}jy� ���5��Hf�ˋ?�z\'�<u(�;���R�K�������+>�]*����Y����i:_%�Q��"�ϻ�t����"���Ꚁ��u�����*�0����SyJu#�q�����}�u`cU�HIo3ʹ���ld�#/�N�f�&���O~5�o�#89h�p�����D \H�A ��~>fb��ǄzW���I�������v�k�f��q���JvY%�qK[��0��Ά���``[sw��<�ӷ	�����$����k�ۯ��]j|��42$X`�>�}�4�t=Nݗ|�j��EMy���4�q�I�� LXW��&�|�S�z^o����y<Z�6��/T�za[4�)���ݴ�H�y���Ge��ʤ�B��1~�To&=�W?R��Et�{"�ʇ��EJ��"?f*�(��z� :vO�y�8����	=�~���<{Z�Y��U�c1���d��X9�C��zR�Pw̚"x�ygۗ�D�&A&m�����.������4�m`���.���_|� �q�[�6Q��/3��V���q���@��Q�Sr
��=,7=;]���h���:�*�rI�κ��a�ѡ +ھ��%8��m���� ����S�4��A*�^U�&b�
�$�7�賁nw�$��Ȼe޴�5��{���[3MK��Lώm�~��v0�{[X8�}��D�䚥�٣�I�߽4��NR�ϟM8-,�4-�(&����n�;r����ߒ�o��3Y�M
�H�5�+f�5@$�:.U04 �2 t�'�81��<��k�G.{�Ѝ{�"Z����Nk��y�դ�xx/5� ������p]8x]�4��{+;%��uP{�ek�ν3����sE���`|ͤ��KC�Sa��)u��Q���N��4�)�����X�E�� �4*�J�
��͈�'of�\q�O9y[�D�E����۳�nr�s]c��lבV"���e�����Q�lF���ۡ�˿<�2J�l�r˫x��/Q��%�ծ�1���,���V����<=nقs���������.��Gt
�\{g̙at�w@w��� ����3�gO���.վ��3�I=D�����4�x�=��Qt6��Q	*R
�Y1��w���j�)z���¾�4�V@�*�7�/�zL���*C�s�1*���,�CE��c�����%6Z@�L��I�ޔ��t��β1=�	�ûPUu�^\1�f���i2i.Ş���"wN���{���0"V������_!�團@���~�4)����`�4>h��7̎���k�6+v���z�CC��>�����ϑ�Ja���c���(�0k]K���eDC�D�b!�DJ���e�&[=ŗ�.&�@�nj�˱�֮��څ).�GD�&Y�hU�L����3Y{kaFN�<��K� )&�B���p��0���#GY6���,�����=�j�^���h#�� ~~A@��F�rk�����7c�/�*�1ǿ.է�� oߞz��/����sȭbt�o���!�����'�Xy��);A���4���Q$Z�.u�p���<��ǓlÞ����A����eg��I�Lя3Xi@0��[R��D�q��M*�o,����^����'Hq��9c��9��A����`<���ggф�ǃ��+�R���s:�O�U-Ea�/A��w�г�d⏯w�ݦRLM�<KܭF�h��G�F�Uij`�\�^�Kg޼��( ��_x�ɭ�U�r ���͠�@3�����t�)a)jXN�'NgR�����"�&�A��!.�a]��=v�g5k<�c5�"��K3�=�Z�#�Cjfʧ��|v6)�u?:\r�}A�T�M�Ѱ^�3�̻9������zu�.w���YEe3.��P3/�{�>y��Ж�t{�UJ �Y��E+��ʭ=��/����]S�3֮����2=YH�f��II*��+�a�=�4�����}d;�\�ܠ���1V�7�E]=�wE��;�0|\���@_m�C7㕅���y/���\t�W7>��L����4U��-%�G�˞���<5@ߒO }C��*�0'��[��5�0D�Mҿ���v�4�O��"o	I֋6�eݨ| _;]B5a
�{ن7kg�����RlH�7��3��O��f�]M6������}�>	���.s�����_=th������!�?Za���Z%'���+��!R H���� �_�� ޶�c5�`�Iܒ��-4�w0k�0!�~���C�@��H����%}G�{Dr,#��@s˝%k!a����%�O��k����q��	��.%�;Aܔs�����<ÿ�6Y`�
�r2��[Lv�	7��۪:���u9E���ڣ�ޠJ~��t��Y2�l�G��+�V돘�;���mp�R�����[R���薕�xgd ���n
����rLXҜe��G�����9��To�p�j��4b4�z�D�����s�w�9��da��<�RO��GԘ,w�_�"�>kR�)�b����́`x�ū��\ي��Z�w��E���L����+ 4�0�(s��l�@��U2Sk���:��9�j �ڰ;T�l �>=��I˨q@y�  ���]�hC�} �n6&��pW������=�5��ᦀP$��J�a�'�p��5Ge�`ѕBk���+"F\�K ɢA@����p짩&3W�����#*?n��'��M��آ��]��=���������5Юwk���0X��������z���a�YD�:C�d+��3��Di\���^jb"���N`�˛@��r��²G��W�j�zy��Sg���{g��w�����>������PQ��+�B{3+1h�<�P�~��SBn� N�uW��
���#K��.(C�y�C��rO�����v���1A�{�0��&F�.0�~,���P�wdK�+��͢����d��*o�ȧ+n��@�e�31sr�NA���
l<,���F�w�:(z�;8J�O�����"knc�lЕ*z)��2[#���Q�c��������G�d�`���Q�G�?�8d��Ā���ny����g8x_�����Ҷ�bw&#�wZ�"�b��z#�ʹRF�&z�F�0���S��?u~�:\����&��J�5K���h�Q�¸���X�[� �k?�|1���ݶ	P�P�9�_��p��r��։�k�_���݄����+X(P��F�E��#5�v��V�Z�D���A[���J�k��=Ȇ�4��9\WD��G._A�n3�Gv�}��%���$�Ķ~�l��l�h��KQ��Ӡ{Rc95K��'�g*���B���CY�[�F��B@JE������D/�����X�~���O:#Vd��y���+o C>��am��x�"�]�K�IT�W9��g������xu��qm� d/C�m*�TWy���T1ů��?��K�6��>W�7=o�td�i��;=�wE��Ҫ0�0h������g���0lM��#������T�9:JLH����/ay�Zn�،�g^û�4�*�$����H�Nr�U��V��`4'�;�B�>��Z���0��ؙ�Lŝl�#�_���xB�\ﲏt&���r�:Ov�x�����/AG��2c&%dӋ�:Gj�����5fS�s�&��p�v����e�f=��,~�汴7���`tUvd�a�W�,�cր��8Z�8�P�����+�S��-r��9�-eoO��0k��|Ĺ��x��d�?�7�G��c�-�:}�R
��j�p�L���_W�.ɔ�o�n���01���:��!�!	��o(�S��/�,䬼Ao��DZ�oB>ѷ�?�p}����y$>M	�^�(��UV�CKL���7*M۞�с���iΈb� � �+��&�V+�WZÅSO�suyT{9� 1��@UK�J�W�{^|wr��2��,;�2�`��4BW�rb� �9��$���!���=2����7����>�����߹���-���w¢`�/s|�=eT�60�,h�Vb���t�˒�>f��0�C[�����ݣ67,]|�'�����M��&��b�h���[�
�_Hf ��+u�8�	ǘa���楏��m������s:���8�{E}�T�+5�?yE3�f��{���=�I-tX]o�j�ĿNֻa��9�$i�r�m�F�鶴��J�L2I�� �u�U)Q��L�i�P��i��1�4D�B���� �ByV�z��_d
Uxϒ���{���1��+�q)μT���m�WM�|�5_0MD�/��+ɣX�-D��W�P����]7���0V`o���dTc��~�v1B�f+�]�q4~�j!!e�VZ;I�t6 �U��ؗ_��ݙ�䒀k^U?�0?���Ȭ�ǳw�lek?�&0�1 ��O$%`j�M�s;o8Ѝ39|��h�ӑ�@	�s8��w�DKu 4׽�iH�t�h�I�3���7d�mf@Α\����7vO �����d�
�p���`����R�����������S��'C!��E�,��<������a,�sf����=�å�����#�sM��g�9I�Ed�M����麜�`~�\�֋���"��=]�Ջ7#ˍ��#�����h8�a���E"o����x4���� J�2��x��(�K��%���&S�4}� 0�5m^Or��mw���W����~�Cj���ANF�耬W��z��33� �T�(5��孅�\��n���Jȇw���K���.ǜ� �5ޖ��J#*{k���c�
�Q��/9�<y�!��(Q.�^H�R���U��T+5n�!i�8�#����f���R��~%��߇+�Wn9T�l��XA~VGn!`c;�ᆇ�CO�$�]�7�DIC@� ����� <�,����1@��vw�jR�V�rF��n�==��CV�E�@��X�x�ߜ�:�3���5�l	����~�{��\�;�E��X'����BLA#���F%����"�v�v���{�ly�*,��E�n��@g N(���y���?�A����7�G�#uD�K�2Q����֢ǳ�~�*�����`�yK���1K`����bF��w@�����)p���~�`�5�F��֔����!Ĺ=�ȥZ������h�؛�P 1�$��xf�\)�6��t�x���$��&B������dD�C�[������|����9��c+{9�1���s�s�a������e�awq]\��8ҀԕT�D�Zh���cO����;*�łt_�EQ�;������F|��J�]�K1*�VU��_ޏ�5�M�IbV`~&7��e�n7a5��]��.���q�;s'v�$�(�-�X��%�yV�w���ޕ�8j�n�k�,M�\��c��1���t_��2��)ւ����Hk����TNL�@�!k�,�&5����$d7N��ښ%dj�iu�3�Ldh�i�����]��u�nA���^�!�e/��j�_�'�
+qŌy	ݖ��b�X�0�M�g�Y��9;�.afy����ךc�PjV*Z�A��Qi?�x��"�������]3�"��=/���cU� �[�y��������0�^>�RX����#q1�bNJ��l�E������dܲ�sۇ4�JM҃_S��:�]!���8��G���M�=�뱥�a�!�N�d�8���fIq:`�Pa��sT\�_�D��J�QZ�,
.�	���[��K�-U�2�6춺{��9����_ ��c�h�q��Qi�[eð�)f�!,��T�6N(	e�1]�劏vwO|�z`�ځp�#I'W�?��,-�oF����2s�=~�	��+� ��,�����o
�<U��iGV~�����e�y��l��HQv�8.�\���T�s-��Rmb��i2�5,�!p,ZE0��~漓ʍ�X켉f��E������jwg���MCL�!�/�U�D�O�:�E�[l�y�v
]A�e�_��V{��^���ɟ���@�qny�>�� �4���C�������7�{dYi�M ��j/.��J��',�� 4U��K���1�%���5+��D����.���NYU�7��c����Ue]y�!����Y�B�Hq���}?+9EAa�yJߚ1�/��6�b��5��p /n�\�6v��)(<'�e�bC�~��/�ٞޥ� v�����y�t�97e&pr��
�y7'p�{?i�^zAN�%l��Aq��k9+����%+���җ�	�w��n龺�WC���+�sX�[\�H�Eԏ@cWDA~��⪘�exg��L�#]	��/B��I.��
 ���^�.�Kɉ��(=��������.p�d `)/Y�/� 	a�*	������};�F�Z���I"�>�7�s�:�]�f�qc�O�Et�vo�M�O�Л�3��ڗ��i�O��l�z�}�� �ߙ���=yaw�~Т�@�L⥒��&;R�d^�!DQa�)%�B�ңybX	M�~3E7���V.-Lܚt�������yp���^�LGXH��+�X�f5�ŭ`����"D-7;�y��|3�@더)5ٛ������}{A?<]N�6�����q	!�z��p{5O�����'Sֺ4�m���M^��/ܮU��,�<C�Gp�xI!��^�ڒ*�1��NΈ���y�t��F-��#�bN���ʿ��C���'*��h���9|~���4s;��輞V$}�OI�+cp[���k��+S;�C��޶�p Q\�s����^��p�b���2�K�X��If#��u�Z����7F��%�R���y�f�����:���2;��k&pS��.,�[$�s�_�-"E�w�:L�o.��3�(��J����o�r#	�9P�� �{k��v��0ho�;W��k�^�����سf�y/^��Yr�ɩ״���+͖�Rg���!�]|�X��rV���>捹EU	����q�0��ٜw�?��D��&eet�iF=(��"xB���ꅊ���;F�k�S����z��^{�2�Mx�z��LGk�x^ǚy�gk䒲�T1{=�w������'��F%�6���)~��{م/!�>���ʚP)d�Xߑ���u��3�)a{B�u3/"�j�0��hE��ZvsV<���3�,���:����� 3���i��A*+����6��˿d޸{�K�L'y;M}�ӓ�FDbB��G$c{-)`�J�n����~G����ữ�v��?�e�����Q�"}�:С��	X�*�Ѩ�'�$C�pyU�g\�j��A%�c}%[��j��Z:p��)�5��ӹd>��<"!�!�j�����:�k�x畿9vW�Hr�mÄڷW�@4�T��{!u/'������@�v�Ͼ�� ���lr��=��_�^u/�|GK��{�G�O�&�lO^u<�P���c�h* �����#8�p}�?��΋�Gn[ipt���6�ܭ��e>w�"��N����Z��XU��ټ{�4vȜ��m%��9q��C\ʉ�5K�$�6�4}�f)0�s:��S�(���Q0��E�b7O��15��ɣ����nPh����z?���ⷝF��q��}�E�����My�X�ҏ�������:@��ܥ�\���u�I���v��/8HD��?Մ{�I9�����^Z%����U+%��δ4KB��O�q��B�~�V�Ht��훴��7���@R��R��2Qj��t��k����|�(�����P��\����1>�-���5�2���Oo�QǍ�Bd	�2��h�r4�I����z5(:^���HPv�����J�RB�v.7����<��̃H|BF�K�`XȁO��[갅RW?����JK�@U\-a�>��v?F-ek7b�iY&��W�Y��cQc�*�?��{����!����r�Z��~��x�y����[������9s��쉧��c��=r�hk�
8|�1ng+Ø��!v! )u��5Z�I��z�t� lFf=�U��C�������1��#�!�񖙷�B�A�6�}Ly%2P�r]'�6Jz���-�!A%K�!�� �w�/S|4�|��mg���B�TQ%@���)�H��`  @�2���!u��-25���y���[z!dZ3(~:WT����^�e���JJ~֏�B��6J�� su�+�].D�X�\��I�D�FI���r�r�`�(Рp��`�
l���ْ;��<��g<��[���]�EzDV�U1�	��<	ُ3���eڻ�p=��	 9V�b@���q]�/�M��vg$']����L�
H{Y<x!K������~
�"�8㸫�d�l��O�2	��}�s��h�$hˎ��:��a@ꄉ,>��~��F!�#d�s+�#K�����J҈>�[|���rY��
)A�j5��\�aU�Z,A-�`����LǨ7��r��aOEJ<F���;G���0��d�N��p�+
YX�4l?�}�N_D�������Ӡ��L�#��)d�t�o�����xOI�;�=TC/��%dh��odp�gƵb����כ�2a�������'��� ���X����3�T�"nOk�W4�rݘ��G1=�T������Yϖ��*<۸g�x���%tF�w��q��u	�}?��k�@��d��r�֨����$���$�v���{���+��^����*NI|���Z>-V�u�Q���G
cS����Rţ{I��H��L4�����q<��y��W��Ю�d�|�_$.�;;Z�N��z�]6-w|C���`�0ϖ<��00/w:��dУ����+O�����v��[К�ut�]�gn�[Fm�;(��T��̗.A*i�)���}���\
��#�+`��0	qc@Q5\�A@$@�B��F��������m攭���ڷ�����Y�$�^�/(&�X�P)q��c����<�� m@���YGx}�#�G���A��4G�8��.-�l��f	닄1 �����z$��z}��iW?�cZ�̛eb���H�ۓ�sN��R-�l�c{�/w�D:]�*���1��������=-W�_�+hQGԗP�|�sØK�^yҬ#����#=|\~/�G�����3PMm�"�0����8@�7�$����Ĺ{lpW��m,.)�'/|%��r�{R5��)��%�O�M΋��	K~���1���)�S�J�(�'����|J�
�w���o�lB_t�ǥY�K;5�{l�X���i��S��/c��M�no7h�y�7ܳ&P�0�R����)���"�&��[�ゴ W�=�9NT�I�-��#5?�>gO�6n��M7ϼ� ���Fu�����x��n�F�D�$�u�:�Nm�qG��А>�l� X��qL8�\��2��s$9�n�ы@&o��M[��%��zuܣ|��r<�G��ݪ���Ȣ��Y�Ǧ�JO�:��y ��K#���v'L�R	��� �j�(
e�R��ü��6���+B�@탕͹�.��g�Snl+��&��?��sm�;��0��M~v��ޮ�6������莠T.ǋ���{�ӡP{�*H�:����4�q Ӆ��ů`6��M/9`�|�W�]�2���,y���$2����g���o��4)���Yh!x3�R��%4-q�/@�T�nF�졮f�d��J�*�n�������C����4,!��t�k�">�#`qt�'�B��=�~�hCˈ��K�X��M�[11��������A�{N�7*����~����Ӣ��K�y�ȩz�W�!e����o��Kۼ��4Ǿ��w;�"�2��ן���^5���������V�)
��Ё���+!@>e�P�ſ7S����*��oOZ�� �ظ�^����C�>a� ��%
J�4o��h�\��tr;�/��q�%x������u���mbǠ�-W����;ou�	�싊�׉�D5��J�d�*��٠�f���YA��r�OP�_r^����a�rL��>���z���&B��
��|~&��.^�׵ �)Wז�+�������������-�Y�3��/��R3�߁4J3H!���)�`&o��y���Q@�3�d��c ���\!b�QMf~9��ʑ0ɡ���mz#�Z�!w�ݥ�9�Z�B/(<�Y3[X�t�/{b��a���:$��~��8BhK�z��NN��T8q�uZ&yUj�Z�|��XӺ���bó���� ,���b�_�,ag���_e�8U8�0���F�^�B�8{yM�k�&���^FLM�,7��q9J��� !������mi�J��cN#��H���%o r�J]C3�t�sxNԔM	��U:O�謶h+놿?[ᒝXm��m���:��&�Ö��<p̼���\�<���&�'Fn���bN]����<r��$���ѝ鸎T�/�Y"�o�?��������`�&��߿}��P&� c͞�[ڨ��uy���{"!��~]��Z ���Ak�o���L�x{�w��71�ےֆ#È5*J��_�8b�XϹ�.�!����Ѓ5��۵��pl���i�x3w��S�m�G�1s�}�?��!�r7��:�nC�pmeT8^�o���l���وvm�� �ɀ9�6s{y�؜��!I룞[�i����x��tW�|�@��v8+�����c���`�^����YEл�P9�jb9}��$��q�%}���<y^��m�<d�������<��;u�S�sv�e\�
��R��%6Zˠ�@�u!}	ꇴ�J���7O[�{jԡ�k,T[6����/�K�$_7}�8�nϣ�ǆ ��*}H�?(' f�t1ڒ{ �;f�MU�p�b*���\�}������ru <"���5�!Ij��fҺWT�b��*�p�	�A�{��L!�" ��G�U��%����I#
�U����{������~�e4q�c~@��2%�e�
�F��09?Be��aw�8+K_�d��`gI3jUS����YY�v�*�Ȓ`c4�m~D�P�lA>P�Cj�����BpU�E7c�B��;���/*�:�$֗]���f�������9kޅ�/�X"�����>����}W�@u�L��w�����$�*H�I�p{�Vx{�y��<V'x�0/*�;����D�{f�O�K��}�Qc�����6��׻H�)k�@0�D1�I�M�p���W��NZ�`��÷����2E�jH�h����u�c���R���Q�J���r%�P[B|�?<�ÔU¶�����ǁ���w��%���Uy�n/�:����X�Q��=�v!��1��������ڠq�맓�8z���-ۥ�<��-ҕ���j��c�����E�ͬHy0X`���|v��7�~�a�߃T~K�׾n�.��i0E�T�����dc���@����"�t{<C������5z��e㗀�g����Vu�4�2yt�����Pg�G��� K,�is�+o��7�3}_R��w�M�R�I�$���}hw��xZǝN���(���+����+�7�C���qӁ���|�ǌ�A�yl���Ϊw�'8���2����B�9���]�y�W��O��� -��4&���[� �7SR��S���U���ڪ����6`E,m�A��[�ၰDz������@�/v���ܶ���"SJ�1��G���`&�^�;6�L�ZB�4�@���&��bx��k�t��Q������Ń邜f��"�Js~�|�KV+�ik5R;d�a�s*�g�/�I.0�p��4���>�I��:���.��.��N2Z->���S��n�ݫJH�_uq�*�%�U"��$��)q�jD��)�g�p;���k]R���
S��t9Mg�]��K&�AAn�"���OϺ]����`���a<A�* �������dhf5�!�B��N��YPN�3ǈA��PO�M��J4@<�򛎏N�{`�����7U@�?ŏ���H�|���+����k2���,}C>=�������W��$�����{V/���B%���r���5�A#�t<E�z�fR�rk&�bꂛ�8{j��S��	~�u���P�r�
��a;��boS���U�k%hۆt-��7���N���x�)�#s�(�[\�r�+�F��iAƽs��T��!�O	��W�[G(��K[�Q�V�i�8]�_(��')��!�XA��g�gny�!���ٮ��gӛ�W�-"B�`��NA���'S��6��$:�'*u Go��`y��1ol�c6��E�$v5n�W#��*�����\�`�P_��`�<�S�2�B��tM�L�&f��%�XIL�Yh_�-+}���|xc�Z����_�YQ�엶ٟ��\��X{��zS���d��vh����q��O���36��ç-`�����g�2�E�֡uW ֆ�(o�xČRr`��)L�pp0�\*]��Γ�����<+�"�$�v8Qb��c���C���+o;p���
�Ix�\P��=�x)`��1xE�M݆<DJW���2$�Z�v"&�x_)|�
c��{\�2���J���#�fJ�ɨ�W�R���.M�)� l$���L��ED�jm���>P漠��c�69LjtA ,���oO�R���^l��V�.��Sn�	I�Y����L|��]��dȗ�%�#� Tr�l$�*싙�M�1�oIu��K��=t���z.�z������~�4��]h�!ǳ�mYCV@'*�������..�A��z1��)�Q�S=�96٦7r�J̑��!Z��58��lq�t��K�g���m��Gr	F�R6��v�&I��oK�xOO`�_����݅���p���d\z6ܧ�0�/��kt�ɹ	"��2G�p8��ȃ�ݏ6EJ^��B^�Y�ԋ���3t��k����ܯ���E>�$�h�^GX�ѻ0�@1�`����T^0����ꟚlK��)�2��i^|K����=z�-O[�퉣�ݙ��X)s��n��~���PN�+y�Y�c�r��=�v��Jb��~M'}�qd1���D�W{ɚ,�e�6�Z��X�3A�x�B�P���6�x�^{����oq�_l^�w������y�;�7�,B�7�.�s���R���Z���?4h�/�Ԉпg�>q����4��ʎ���������(0ޥHO��<b*�nI�C��IAw���$��l�q�/����,B��f�A����~�|}��/NS9�~#Ќl�R���x�����*j}``�xfx��^�׷�e��I�	�&J�&�!z�C���4l��Ә�\�c��c���F��G���؍MyEZM����\"�e��ָw�И`�}�^���1L���sը�6_��_�t��)2GfDȊ�(����+��?�y�G����iX˜��-i�٭��]өh|˨����`�1t�-�-2I<�3���qK�}�ǽ���r�h�e}�٠x�.7Ǻ��P�	7/����履s���v4F���@�#�G��j)�[;wױ"��5ZՉ��n��K<�61H�gV���ړL;<td��(`l�m��ν�o#�n1����%�xF;?e�0;����N��X!Ԙ�h9��wYd"�t�V�L"�g�n0T�xT��lg�9-ڟ�PbO�!��8	w��t�� �+�.ng��9N�,�i�m�64���Q����9���/�C�.YL�L���%���K��"�
87ź$�0�s�I5��+4v��~���:"�e��|@�8����~�M�����A��/؈���ھ���a�^�j/���Ō� oU�� n�i٥��D�XG��G�.�>�?��b���[����l@�0
&�(�-���`����fxp
WwLӒ�Ig�s>�b�bAl�!�i����:^H�G���3���̣oX8���y�;��C,J:y�cH�t�T��@�%��S�;�5�U��`���I��K�����C��SR{�̾��������$���<I�����G���^ỏ���	��������WJ�&ȚڃzHf1�1bo{:V&��V�A�Q^��=��O�{��a�d��?�~z���v�����o���S(��N�C��y�h"��Ņ���u^�����DpS��E��6�g'���W����ʶ/�s�!LP�5Aeg����h��>��u"u����'���`+�Yw�ʃI�����B''T�ס���j�sf��'v6D��3Y�BV���z�!h��(u���vCyZ�C	� �#��.�����D���^���9,�!h*~�[�)�x�H�a�����	��T�� 2kEZH����q9E
�k_���I�S�_��A�ɦ��F������g1p�w��?��ke�����[�%�i����a��	�K ��F 
ϼ3�����AKƙ7�4Z��|��WQbr��	�	p�Ob�BFl������m&[hc�փ>^���+���K��yd-9��HB��6H���K1��}/��T�=����W�&N����O���َ6���nE�ƙF�]Ki�@f�֖�����*\�V6	�V����8t��u���Z�܇`o�	/�-X\ö�y�Dd����h�ˆ�%���Ex��a�OD��Άf+����r�� ��9���`�	����ݒ+z�+0���a� H��_ߎ�T�,�h ]��i=�>��դ8MKb{�T�S�l`0�W$�\��U|�>��̭��]�`��;���{)����пa�c�S<N�zϬ��a��T����	y�D�ZfV,�����
��|��`q�`�9��m�f:�i
7�^�+�#o�b�@��MZl�ҝ��a��^x��ʶ觌��Yj�ՙZ%|�[ݸ��=��Ѕd���>��Xc0���GD�96�1�a�v�"�#�ZY_Ӌ�]�y�E����:��#T")�~)&��FMB��(rེ̲|�������q�����M��=�N�2TL����:%���^S�~ѕL�zP��XY �l<��=N{{-ϼn��G�~�c�߾;�́�S|�&�d���0�b���X/��脜l�!� ��l_�EMrn*c���'�gj��qCe|?!��Y�<푘�'��ث5opj�M��	jk��#��p��n΍qn��݇/��w2 }|SxOa[A�j�$�J�}�_+p���[���(1P��% s��/^ �]O)uB��V�W��h:d��$���i������G���g�Z
�x�$\Lͯ����{=#�nE�
@P���I���+ �=�[>78[jԒ�_�ӷ{N��B��2�����{+�)/|W���:8�iVB6� �̓��]���X�1���b2
j�p)��v3��l*�
��������J��p���l�!M��7#�ii��������f�����O�W����ʍ�d��0k�ّ�@G��3 S�|���?O���"#g�����*����_���J��U����@���9�T�� �U��F�"�NV�9��^�ؾM�CނEk��n���2ّ%P�a:d`�׎��&��P줢�g����	9Gߴ�N/���ρM4d\TKHj�6i�sa>���8��(de��E"˗�PZ#����g(-��2u���#?�lSc�9i�HA`&���낚�lt��������+��K�Fa_Y��M���W�u9~���f�SP�tR}Pt~\�l�K|�L��Ou�����_��_I����3Z0��Ŷ��$^,��u�Wf9N��T�䞫����߂w��t!@�π�NEi'{���N����ع��6_V��uR��U���bk]!��6u�>2k!�'�;�������uw��R��a�x/Q�ꕈO��[�?�K֚�ط�1ɓx:%1W�����E�����/�=?p�D_���֑�۰B���:�6�N�b9�.z���F6��n��98I7�ת�`��O�h�	q�Xl%�us%)oڬ�g�����͌9�����t%?�'�)�n�:��2׮�R�l�����c��u�}B��]/�$������(����R�t�N�7�x�;PY��Py�PR�g��nz�]%ŝG:R���8�|��B������=�z����N�1hɢ�W�2g���٨ڛe��;�^w�nV��6�0f,�nM�J�4.�Ȫ�6C�^^y�Q�A~`��K�mO�dsT��E�b�^�~~^��&���o���j�_�`Gu����SM�uf=�Xt�X`R]5���Z��/�a�{e�-�<�Қ�p3N�
��E���r�H�f�L|�a�d�MM�
�c�ۡ>���������3 ����K&���c�dǶ�������~�UeR�� ѣ}���8=}�����_��1����Ҥ!��
��a���g�!��뢮T,tGO��K��ƚ|2`Nk)��ʀ�&��c$7�\ܟ3�2��Y���uG�q�h|X3wh��"n|f��!#	�)v�;[�NRK��i�x2��b�������=����5�.�*���mh\��>���d�xTj��� �C�h���W ���	���q�?���&٤�I���h\lBHD�M����&�yf��h�YLw�u�P�D�Nn����Bs����!���ERH�eQ�֒� A�qr�1!�\��Ԟ��\�W]�,��6��������va���Yh���-7=�{?�O��tN+NO���������.=��6����{)���	���x� 1.�n>���	�s����&���d�ys!��I��6��Az?{V�,�A�"ȥ(H� �]KC3��x#}�tA�����G��=+w���g &�`'=�I�q��|�ʿa,�&��R��&����G�ф ��٣4�"��B�Te�����[�악-�#K��R���12��i�N�J?e�r�N�!:J�L�z�-��.g����e�CCN̎rX.d��J	�͙yVEY^+�db�9�e7����]�һ���v����?�r�yɪ==�T�L�����Q�tl�r-<{��]Pc��	����uMj\Kg��r���}5y=G�l3�~3�V�DČׅZt��$���ȅ�s��"j'=���儲I����E��:��:����$o�_���^�G@o}���}9�^��+�����bh��o����5]��-�qe�L{
���/�=u^Q{���'�Q�ť��Y�`;+�!p��)�	4��Y	Bj�n(Fi���B�d�c;�YÛ���U"���y���XS��%5	��1�!���^i�]���Wκ�rd�9���_��?���_I;J0�ץN!=���	:����K�ę�� i\l��bDm8C��@*��E"�=L#7�wKB]38�X;��#&و�S����N�~#n4c�	3�JR�ƨ4�B���7F��PKU����/���U���4}��|���t�V�!;?;�f�a����d�"%�P���(���q�pE�l�Aǋy��D~֯���C#ڜ��_�
��2J�mLcQ-<z��L?��ch#,n���W._�)�#�N�Gw�����~_����!O�$���CD�;�oe.^}�H뎿��;� 	1>�?���%��F���,r���'qUp}�IO��;k�
�:Be������d���ӆ'�'P��^(�	�z=N�@�o+�� �^��c��H��o2��zq����x�̈KwO|m0w���F�L�?�����٩J:���~:=J�OQ�|�#���.uq�_�9L:Ĵ
"�E����{2n�x
�4)� 6)Uq��O��Cr$C�X��Z�1������1qkbb���u7�d��x���>��5�R�]�:1��/xOխ�q�C{�wH���G�۾d+��ۢi��S�F���5�i���f��`�eK�Q1�=�ј"����^�Qz�����Xo�P������p_,	��c�G�_�?�&V/�}�eفj�_1����������N�Zf������ƻś��]��n��~
8ũtw�P�S�;w'r�t�6���7�fh��M��-+E�[�~�̝ޓ>Yv���q��I]'F�>m7A�E��xâB�97r�(l ���L��*a	s�5������j�3V<M�`X���ck�ui��+����w�HЃ�>.�e^|���n��|6XC~���EI�*�������'
�q��m;���xZ�C�IJȢ�!l|��i��HF	��u�?���w�������5y�$���6��v݁�]c�S�`�ܱ�Ğ"L?ˈ�R��1/�~M$���m�#����O=pԏa�
%����0���%���	��+�����݅jϹȒ����@�^ޗ|k�S��ujBLe|8f.��/k��4Ͽ��Ϡ1�����x�� �|h& A�>��<���V��ݹ���[;�o�v&�]��]�3$C(=��YG��H�+���;Cڤ�_�m��#��}���l�ֵ��f���Tm�Ñ���~���15���ѹ�rs5-T����f��sS�g��݌��9� ���k��}Τg`w��\ի�l�*,�}M�i���x�b��c
��;�a�ߌ�8W�n{���d</��ˁt��.~��ab�A�e���Ґ�z��UfӇc�aŀE��+��{)(ڰ+(�\��&��۪�hVn^&E��D�����6��ݲ }5���.�|�#����_g� h����T��7`� y�xȕ��������������S�^�Ѫ(�=-���HX��]+_������Ղ˙0��;;D��@��ÅS�Y]R��H-���B�Q��B��)?����&mI�z�|LҠ��%uR���mA�HBj��^A9j°�؋@�Y�D}n�!����應(�K�rc=��(�7D����(��X��B��R��jY�⸳���u�!�X|vP�CHS��ِۢ�3�j�)�Б��o�q?�$eg��Re}��UL�� m� �c&���sP��hJ�V���[V�z��g�]�y\}Rr��ޱ^ھ����%|�2�[�(?"�{vX�{��GΨ�ҺMH�K�{���4���c̒���S��@�C�w��؊�1e/$����ѱ0�^,��!i2�>���/��El�Km�ωa�L�N����·�xX�~Zd���&�d��.�L�L˭*������%G/$�E籱%��E�G����p�.S� �+7�5d�+9�/��̂�q�]d�X͝�ud�>���ݲ�bQ��F���%dL�a���
�Z�),Zo���ݲ�����'�-���6arŵAH+96��E*�