��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�_���v��	�������d��i��HO�4�H`���ul]����_/���g���s�K�7�,>�Ezr ��~�'֗��O�( �,Ly[�Ლ�@���f��4���fH�M?G�f^q�3����&�P
��Q�=�\�1���|��ס��j�/�U�xHg]F9��E�H�z�O��$�G�pR��\�`3��_3��ߒ�#X�ŉ��e�� ��c( �#��+8KE��X�C`vθ��m
�מ�nA�s�.�����E��_bXӰ\�Olj
��Kݦ�|�a0݇o�s���J9���?#����W��}��T�7�/Ȓ�A�Ma������0Y o�S��V�a��k� A7��R�M��Ԝ��9<q��$=8��Xx���^��̙�>
��t[�s	ogs%|���+U��:crJ��=�_�`Kf�YA��/�ev����z��{�.�G����BsX#n/�X�N��	���B���^t��}����ҭ��ZN����� s���S�8R�p��{�@?���`�ؔi��(LTE�)��%�!o7a��6��.� :�7�Tvgթ[�< �����!6�b���>7�AdY!&?}�$É��z��OE,:/(�>��/;�3QtKZ`?{'�`~�Y��S��6�9i�a*!�`IY�����T"�8<�y�o	��m3�9B[��չe)�O�C��:r���8JE��S�7������W�hǀ͞���ʃx�?�s�uF4�A5�B�x�A���b��H�<�'���$nuL��f���Op%��G�����+'���Z �\�N�?s]��ۯl@�K��_�;���bQ�p)ۇ28�X^X�?��Z�U�y���[���tùm�aQ�G�*9j�� qcCп�G�=���E8պl�+̑:kC�\X�7��h�(vg*
�䡏��T��|����.���ߪ��9Ӽ`>mkpA�B\!�ȟ|�]�2���|�rZ�}Vw���M\v&��?�����	m>�&n���G>���m<SFG������]k/7��Q�vq�a������.W����N�=Ӵ�G�ؓbyc���b�v�q��We�"�;�r�7������Ir��T�������l� eb�9�K+��<��`�m��E��9y�gBUX�{��f���Yi�yMh�����޽hvQ�L+s�e�Z�DFT'��5ǆL�� �%�S�b�?v�	�E3݆@q��Ĳ�]�n^C��5��zx
T@�s[��*9��YO��
��m2�u�%WF�G|~�����Z��,wQ�T|�~��d�.�@��2�$�����OFj-���Ŏ�f����P)�ㆻ"{�^ E5�(�**d��pp%�v�0ټ�n@�%��O���9�af ����o����P�J���+�#$��4��A�v���쵗�H-�"�\9f4,��ͻ��	|&�)�L���JB��ib_�"TB����p��8��Q߰�լ��QA�c�M����W��n��<�)�>}E�{V��yd�c��v6�գ��
�US��*`ꤟ<���e��7<���N�}�m~#��D�k����U *B
^�d����)c꘯rr��g�jN�ˎfJ�x����"�&��� �I�Ô+J���$p,�:��&��Q$�N�|�g�ۂ�LHhS�ԡR"�?I�BmD��j(��Tg#�ClU�~�����A���d�~�/�O���߇�Àb����a���� /��Q�Y�.e61� ���Η,kF���ߢ	@�ӭ`X�%RՎ�J��4m�ty�&;c�b�U����,Y�.S��0&.גm�+�8z8<j}5�@����T_r�y��.(��`J��.�n/+�kh�QK��؝<S��z&������8�̠�P���g�C$n.s��c�h��H�kA �oS����	���8�7["Ym�~��l<W|\Ef�Af�^'!����>�{�5�x{*/���ũ`P�J��ea��a�+\";��󊉽�O�4yD��J��6����5pᵉ/�r�k�D������B�t���='��zw�l�Ջ���l���\�/��?��J��i�O�}�**�(kԙ�Wm�MM<{�Q��b�����)��̻e��VL2(5rZ���ŋ�����yk�:�[*�M���D��v ��Q)�W�=T��7It\
(4^�KbG_=r�h�h_y���j�Y�Ƭ[JN����y���_�rI��p��1U��K�*�rc4�ݸ���Xʖ���ũ��lХA~��B��±J�)E�j�E��X�yw�pP�<��Yhܭ4k�Ҡ�_��yu��N=ܭ|D$K����g�+���9��a��BO���[rC��O&�~��G01x����D�4%��l,�t�Vq�:��"��)�)&�]$�Hߎ9�k��?��a�͉�v�k���8\�r�4��՜h%l�H�-n�*�-���.��}!�Lw]ew�.д^��Wo`��J�/wCi����0�vHn-6u@�)a��01��
����s��ڮ%�kg����FW�HrQ;'2��h*��u��Ҙ�W�8b�<�X1zk�n�)�5��K�U�+�����uI
d3�P��+-���qN�DI�ķ�%��i]���<qE�d\��+��=�u�䒪r�C�)eP����2	]T�p�emD�8V��r�-�݊��Y�_|c����0.�M��GN�'qJ/1�nxuO�7T����`\��*�C/�ا�"�+;,�RՏק��J��e���r⟜�N��w؄2� ?5݊�$v����nM���p�?ÐVҐUA�jy��|�����'��eB�H��i���y�N�.�l]+ln�&sc�F�D�e�.߿�"�O�+�����_)�m��"���#k�y��J~8���ޛ4��%���f#��ǈӤ�$ݦ���pE�䚯x��
�!�_5�Lt*��c�Rb��~�.�Sp�|Ƭ�9�;�<D���������VW.�ڭ�*v0n�����\M�s�`��kAԖq�r�j�b�MR��<$��X5)�n����ю��Rd�M�B���/��Pn�.H̩C�[^ik��`�T�}&�y[:\��z$�C��;D��eGPJ��13Ǜ���RĐ�?��a�^Û���
�Wg�`E����q*����AP\s)��7�%?����|�C -�p�k��z�)�O$U�Ng=�E�Ck��r�y�1EV�ձb�}�q���h�]�ao�HW��f6'�@��9V�_q�����3�Yz"�֯=�|ҜdLd~9v8�$�+l �α	f8Wy����dEø��ʁ�����ШfR�k�C�[9���`c��⢧�bN)�Y&���ҏ�d�vB���̊'���ƖhE���̜nD;��}�����j<vXe�>`^����cW1w��@P�LO��a}���T�G[6GѤ�d1&J��֌W����4o�,ow������oN�cp�P��&3�����M�%?����~[�!n�.VȈ���G��wGz
\ءHz����t���#~�=��I����&����w��.%]#Z��J$�ұ�$I����R* ���ylG�;��s��w�`�LX-x*5��B)�-IޢU����m��z�h�\����p�_��ό������|�J����zИ�:1�,I��9v3T��*�q�4\ih���Ӷ0ȮI'����Ӹ�$b]��ޤ���Z. c485l�$o'��Nă����Fk��xg��T_�����t�Z�������tKir �����@N�O�����H֜U�`�!_��W��w���}Ey��&��߅�>Mհ�g����_;��$�a���i����D�_�iF<�LA�H���uq�6��TK]N�qYL���F���V�������n�j��?-��:��HCV����^F`/Bl��8�)+V�(Y:�tQ���~��q��R�}�����<!Qp5�~��#�U�@d��7�ߖeg_4a��s(j�1B�9��!/ޱ磯�����;��Ѩ.�C��h�����I����PW��5uԀR 6�NS�J�kK�ʌzS`Ib�0��݈�}�js����>�KKQl�ˤɩDw��0�o���.�Yj�S�z����Ѿϕ�e��899��SN���{�'�y�]�R�ҋ�G0���2#F#����i�0�v5aT��c}��⪴){z$a5~XL� �������<V$�n��	p�tj�^�ԅK��kE�q�1X�S�)�e�-�m]��	�,��n~jq��d䁯ڣ�ÙQjpi8��\IyD`���ک��n�=U�S�ԧG��-c5�jY�K t:�e���F��
�� /��\t�g�ҸQ�s�W�t�C��p�{�[>�͜�e�ޒ2K��o�)㔟w�W��jo�q8����ȷb�[zHѥ�
Zp!�����.		��u[����[�?���f��}�=��"Ѽ�����$7xe5�30��}���x�%jߟ�*��5E�T&ìǛ}o�����fn��� /���~�Q.l`�&����F�1)���y 0����)�a 6����Ǉ�Vq��=#4#h�<��~T����a
>�횤,k��+���4��rjvt��G'�ߪ��9�X�M�����q��?�y>�N�����좙X�_XD$��U꾘 "�NA�i��;���e�96v�%��_�L�=��^jI�Q��m�3a~@��Y�H��|H�� ZO�X5�s�����z,7������@��z%4b%љ�G[���Dؘ�I���g��#<�L�&KO�$����A)���ok�mE&�v8i�f������_"�&��s��0�!��WR�>��O���G�C`����k�*�O�dG����F��b�N���|��tE�j$,�*��1.B��[���ݝ�d� �M�[sj{�C]��N����Oy�����r���Д�����?�d���k�A����[�6�u,z#�$�k����
=Gy5![��|b�b!L%��`q�<Ć�� O��Jt����Rx���'x�C��0/<�f���!�����++�� �Q(ZH؉A��ؑ6�X�B0Kҟ$�[�{h�p��5��{w
�k����E����) B@�87� �����R  �p������������uSE��$v��VhQ}ng�����@���si�����E�
@f�|���Q����D�1s�R4����I,z���8`ixh�d�F��|~�=F����b,��z�z������W��VL�u!��-��IQ��TPG�<����"Gú���/5KC2�����-��_�����x+^A&׿Ց;�!�@�t�q�T��(e��hқ!�3�~0����flt��@rt��c6�zu��2�ٓ7��R�{�F�5���h�I���NC��'M�2.J�Y��bj��q-�=��:Dآ�Ӷ�"�Z�2��߳�q���6��O��?�9�j� *�ShhD?�
M����Zq�-	�9�s=o��6����cY����.�W�~b�͍ H3�ɫ��V�c{�J�%B"���"�ė#X
�ay�9Yp�vnW�6|l>
���*�0o����u,S�S�^4it��G{I�gɽ1���Ah���U�5�������K2T��@9�"?s�mg�Y�]k��P૏�H� omƿ�j�U��h�|�7ǎ�������?u��4�۩���;a4�.�є���`l&�5\���,�0��#x���߰�z���ɼ@��1}!n�2-1<^R�s����%�8,OOO���Z+Ϸ���H0��{~k1����!��g�*"��q I��J����7N�er�� �x�Sh
�!��h#�؇��U��p͒����䉿an*�g:
Q����j]��+M�s�vC��w[����V	t/�3u�>�r�H���.m^Ճ1@�Mg+�v�Gtg�A��2�E�;���J����>CM�Mו+`Γk*D��:?�6BI�_�t݂�{^��#ÌDL�=��!�͸��캭��ʏ]�$S�uuϹ!Ɨ	����Q@� ��?��J;8�����^���QC %	X��_P!��<�i�|�����R�3�tdԕ2\�a�h�a�ZG��3�S-�t��Bl�%8iA��Í%���^$&�-lL�K'�#&����ny~�,��aNS�g�~Z�K\�~u�=6Tz{��\�n�S�A֥�H�h�֕�+�tJ2&�۲3^���9��6I|~���c����c[�n8��}P!��?דjә;O�Gm���eA=��*��*a�^���,�z.��ޔ �bښ�@�Gl���+�U4̑[W�:*Yx7(�%<�zm������ΰ2\%W�F�4}�v�G�������ʐ[����t_�	����'�*ʝ�k�2�aB\Ƿ����IGe(��p������v
{9��m<�\Y}\@o0�n������t�j�F���[嵒p �~��w�^�%#��m�����0�`C����H��6��S��4j�!WQ��F��+�gA��7K}w�p	������o��=J�1`6�J{��}�ɽt����{#�lP�d/L���~�r�z��sb� ͏���ى	�P9U�%�쭈})I��dz"��#:(hL��}V�}ŃO@�&6�����:I�w��!�U�^f�F	�꾌mY�^��|����xx��Pj�A��"T�E\l�iD����Rz.��em�.{4S-!���["�iE��Y�K�;�M��6�%5}�5��>�꧴��� �k7V�E5��-(��A�cۘߛ��Ntc`�v}'e<n֮h�Q�I���BN�C����3��_'6c�{ق��G���Y]����� ���a���������u/�������
�kI."�ܖO1z�0����(�H3Qу�R�rZ����5��_�:8�=Mk=d��R ��U3�fpTԴW�q�/-T!���&�&c�#-� �P�uR���#�o%rB��X�:�e��t�eF�
��q7xvȿs�d �jM�։��R��s;g�gT=q��n�2�#i����sG�[���KD�8h��F�J���󆣊�m<BS�C��ߖ��E;>G�o��-)Y�B�`*�اI\�>A�_=�?��w#��	�{��F�,e�����7�H��
��K�N9���	�ԫӊs���m��l�m�����&��<���(�3���AZ��&�/i�pC�T�¢�s�0c!1}���;T�������~]��P2Ge��xM���04k�u��&v�;�xe��Οk;��;*�Br�ڶ��ڞԃҧaۢg���T��c�~b�⸎�l���c�����&���A���IkT飦�B����'�{xGN��������z4�%�����+>�v��_5��V��O8�c�R���߮#��a^����e'!^ia�+��"�������ы��Y}�D��H,��7x5�|>��XjB�����Vo񷪄���#Rk�L6�!/����U�b�K�u\Ԭ�j�kut#l��8�dt5zSn�:��C�{Y!qF�PB	�5��7���I�Ut�g��HM���I��Iq[WO����(�g�Y�fk7��@�=�@#
���W*5��t�2�H1����K��W-~9S�wF�,6�&��V�_�/�� (�oS�ሳx�Ǯ ̃�K)7�p�;Z�����Ⅱy_�ŷ| ���<>��(N�M��W
KƜ4Ċ�V�~�)���"�$�Mh*.�I��$.�Ӿ�C:� ��|�5l�N�	�=��xN� x���MMڐ@puS�B����4Z�N%�����_z�-�~�]ݤ��e��O�ř%�ò�K79�w'�Jz|:#ERp�B{�~l�Bj���b�����0�HcV_��~;�ۋs�l��l�$\|Vco��,�)��c�Q	��q!�3����o�3^� 	�Q��Ѧo��	���<�x�B��Ú�`(!��*f�C�s�:�J�����/���,3a�ȃV_���r��ڛ�������-���-	YΊ�l;�A6p��i�e6��S�PbPox=R�wft[I��R-I��<���$��<�j0x´Y��^��A6�������1a�'�8�6���e;�U�����-��I�\�h�������4�#��< ���(b�q7d9��%�xD{9G���W���!�r5I��ߋ�p��=�`�nQwV�mf�����s(�s�%f�D�}����cNG���`���9Ձ�#�����p����5D�[�`an&�6��X|s2�s�;�mW6]������h�C�Xb�s�n:5n�v3��\p�]kwp�6��Q�#5K�Kj��J���{���;f.��$�W����';�\$�<��� ��R=U��jE*L�1|4+�[Z��m$۱�����X��sֲ%�Q�6bXޮ��F)�+U%-���Bt߂�4��?�p�T����\�xx7:\bW���8��A�;v�������Oˈ51��X��Ǝ���
�v�	��X�`����� �������lA͐��5��{+��z�w�QZ/�L��7W��Ri~�c&�����v�Oa��(��#�0e��F��~��7t,ҞJ{/{�-����o7Dh�����?}]E�F�k:u�#v�љ���	3��r�x��T'aȅ��H'�W"�?�1��q]tq@7=ş�3qwMowJ��RE��3aG"%�#�����&��)��C��a���oDֈ���|��n����){��dG��[� �"I�3@x4\�/.*�\ �YP|7���� vA���mT} 6	�4�E������X*S���<�1s}�Ĕ��-�%B$Tq�ZEL�0�#MK��z݁¯��ԃn��e����2o�d4s8��7�}&\zT�L���<%fu�q1Z�;�YҟrS�BÖA5��=+)��0^�~eɀ�����,��j�6mo�E�\�IR9���������2��l�/�<�[�]����>����v��Ukj�1m�>�C	�C8��*O��E�(�xN'X)\�?��<��3���n�4�=�þ�یA���.�%��;ɿ� |�]�R<�x��#����Z�=�1s�q5��?3H��[�b��0�4Z���ًA��Dл�$�rJt	i��_�	~a5�F,_j��.�n�`��/��u��mr�?JT�%��w�/�����3��)ED �dNCDf���ĵs�� Nݪ�!���`C�@e5�OރO0�^���Q�W�RVO�֩l���n���0tz�h��T�?��J8���Wԭ�"���_�{
�j�^4�:er�ɤ����g��{����j��S",V;y����� ������dT��n�D(=j!�V�q.�#�Hx2V�-�t!����m�ǆI_s�LcE]!��Ob��6���6�WѺ��9p�&3�T3���sox���C���� �q2D�D��NH�[��B�Ok���B�K]j�~3d�qޟ��Ƨ �&$[�d�5p�ʈ�����r �q/#���Fz��i댊���W��5T��BJ?�bq!,���]b�ߧ5�|%�pj�*Sٜfm��5��
����lb6��bz��@��O�֩�{e9k� �'��!�J��y�0���lݝ؏ 8pk��#T��]�o�Lo�{L��\���5RkK�:�~��Jx&�(1�W�0���y��ܡ��zo�_u���d�i[���`{ֺ@'~�!�|e�M�79�0��k���̒�4XcC�����m�mzVD K�[]#5C�b�eI�"
'�Q�zX���3\�t�3w�};o<�Y�o^�.a��S�z��܇��`X�$*�[�n�R�pcQ8�8��a?E˝,Lｇ+��S���EG��LE�yÓL@p]�\�ԥT��2�vW!8d�^kNe�p��2�׿��!�԰�Lc��0�
�#F!j0/���s�CTpI�y�ؐ��ɼ��:߮PN+:�������!�����Z�X��Myj��j�$^��g]��@�����n��b�ܡTa��~�@1vN��0-.&A�@dQ�����7.9�sPD�P��� 	n,-�����emf�S���g��IF�1s�%t��z��)�Y����N�G���x�+j;���o����@�4S�t@�Kw遢K��(���8�+G���B'���J��w}Ɏ4�\bi1��Z?� �:tIG9ā�>�W"D���7��&	j���B�T�4ڝ:�ځ�VS�E�ZgZ@>���B����N-�ﰍz*=M��Ҍ�X����;o��B2�9;ӦB��^2�����B�Ǐ�/aV�l�I��|b���ˎ>Ǉ^Knrz4p�O:���A�F#�Q�1�>�L3(��#�|����s��H
�����v��!L=��O��	�Z�JOg ��m*�?͐���-ȹ�6���4KrHKbF�?m2Z���|����a3��f%��}0q(�JD 1��f������ӂ[lP�IBc����Ͳ��6jkE�#����a�^�7����#	4߱�%A�����^�P�j���ӫ�D6+p�m>��HK�[`�i��`Đ��ή���ԫ�p3���*�P�J`�)�u]�¤R���R�@NV�w^�s}<N����ϥb� ��f핚)<�/�8t���M�L��ęVE|�}2�B򫑄ib���(o�гH�G1;z�:1c����1LD�1.JZ�{CD���W�8�o����{΀�I_��X��:�[c@��a�\E�7�'�m��0��Z���L�N�V��)I]��y�8z��XOC�I���٣�mz�-N���*q� f���!���ݧ�Ӆ�;�I����r8�"�̠��(��U便�h%}����N3%d^R<�]�jK���դ�#9���e�`����ɟ�U�ƾ?�oi�'� ���/�u��Ŭ�!���6�e��:�T��@3�?�4M�綸8!�����|}����]������ͻ��g�����ը�.�o�]5����W\�l��y��?���� �&6������ߜޫq���U�P�5D:�BV��G�!Ӂ�Q�����θ/��;F,bV��.|�9q�菕��آ�3<4�6!�i�D�� e\#枾n��/������ɔ��Wܬ{���פG�M��
�r�r��p�� y� �n�xd��Zq�u�.O:X2��u%է�^7�/9��XI�e�E�g�\�)'��}|%�ŵՔ�@SU����R��B�h���_�0���?u�|�+�A&�6��}�a���,�ȓ��[���b|*x�{P�W��������'�k���,ysw
w�FD�p��ж�
WkU���-e�����r��K�L����̧��,E������ɤ�T�$&�E��C�K E�A��;Z�ɋI�����C
�`�a��m>�b��#�� ��ڌ�F(kv��-���21@$���f8��R���`L�v)p��,�h�gKQ�WjW��5�_�ѐ��E/�f�S�&�E�3�W6�T`�F�@:T�V���P��7g�n�Q��?������)M-��V���y ����204�~Y2��c� Q�^�%�>g�+?q�![\`�o4��ܽ���o�d�>C�!��s�}���e�S9����*��ڄG�m�*s�mS6YP)6]@�~O]~5ON�횜AR�UXv>Ɵ"c�n%�@�Nܘ���[�봅U=�9j���֖Ya�~��&�O�I��6nˋb�~W��P�X�}/H�R[N�=�S������]��)_�<�g�Ӵ����Y��t�$����$j=�v��I��&'ͧ�@�G:�Н��A���&��O��h��	�j��y���	��8;�K������r��8���}r��Vȩ>�/�������s6N�u�d{�)�dRߺ�l���b�KQpjg��.iyۃ>�h����	�%g��w�5;�Ϫ���,�h��5V� ��W؆ �J|�	�����(1~���<��+�D��)U��ʁ�N��9�XM�Ƚ<JV��ۓ�G��a{Άg�pF�[���߰g�ݤpH�
���m\ٱt;��P4'��I��#Γ0�����U����s�deM�h6��9WZ���t4D!L�|�Fs�iI �N.EAtu(�j�Qo�n,c�O�n�&r��#�}V��ٶ�T�T��fq���%�(@S�(@<e��/��o�y��.H�@�p#����Cg���|��Jt���z��̵j]Gε�k��.�϶�a���j���.[���>���Z�uB-��v`���}K(g��?��*��C���y�Yuӱ���W��#�<����d�B�t���$�����v�<L�s&p�7�ԙ���;^H��y6Pf����n�Ӱ�,��AٙW�|k����S�-�У�,SF��(C��͛s"�RƏ� ������%�ԮI)��p`����
����`���?�KJN}b��RXꉼ��٭v��E`�������3q$!d%Ҳq�N���Є6Y��;P`�K�Ԣ�q��Y�uP4����VYy<�c%c�
�u|)	A�g~�+(��FizMk�*$�ˍ��e�TCs=�$�j2��X�|ԫK}�cOM��S�E���?�ÂoYz�~����ÃF�ޡ�1�P��Y2m�{��q]~)������5G�%��w��B�v�+�/��7�؇-�J=�S�yV�6���%��>x���8�����(hH��%�/�\[t�&�$��s��h��lpO��$�I>�0��u�ȜۅB�K��=������$��c��?0Vׇw7�qI`X���hA���}�*$Q��#z�'��=�D��*�;� �܊4q�>�Ƌ�5��a��X�{��e���`�ݩ�Ҥ�͈���!����^y��~���zF��*r��0�Z�4|�I����������Z&�'�/�c�E;��H���c��nE}�єM3�	�y���_�Ճg��CT�8�_�a��7�,d��~�c�Q��	=L6����t�?���'A�^�]Ő��bN$ϓl�m��y�AOo$�=�lȿ����;�5G�>��0W�����|�N~ ����k��C�J_��O&�3S�ݮ��n1��Op�jB�fO�AW�]����h/n�4�rv���3k�"'	�0�Ƃ���� ͉��g����Ro!]~���s�f3Y�$q:��_%0�>(��S�`�_e�q���� ez,v����.����t4����7L�Bl���݌]A��	R�d�(��������ʬտa3��[��w�J�ϴ�ʇ�h�C<8}ۗ ��tE��3Y\������o��0��f$�Q�S��O��?��C\+����`Hu�}Q1�~���
+7�U9j��<��!��6ۯ�ea�sn��>��4;��r~v������v����J��r��6��o�A�_W�敀UB�����A]��Q1�nI��"2H���9ρ�4h���7jK�SȲ��q��k�Ȣ!/x.AF��P���iv���������|�%�i���:��:�ч�qG<l��){�HP��$�:(;��A=�1��:������(�F�/��^��q���/^}m����a������
����a��:�7�(�,K��|U�qJ=���ŕ��DB_���"*D�`�к���&JxsM�_�"��/T�j����.�X���%.��ÚOy{��`��9{�A+�Ƨ�/|�N{�M+1��*S92�{2�]*B	f��'?n̺�R�7J	`�T88oP)����1e�g�Z���(U��u�rK�M�֣5CIc�2�bP/�ݴ��S ���a{#���IR�D���vaD�(�VU�� ��u�H��oC��;� ��Mh$�n�� ��g)r�Ox�(�U��,.��i�����M7vgd������u���h��Q����U� {�]D{W���%���\tT�����TK���+9���͎L��?��j)\Whm:k�(6$��l�rDf��{j�nݧ��P�Cq���̶��k��Z~�=^N���O䫦}�"�I���3a�]5���B��]��X��E��MW�8CO̗"��Z�Jb�I��>��P{p�WO�R8�6G��V�s5�Ы�5����.������p�
O5X�Gt6�?�*R���'fK� f�w"��1b���c�>�<$K�a�1phz���9���>X�n�/���	9R��iIg� \�e�?{��Ǎ؇"�.��s�G˴����[�ʓuW�(Հ�{�J��X�j�P�QS�z;�
 aż�R�[�݃P����w�5m���C���x!��{"&��B�m����+�7 R�;R`��?�#)$�P]���6jֹ}=����v(��|[.����rR"6ty��rM	���D��}�&�ڎ@_+�$sMI�w����)�Dg��� ����m�OAܼ�9�}�"��9����muz>�.�h���J���Tʩ�k-$�j�S�0��uh�ެ�WT|:a���|�"[T@/d���ý�w߿���,�D��m��M�DيknZ=��c���H���9�ⅫѾG�X;���'%�[��m�S��#,i2T"QVŦr�kbb�pU�V���j��W3L`�;D𱈱{X�1,��h�u�2� ��J��zS�a1��ZKᜄg^5v��q.q��)��c�x7��lf��IHǦ��Dix����R<m�����)��_���C���W��`�􋗥Z�a0�"Q�gyh`L8�&n���4����k�yE�� ��ଈۢ�L��獨�Z�]�\��w?�4���F���n�3%X�#�Dg� ��
�}�E��{�LY<a�Q�&�	K��*Nu�8Ǖ�R	�SQm���ۦB\�{�έ6���d�{�V iӍ.�$S�č-�� ������V6w?4u}�)D��X)��U;*�YZ��G�5��f�51�A�K@��/���"V̒m�M�[Ȼ9��K�d���� 2��W	+k��^j��ǉq�㯞����i��t��H�X��[��"�v�F�?�M�q���$dhH)j���牞7B4��(޳�����p�88������,�#��@-�##�d[E�Sؖ/�9�4��O���Co'�7)����"S�CQ��"�!�i4��|��{�P�D��ݱ�w�]��J\�"<C-�p���F�Z�ߓ��!D�$��@�TL���W_)7�yC�p	����<I�j� ��wV��C!�� 12;}*�]Zq�ǅ��@ЕM�h�"c �[:�CR�g��Q��L��ܶu�_�����G|o�ّ칾A^�S;4􉁛�+�̘ջ��]����em�<Q
s���B�����nϣ���k�JM��ĺ��?�����P��;��پ�n%���GλF��|�J1~LM���8���o����D��R��5M���qD/�ܖ�H6���x��ݽ0?\]�;�{(N�=���@�v����]�Ϣ���L��Vo��v�ǣs������>����W��� �`}ۢ
��K*��P+9��"$��0kZ���Ǌi�
L��0?��T�xp��5C�ȢFOސOG}��;���>��`�#w?$�:�r�O�53�~ sy��Qs� Z�ۧl�R�g���'?G,�L���15���\Jk��N(?��H��(�iDU[�ȟi�3A����/������uQ"��~�M�mo.یi��3�vL� �x�ay<��9%�f%z�2V�*YH4Z&���
�~ ��ˡ��!c�ȧ�.�(�!e�ȁ��;���3�L?׺5z��yb1��)�'r��_7�E�j�q�+�F&x�sLʷ����
�Z���&Fa��1�ώ�]�M��|���o��X��#��aٮ�j%=Qr*a�se��a��ģ��e�Z
iRѢ�}J?�m+�(a��+�q�g}�͏��>� 0qKe��wh��ce�}Z�5��}��?��9U1��c����U�`�,B�_;���@j��{�F���ʙ���qn�q>�:�P	Q��{Z""��.�h��ł�c�~���'��?FRa�"!�oC[�����dB�B.�]�WϭMl��	�59����-����D))-au���m�*]-ڂj�xB����?՗dѠ�,%a�RMo-��U��9���(�K�J�M=)��U��&0������i#K�&�4F����AS�¬�4�R,�3���{����7�b�w���=�|�SS����u(��S$�yg
��w�S��-�R*yJ�4����;F�&���W�ۜ8s�/�>A�bd��0T�-�a����7/�	�eIգ?��~�A�DԳ��S�����,V$6~���qHf���$0_�.�"��r BAU4�U�����;Z��h��{h�c���`O`���)�"���	���0���.�c�S�v��h�A�$m@`~�VJ����~�j���ě�2jl�]}F���� �!�q4;34_�6� '������!�[��X=�}Z$R�e�lX�����bS�:�#���Z`yn����{���M�������]�ȞL���Rᜉ���G6���-G��fF�8,���aW�������<�����#Y��>�=n*�}���Ucv��3�0"��uk�5�$C���Ns��s�m�Z���>�-h�4�d����[$+�p������J�C0�Kȭ��LC;	��;����s{/��R��O(�Hsehw�im�.�u��k(kIS4�w\ki�������Kc�胡��^�N�{�m78���=������z*�"X�6�ѺB�����锪&w$���ڈ���'`'~�Z���4;Xg�/ d^�؄����'��3��uN���_�WE��:*8O��m>e�2ߔ��o=z��l�����O>8.x�7����z�������1�M/��G�f��'-Msgu���ҳm��@�{���Cr���ߧsWp%:G�]vM��q�$�v3��T��^Ɋ�?��r�U�X�~�6d���x��c��֧��~��ԣ_�D�U
�ۢ��"�|�c�8
G�C+k��g.��59d|�K�GѰ��%���E:�yiD�hp$��EТNǘ�j�_�ݿu�2���\��I8l>�o׸�+����y]�,M�yh�VXxD�T�\��?��d��OP�3G4���o�GZ�K�mV�brp���2v,��`v��7�+E-z����o�3 �b-�w0S�'�@ǃ�4�K�8m<��Q�Q�#���6>e�I&������I��<z�mn��܏�У��5�|��p��:c)#�1Q�4p��(	�ta�v�9V��B����wZwf���8>`��xMf _k7�F�{�V��u��ܧ�%�0�s���\�N���~��-���I���<lf�e�
�z��'��k��㌊ex���'���M�nCFI^���.��"Fo��Q�����#���ȱp�^�4��� 3i<_a��5������$.�H��P���-�yL�B�(��LgRr�X�8wJ�6��</*B�r���6e4{�����T���tO���ۭ;w4�
"m�V��s�џODS�&h��L�ܧ ��&XN➪�V��|�I�u$�����Q,�i���hD7�F6�A�2} ;qUn�I�<��y�U�&!r��!˶0���s�V�}_%��ݣ���`�2z� o+�p�sw�|JG�:=�d�ma���?[�}EKl��!!��
��x�i��@/p��)�D�V�/X�4��� �j~1)=Œ��ֵ��b��yNkȝշw	�EI&��O+����xE���/�A��B��C�12�Q�=Z��J�W`���{�/xO[v-f�	Ł$yl�]HȨ'��x@f��^��K����@�b8^��.�|��-�n?2:,�ܯ�%���^(�~��$�|����dv	���a�9�ģ���M�o}A�B�)���0�c���;�)^�|�q%[1��K���`�����0\���NYhv���j�Oa/i"39(��0B������R ����m�{Z��Թp����`�X�8˘J��Z�=7���7��ܲ���x���^Tiڀ-^ e�U�S0�3 �A�|�D���>n��X;E� �X�o��˭�sǇ����p�,��^�㣑�M�� �z�EHK\�����{m�6�:�	�\�:\ݷ�5���ܑ]��(���+��^Fm�LX+#G]���n�]T��S�}E�z�yl�{��?��38>�D��W���D �HMuKtub��~��������{�+!�)����ԦP�P�x��L��Vpy/�:�^�jS�1H�������W*��S�#��rUA����(W�Դ/ܳy�p�q��[�\�B�!_aVd��(5�������N��o3�4�!ID�{�潦օ/Y��(��o'eiL����~���&3%�H�%�ɑ?�9���y���#��t��*���:0�ծtm�Xc��_C�ֶ�Tn���by�%��R%}����꽞-���5�����Ħb���%��%k��8_�:z�}zu�A ��
;�M0;�; ��o
d�c^���b�5�wVb~�_�>]��W�`O����^�4>#:9����1��#�=|:Wbȳw��|���Ǣ�7d�m�@��k�Pk��O�h�3LU+x�sQ�|��V��DO�Yq��� �6**:dE��&�s���-[64�ȭ{�N[u�bԞ�+���x��vg�~�ݕ�(�'{�ec��ks�u�UV|_P�X�)��J{����Hi�:Y�Q��x�XВ�.�O�-2�$/TE���e��i����+k�W��H��5�KDv���6�����ϺrV�-�Yh��?���2Ip��e|)O�Kl�djR�%'k�9��{��Gh�4�"�Qjy���k�I�2%iu>�q���ǈHI�-�څi�hL�g<����+4<9���)^���t�[��.�0�Sr1&G�tev����a
�[K��&yA��DN��#�M���ue{��zш�����墀��IDu�(�'_�#e�(?w��$�,��ϴ����A ;�6�2��@����_��o��rW�I{T��8|C��|�]ګ����?|h�0�O��� �k]�0Ȳ,�)$�51�W��m������1����������I��ה��6��L�wX���8�	��U&R�*h�
�f�>���%���p"*Fv�e%��&�AD0	6�D�ԓ;�F����1��MmTJJ7�I�$��G9z�{^�'f�k I6%[W|MA�o��i�[X�����Q7Ü�����
4���D9h)���S^uA�G(�͗��Kj��o�s���ݷ�7�=Sd��C��׈)%�L�DY?�aV�?4���V-�VO� ��EBFI'���8n�!��6M������$2�mʔ�
?�j�V!:���őyO��v�!D�?���+?�'@��WD������ 2G�Ԏ�2&z��^��Ν���=X��R���*f
$9HO���6��|�:��PgJ�>���� w�]�U��+J�e&����9���_��Br�����	G�M6R�){i'E���wY.y5�������k��ʡ��Ac�hm�G~�I��]#�ã"W����x�[��RP�V 3��"�A�^��	~OM�1����)ٖ�ȋoA�c:�ˍ3��@�.��3����Į��bIW�u��5�Ԫ:��J�f�����
��[��X�m=��LJ�r��!y}N�e�����P�ҜS�)m��V����WmW�p׶�Y����stw�߷�Kf�g��'ECuU���4d�#P��X	Жl$�ӯ�XVsI.�&�T��v���b��i�ya=1L-���Y��S�� z����9�b�� 9����p-��&	{Y�r�E��_��evy�w�d��ol� ң}�Q<�"l����gE|(�>45������R˾�vs�A�YH�t�.m`\��"2��꽧eyRء>YO$����4bsw��Jt�g�p໏@���m�u)�m|�`�D�He�k���c�f��9s}#���������̖H����{�y}���W�X�B\cj�~�*�g�A�13��`���7A]�\n��.}��+�Znh�7��`��-B�S4�gX��6�f�S��G^z��Ac2
z/�eUS�]R�s��+P��IuJ�OtF�Q,B����*��Fݪ)R{��`�B�i_����������s�~T�y�%N!�xd-Hqw�˩�b��#�m��� H'��W��xR��@��?�t楲��>N��8�r�1!��0�b��_�	������>������)����Tr��o�m���	���{������L첦:��ӊ}������9Ƕ�P�Zi�k��$&��0q��PeU���������,0N�����?�ͮ�i���?����RX� /+��7��FLhQ���1�N"k����k^���4q�3#�7M�,e��ZG���W�!���b�I�+"t�����$��d�'���NZ����K�ۜ-�7Z�E�#Qi��_��*��xz��DA�N�J�k����)�$L$f,�t+��XU��I�9�ԑ�w���h�v�Nә8LDX��wLw��C�V�c�L����䠤N˨���\|W�o��s����j�俍�v�����нw��V1_��?D$��iw�TvJ�[��@�Ws��B���9)�th���QK�n����[Z��MϷCHۯ����~r�?�j*�)=��0'U&�V��}��ǎl�=&�Bl��S�~<o���jd��x�@<�9��q��{������;�^�X �M��G��ˊ'F�ܷ��?.�H"j;W�������W7�o&E���Gsz��	jm6�	J(z��f@R���y��X���g��e�'N�U�܍<~_9�"��^�z���JJ{����N覴ƇQ2�q��5�������T�����Y7�#\���ᆙ��~^h���5�o��5N5��I뱪���np�Xf�'v �������dP��cӓN�A�b�!_?���a���x>oԄ���+"�ה���RZ����M"#���G^6,�4o/�� ��������n��⟥�/7�>�y����RHe]��G�	�w�K�(��de/���~G����O�i��갥�OW�Y���lL;a����z���J&n�$"��*�y0�8.gz�3�J$UAoo����"#�P��0&u(oY��Q�Q�*O����DjDة�3��
���I��<U�Ⳉ]���o� (���^_,9��+��P��'�:A����Rt��Ң�#|��]AZ^Y��z��������X��n(	;���]'K�v�
�!_�z� M�O%1<�����Af]�Aj �^��5��I���CZ<�9�`����>p��N�m��������3N����!���y����Us��KlTɹR|��~`IH5oBL��pF��4}��b鴳�B�^�J5ۓQj�V&Ppr2�G?���c� ����6U�y�CL���n�B�]��~И��*�8.oa�#��D������~�5ā%x�X�r�3��q�r�P6�Kb�\����l�x��!�`���n�R�0��70L9J�&��:��gs�V�I���k%�I�c�ɀ������cQ��w\�͙���_��Ա^A�:	)� �B�%y'��^agM�/�|&��\8	`�KAm��m'�i�p���c��a�%1)���+�<����0;�^�v/���q"�w�j?��tgv���ڑ$����eJTP�<)�Z̼�����&������2o%?�ὐ�ЀW�\�/���t��TT~�
R�*lY���q��;�ݚ�9�+��J:<!T}5�c�?jܤ"�C���g^�٦>qɪ,�!`.�8&:3�j<��D��Zu��h�������5�shψb���T�s���ܜ(�u>������uw���u� �����W�[zAy�����dZ {Ic��h�פfĉ�ܭ���ۘ����XI�6X��.�lƬ�q�Fz]�6D�.�ύ~x'���e��Z��1=����`&E���(�v��~��myj1�	�+e�8��%��$�I�*,�lђ�7?E���$/!e�ƣǪ$)�^���s��$����շ�nV[ׄS_��>�Mʧ?}����B�MZ5	�9����_iA��S���C�-�9���&)U���`SS�y�#�yґ|*�*�GZ҉��W�#I%�{q�З��~��G��C�t͗5.z�_��	j���W4�z`������։��y��Z~�@�w;g�D~J\���Ԩ��p/ן���36��3��[��"`�1c�GÜ�Z�F�k_�"�۳3D<���2�o�5[�c\��������4�02@��q�%�v��XX�G	"���:�p'm���"/<ȃl�����`E55� �k�����q�%(��I�|�D�8ja�2�a��+����� O<�μ��$C�]E��~���b1Iڸ��upͬ�A��7�n����5��&��ʽu�[���4�4�����Q��}4gҒ�j���v<��ǂi��ޒ8�����%sdo9�#e�<և���7'g�]O�{s5�rѧ!�@N\p�O�t�6��"�T��
)m!�y�%$����S��m��n$|�k��x�y�I�7�*���d���D�_�Vw���K1�W<�K��7l,�_DN�l�t�°�F|���|O��E�f��
���,��nZ]��d�a��*��"#�/��:�*M25��y�����N-���=�{6姟l����y&ƬH"}�ٰ#�%'�6�q��X�t��{���n��,���;7�iI����_P�V��d�,��Ԍ��ԅn�x���Ҭd��zp}B�7{e�������<5o^}_���x|"� ��0�lO��fb���Јx�0�{�����J�*o���_j��5gĸ�����C|��f���
��l\�٧k�A.�,|>�y��K�V�GxЂ���?R�ֈ+;-������H5
�q,W��ve}"����=_�uO�?�u-A�����P�6ی������s����e��y ����I��d���^�� �4�`���O5`7�S����cZ'�v"(�]��E�@��;08�_)n�&Mk�7*_�㶲�p3̦C�[��L�ZOrd�&d�r1T�׹�8��*=��}ĵ*�:����Yq�W��Ö�D��Z�_#�рj��+��@�%�}s��+�P�#Ӓ�Tq�>�k��	��,g�%��xj�8��i�E�s�t�!l�3B֜P՟�vǔ�?qQL�a��I������1G^��O���U�\�hd��/߹��~C�'���k/i{o��E�A��k}��sA���M�lCB����'��L
��X'�7�F �(Y3��J���Iޚ��pԳ�$���!R"lۨ����qE�`"��L���> M����p3�w�Z!�۸��aA�yv��~~;��c���x)
qzm"Ȗ��j�jp^�z�8u���(hqJ�󋹬\#=x�)&��&��G��a�H�u��8]n���m���=��}�l� ���DY�d���l��v���-�ĳD�+�*�|���3X��CE>�o�:)i"�)�H����)WVR��G��(%�� ���J���%�ĂC�H�{d��%�PE�����r�~��}��� ��^�0��XZ�b����.`4�e�.��K����l��6pQ����n9����]I�Q&u������n�� d��/`bf�#9�t�*�	���3�r�YQ	7I�R�T����0|M�n����������G�27l1������@�~�`"���8+z%����t�zVCA��K���l�BV��1m)�H��p��Xf-�,D�ϭ�>�d@�Zj�+��L��`��xwB�῔�A�*�2[P�~kK�]h��}t�#����n)�(d�q�_䀄�}ǀ?�(N��|��ʡ���c`*-@i��)p�I���Z�K��?����0"���!�?�_)vMq�f�������0���9� x��9~+"��C��B�p-ye��o
+�h}��(i�3�m�l1:�qH|0Э���o9�X%�7KPφ�4�z�:��v��B�6]Gb
��%�L�!�}h��̹Iα��l�#A�qE��'�����u!�g��u+f+��L�Y,��j"��{̋��jN�y�G�<0fean�#�NWM	@Qh���+Շ� _�(Ӯ.�x$p�:�X�W&#Ey3��5uN�S��n�Q� h7���h�(�7����:�߂��p������z-�<�G��z��.��F�?�:�,&>�>�w�H�㷓4��j�{��`����*���&�Z��μ>�r�:3��R��{V�N�:}8�k=M�O�ܝ,Aΰc�cnqr,,�M���M�t[��'��>y�:���M�����2DjSkTD�Ӆd1N�=�bW�gR��1��/dUe���8쉕�1~~���"l�dX]�x�k��Ⅱ֗;�*����MMZ-�~s��K̥`:l�rgP>N̯���L8���b�:��jDOk5%�^Q�8�s�����eBg~^�=�)B��lO ��NS�t)����B+34'S�J��h�����Tԫ���c���
?�s��PQ�(�����~�d¯�y���0�śx�]��Ģ�X9rRy��&���Xx��ir���~�~?r��#��0}���9�+i�*�w�xY���j��s9�a�a ��\r>�/"1J8�ȇl�J ��>��I."P�>Aa=|NP��c���a�|��q9\��
p4:NIN}K�'߿]�^`$������xy+ڪSҒ��|}��{��T����#����K�/��>���|�VS�M&/�S�'c���vꔣ�?ibx)%������m��UMx��H�p`i@ֆqA���
ݢX���}�Uy̿Y����\�� �?�j��Qf��j޵��Eꄳ�����J��ERzEĺU&`���;�C$���	$�=�
� !��~ �[�*�B�+��d���Ɗ7)��/���P?�	U6��n^v�j�5��y���Ђvr�*��.���;��^d��'5YEo��L�w�3��X�m%5�g�M�p�+��n�� W�^"@�'*��	bF�i��$8l��Q�X�V��=��H��$ EIE;�T��cr�$���I�Q��q�U0���dw=�k�ck0x	m�	����M{� ��m�.7d�g��D�HMQ�G��,����?�
6��Wb�?��12���q�bݷ>��N��I�S�	���jW7R��7 ��������RF�>�n?LM�g����%f�,�E�QI��F�qd��h�gY��Hi[�2�z�]��t���5�w�C6�/����;�Ug�cp��|�JH@kN8{�m�B��D��&�ʁ�<ϋ��٠����������]�9����I��ᇉ�K����`oD3����俜�J��RǗ6U�=��~��o�0�U��e�XkYЈ��B���b��������_���+��n�赞qL
�eU��0������"x@����i#/>"o��p�F��WQ�����Yc%���F:yI�ҺZeWI6K�E�:�������gS�_�N���ت��e��hKՒ+���)
7���3�W����EO!}�mn۪N���y[Yv�o���i+���&?	距�0�ς�&i:][�z�q'��]0�:F�h��W�(�,� �5�|��,�Gڰ��.s�x�Vk�3oϭmd |��O�a�oW��Xev2ؘ�-E�ީf+TM��Z���A��>|�1Wo'R�D�R9�<' ��,��݋\�-͆E�,��}k�~�=.?���/X8��'������3T��7��rW�Hկ�IC�J��P}��ߜ�\�{��t �š�]%��7���{��F�ތ%Fp}u���x���i��FR�ܺ��A_��B.5�{���W,RI-�A`�'�=��ʛA>�w<�X,4;_�|iz�t\̓Y���Og\hg���ŏ�i�K�B�-�n��f��n&�Vz(_#�d �>~���s�M�7�~����=�Ɗ��+)��v*|h����-F��x儡yL8>�Kgu���=(H��}��=����J�x[c�j�).(����Xg|�L�Y�*]JMJ�$������������;Z#��XBvU��	�|J�Yu�x	�
�ʏ�־���)�Wy�~>��^�z7��f��sHԞ�~����6mlK5eo�-T{�P�!0���þ��3�.���K�Z���⤡˕(������.�vCw�@��뺦f!#�}G%z���!/tpӱ5�8��K-�4_��e�̈���
�zeb��<�]��͂B��5�����¥��7v̨ׄ�ߠ�����2��NCMX�b���v�)��7��鍙��PC*��a�Дʴ2��<��y�!�]�yƖ���6$>�!�^�IϞ KA�OmΉ'\�B�����<P*V���	 �|�6V�<����|J"��4�be��{���L]�)�}&���L����;�����/a����QP��?��`��p�Ì�>j�/�
���[�a�>_,��`�'���n������(�T��twtfE����{�BHJG�7OKhxO�{ss��w#1+p^�[�d�Ε�ƫ4}L�����X4R(�5Z�;5</<m$̒h�03y�iMK*���<�ۍ!_(i~��O�Xn�B��Lu�C\�?$)� ��ʟ$a瘓3�̇�X�i�M�=fzW�w�7���c�b���>��k�E��'��U���5Z5������� ��p:vb��c����q��+��д���D�S���"�1����Ux��ا�	=f���LIk����:-��-FCw*��	!���ڪ�$b��	��݆��)�,��q���*��c޺��""���\|�/��8�ە����Y_T��bEz� �^k�:�XN�f�B�)/�E�?�Hxt��I�����९����n�+|QkiU���Uʮ6�?�dHr�gj���u���M��3�9�C��k�f��>U�kD�3��GZ�_2�qM�x��sŒ[	&9�U����u�Ӝ�J_Mw�B)����n(��:�RsZ����&��ԺY��$V����Y��=v���l8s���ύ`T,�$߷t����U��H��L]_��~�4~���L^��<�I�a�(_��#�|)��_�]�tn���4(��|D�k+�`i���ٝ%O�|�oj��&�DH����V!1���w9g<m}�\�w��u���#���ML#L1��{>�Q6���U���/�m�KA(L����;�� c�����G��S�;�U%R��^m��L�2
�n7!>��G� ��B�PC�*�	P}��+'jAS�����K)#�w:˪}��twm�߲���aJE(���		�a�j�{}����cZ�rpo-���#���.M�~����N�&�|�����k�F�H��H06(�P��xgd}�ݟʞą�7A$����ɦ7w�Y+fS�HHGJ`���E���E�r�(��Se��ʽ�g��h�����[��G�'�W��k��j+-��Gǜ�}��l5ð̖�=�u�<�l��4�^7H��[���5�`�]W�	�ш:e�R?2��cI	���k����hFV��tX@����a�����2�ր��yѯ��%n��z��J���Wh������$B�TRI=�([�v�fyٴ�\�2���3O����٦��.�P��}�O��g~�p����ʉX#���⒏� ��Ei��;+����j�\^+�Pg|��j���b�h�i��*�Wp��?�O40xB�t�l������vQ���zNU�0��);���0=�J������0O���d�BY��0b��m�K��.����&^�^�^�T :q/���H3g.��a������a�$�kq��o��ƚ�(�Q��J�·���^�l��P�
�ؚ����@xo(X�G��U��k(Wb4=s@W�Z'"��/�i�)j��Z��w8S�0� kd�C6�p'z� g�|AZ˕+�(&�-FY+�����D�w��ZL�2$��Q���7����Gd��;���Q�)���e��YQ������@���#v,f�#�ȳ��s���
����� �7�9�����ؔ[���<��D�4Gۼ5��#g�/�Mj7[�O�(!:	dȐÿ�Հ�n`�?z+;�u,G�u��.D2:S�IH�	;�g>��=�MU_{8���!i��Q�6�ѧKC�?�E�� �S�G�a�����Y-�Qf��E�2=Ι͎e�(�^f�+��ә�|5���D����:�<+y�Y]��Ó����Cd��N`�_>�1���T��2yq�б0�0D���K]�!��������������=�Z�)�VlKJ�E�*�"�ٲGI�Y�k�#�3�uq� r������P�beo�$Y��U�����q��4�� ��y,fS ;[�?�V����?Z�=��\�s�aP���ue��q`$�'3G�.j6ũ_������+� =3���M�z'yL�.�+��7�_�$|J��(�}juc���!�=��H�f��5OF��f�1uJ�L���v9���gL漝])&�h���~�@$%B7. g�����F��z�U�8=�_�#vt�����_(U�)����`:.���im�^0�iJ*Qۼ�c��{a8B����4����f�݊�F�+7q��b��y�tk}+���r\�$�b���|!)���}%�0�6���a�qb�Эm$6Õ�J��� ��`�::��n��-�Ϡ?�u}C:A�2�Z��I�Ѳ��{�uu�ۗ� Qt��������b.hM��q�Ð�/B|�ȯ���+�0{^g�Z)dw��H>�y�9��r��2����ړ*)'�@H����j��V!1h��@��i�<�{5X��������sZ��<Й�5����,!��e���!}�ܔ-Z H�,�����e2B�
��T����]�i�Yd�j*OB�j>�]X��N肣�ix��U�����+�^g��,�"�=Lf����Xq��gC ��71r�	��")7̱���uW�U-˷Q�A���P�2\U�����U�f�u?w�b֨�c{&�؞��?S~9D��jYo�@�����y{�3�1Dlyf|������������H���|�s���$��d.��2���K4D�gk'�SQ����<"�\pH%�+������*���9���j���0A��R��>��� �.���=�8z=VzK�YD�ٟ���2y45h�տ�q�}�6Or{x8����Q��� ��T�	$�|j嶤�������� -�v�1�z�[xrUhl�:.G���A��OU��j�も���}�%�$���WMYc���?0h�:#D�͙�i��e<*�ߋ}*�.ȷ��rC���ҽn ��o��S��ڕK��y���ibV)$�ԥ.�t�t�,dW%�����f�sRL%��~��yo�d��^���!�BG3qEj����RA�W�o;�Jx��0�I�W&gz��1��q	F�G��	�o�	# RV��)mXS�PM�`0�44�}�~��9�e����,GF:�KY0�}���P1����0�!Y��Ѓꇍ�0����������TL�GNVhOk��Ǫ!Rz(:>�F9@��l�V��(ę���ی���Xan0�[K��I�aV���'I��y��c�g��~#�xꇝh��U�G��$'�;t�8�F�!��`���[G����_���rh�w�j��x��̌�1;g�Cx�un�I���}�N���ڇ���'�5#�q�j�~ߎnU����ҁN~(ovB$ ^��t�>���3�+ic�'���L (�h3�RY�a(��o��+B���
�e�$�k��i���X�\�f��Ƈ�&G�t�l�(ߟI�G2��N�L�"[%���YæC>Ʌ��_c�:$�wX���BK��dD�: H��H+��zP���ĸ�_	H���zWi׼|������
/#��a���C��)
<����[4�����tL���xO�5�Y��A.̔��V]�Ly>!\��]���A���f&����Ԍ�&0�����L�?oS���[�Y!A������YY�:q(�߱���P�;iK��YV!I	��]d�]�����_#2=�r=�p:{�¡�S%dܾ�Xb�Q���V{��*5N	����� ��;|j����6{m~�dׯ����8��h���W�X����'��T����Z/�H���G]c���ңx�f��h@(b�� :b?ѷ�xPБ<!���Qh�]��Au�K��,�h |�6�e��ή%dط�m��Z��ht5X�"of�
�h<w��z�I��=���ɢإO�:��i�T	7$Wf��&�(��b���#4���������]Uʀ"��>O�w�Σ�~��y�!��<&C	W�����Rg�bK:t���:�,�U ��{\��� .��YZ���b���'�ܛ�dqJ��U����� ��pU?���Qca�Cx�������-5Q�Jq(F����:wN��E,J���P@�A�:���(�:s�^�o��Uۗ1���$�`dy���3��S�V�P� ��L(�5���D&�oڟ%�KXߴ��LE�c�.��M��w���xnv����2��V�Z��ӧ$�$�xj��:�糅�$d�*�m��]��>�M�\�,Z�f�FXJ	����X��z�ԉ?x'��8���f�	o�����o��u�;qK� ;k�?pw�ܹ*��w�
o��ަ
�EZy0Z� �Q��,^��� �t�L�z4�X�_\��`]
�M�|�?���