��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��oA���C�y�b?�Y�u©;l�F:I�N,�}�	��@c����d:��W'�8�E<
��ԐK�ĲkQ���=�-a���-6�ć@L�0!b/Q gW'4��19i��&8�B��]�h�;��H��T�@��4�3>	oB��m��ҢI�қ���2k���c�G���J6<� [�}�2 �@����D�*p2Ls@��2���e�A[�2��"q��f8Q�\Ʃ	(�FLaӦ�fr���:q2�mW����اs�����#����g���^���Y��fI�E`<��ti!����ӂҀ�]��3�T[;�3�kVغ���1��_�7F ��-�09�-�1���elD����I���Ƣ'd�06;c���F$�M�+~AP
yw�7v��n�Ā���f� ���3�XC90@#��Kp"�B����y�of�u^'��2�H5Z�{}�iW����w�N�l��tiq��q+�cY+�A$g����~!���!�i�l��	.�}[���
���'p~Yy��}]	����g��ym9�v�V�:�b�;/S�e�=n^�vk�̼W�+Mu�O(Y6t2�K)]����[��H���w������F��%�bi��ɖ��^bWw+g͡�`�:�������X��ک���.�6r��`N-WP�G�ŧ���]Ϊ���[D4�r�S��
�䱱�u���9�����=���`kZ�>�2���_�\�!y����0]NJ0��%�|��	�N?A�^�����p�GE��
�%�՗����"GAP5���aL7�Z��B\����)�(��>���#�珍�=�[V��O#g%�ؠ�b��)-��No
~�Ē��%����O֧����׻����Eu��}��d����S��Џ�1kIJֹ���u������A��v �o`:�j��&)S9b��?y�D�[m99"�_�j�/�yO��Ff�T��/�ɑtQ�O�k�������F;Z��;}�.�SL�x�=�-�ڂ��9���2$��>��$Xy7�"�)��IZ���b�U�u�3�eX��"�ڕ�B{����>��г\yɃ$qFe�}Q��/��Y��"2�D3���������� �=�/�-?�(���ūȅ+���O��0րS+��*_�Pi�^
C��FpKk��X�t�ޝ�y	8�bD�:����^Z4U�:�*0���7j>��e?��`��'��LQ��onA�Yӌi�
"���{�R��<.�_M[���{�C;�ֆ��F�Ȝ�@=@+<~jp�6k����1�c9R�{� �� ��&z]�1""D���i"'^�= S�� ��#��V����Kl&�)�rr���+�a^l���  �po�KQ�Ӟfkw�Q�Ҁ�GJ�$t`=�*Meq -e�}��p�j�>����ڔ��5�fcŰ/��2"�D��9���r����o��}����\E���vw�Q���vQQH�!+/1�丹/�5��p��Fm%^��|���?��s�࡭���e��s/��/����)�~��]����yi�h�IC��J'��;��Y�^>�
5�g�!:�h�q�.~� �L���
�_MRi��G��իP3Q�m��Dv�$'H>��6EM�إ�1&d ��~�������>2���S�O�g�4번`���=<�0�[��@"�O*�y+��;Ϳ�0� �ܹ�f]¾(�}`,�^1��vy�<a	��a'n��["�|�g�-�?<��N�F�6�_��tFf#�x�e�~�H~
��<)�uƞx�G����+}h�CH'U-w�2����ܺ��ccH)�=I
��#�}�rd�"�o��Ž?��	�~#��?�1�n�>�fQ�_��HǴ��������^\8��Y^DXe�3���H�)��~O|��N���5���R'�"w+O���jd	�Ų��K�<�.)�%�z�:�����[���Iǜ����9yC�5��.�ʬ�i"+f�Tq~�vH�d��چ1��O���U�y~$Lwl�ɭ��E=kb^G��Z�X�x�ni��hC�Ϫ����o���)�9��\$��"O�7��p3��;�0�q�~��/��V<Qt����zj�pZ�"���T�p�j^N�4��Ђ��VN%�W� ��?-�>����
0ac\��Pe����Y�W>J�����|�y�����e'����N��M�����f�
�ދ��4�S �p.Y���t&��ܓ@��
���!V��0��гfp]��B��$�F�,qɹl���Ə�izI��N�Rq~*5�.hn�ܨ���m_v�t�!J���x8*N^�Z�ߡ*,ꗬ5�����Yzj���8 �<��E(��@����(p ���*���u`<���pU<�*)�����;����IЗ�������<�c�0���\,8}����?�R�7�DbJ�χ%���wލ�G�M��v���q�30�hl�W�ןש'�Qq��4�ry
 �!q,�(E��e�����^�f
�#����V�N두B�ͱmwP��a�u���ȚT>$f� �U��촇�OrrR��/��c���}6�%��9�6�U�JL�y;���"Z�s�l�3�<K�������"$@����uA��~�� 3ό��l� Á:Jp4wJQYB )���X#��� 4ƂE�ϐ��ô�4��9B��a�_6�y���8~[=�0�!��MH�[v����y[�]
�H��X�]�F�w3^���R��c�R��8�'yc�w�������0�^G��6F`I�����
�B�A?���Jg�4yU��!����G�md|���3J�N�vC2
X�0$.�Uu�p������io���8j��4�����d����5Ԗ%L�r�q�~�e��`��,�-�lq�L�zkIյE{�l��m��
��G��to���wz���W��4�Ƶ������<���L��u7�ʷ�ť�]&�P��.�k�W/�����p�hx�Tt��D���B�Ԗ�/�̣�[���þ��K����.�s8|�o|��c�T�e;�	ϣ���ϴY�t~�XX�TL��ĥ%���6����m%V���jvI���"����n���|u�9��cxj������_��sM�(}�_m�||�?6n�s1�bK��v8eA���A��VB���a���/����W/�����{�Љ~�Z�_�V� [�ܵ;G��D=Ykh��>���Di����.�}P�'����7lt����1�F�)����SS�$�iʒ;$����<6	�7�~	\B&�%ό\O`G6�w��a�4�X�~4>˛�aj��cl� *��4_�����W�׶��8c_|}��|��������
	0IC���Dm�n�BU������K5��q��^��i(��*w,�!��|���T��ϔ $�Ng�d���V;۠����;h�k���<��r��J�\-.��a]v�#jBU �$X���j8S��ȷW����3p�[ٲpd�d��5�m�&�bzV��o�$��֞67��xG�(񜳪c��N`ox�W����y�����r�峭���mK���FC���bb�G��F��k�{�9a���-[d���	����:��wB��Kۤ���Iꍙf�On�1J,������N|i�tW���!)f�M���� ��ΠhQ�\^�X��ad2ɠ0UO�=�=8��z��E�lI��SY�Օ���SR٣��O����cEH�O�lM'�.8�oi��G_Ф�4������R"��m�FX�����l�b����ʚV�`��
��=��	D�<�QגJ����/q]X
l(s?�hV���Co�K0僖��,�a�{C�i����Zߤ��P�"�K9���&��O-;�Y�=�uZb��i߀������
f@R�s�*ֲ�G�$p�����ötِ�`�T��K-���-���a��޺.3��ā�ސ�1�h@��`�*֣�C�ĳ�Z�aĲ���F�cL�i~RȱS�#*��	7>)1��N.�����ØEr��h�VM�P�8����;Xx�O�f���� �ukr����޿_���8��GFy��W�S���N�&H��&�q?RC���N�Z�iB����EH�ç:��K/����)o�w�Q0V���f��4L���ٷ���#Yۧ�x��i]j�veXdȻ��N�=���o��B#�xѵ5����Ū�+��5���|���y�r�?��#Ŏ-}�ݟ�zV�B�b����d�����H3�u,f�d���P���Z0���]�Ӈ*�Ҍ�Jg�_�.�)0r�})�4&�d���y��y2I�	���S|9�Z~� �~:/'&��庢�c���ME��;;xմ�����s��q��߯κ��T�ԇm�34D�K����[ݗJ	ت��?,~<�����^�`mu�z�����q�%�F["�n��h���ی�	R�[���'�* 	6�}����(�X����M�}���(#��d��z����o��� ��@7�'�p�'���\Fi�{��x�l��V�GĂD�
��ts�kҩ�Kx�c���?� g����4`��xU���$h�T��Q[-ލ��/ov�ԡҶ�X��f[��C�Zj]�G���18�&�Gl����K{��O����-T�692�%�>MA��k�vI���	�2C��9�l���͆.*��n�����0���s�ZtM�GAwJ@%����D�+ίYy�&�vMj�z 
�����~[IŚSP����B>	ܥ�q�&0X_̦gj��$��S@,�`�ϼ��"o'�S�u�(���@, X����S3���>P����/�8�뻏.aC4�`�^\[f?��x���xS���թ�B�/bؼ̛��s��C��R��Ze1��#~2����9r`�e�0aza;5�f�b�~������e\���j���b:ZTa� ���
�0�1�*���\��X� .pi\�76���k0ߧ*�5 �e2��r�|CI��taG���&�&TZ�t��'.��ءM���x2�������q��
'�)qf/��D7����N'��^uG�����L�s�� ��)9_���e	fk��ujr�#��)�$�	�\v,ɤ�2��=�Rʝ�]�lU����V�z�'��X���@�ı�&4�V��K�{J�Yz����%�)բ�����>� +�B�%.Z�%�{�҅��5{�Y�q#���(�H#�^K��[�n���O.4˪M�$GN�x�����}7�S\�˞��!������8�c&6T���k5��q�t�j��"	�k�vN�X.S	�>O(̢�z�`�D�4bS�ϲ6dQ�95��#�/P@���}��\}�G��ɜ��RO�]�*�Ԙ��ȹ\�#*Y��ŀp)���-����ҹ\�1qW�
���|\�W&*f�w�M#ђ Q�$�C����"9���nыOՔm[����w(�k�ԋ�6=ف#������O~���%��.�7u�-�����.T(���S�W��/#�����n㖝�eI�2�Q,�i@o���?�᭾_O�_g����*%��c��]\_Tp�mN�wW�TM�L�	�6�=���C㈴=��P?Ԣ{D��-v���k���@ �P��@`���G�3o�U������/g�?�6��a�17�(���-����#������ j'�>�dO�f�w��r�>9��B����eՓ[�s�a�{��6�P���]�jh�şPL�D<�Ñ1�sN����!�;R�h��J������X��ֺ�P��t֋V�v�_�_�̦]�Y�S� ��xG��J��204�+'ˌg0� E`-�/�N3��� �՘t�;>,sI7g<�a\�3�����[�l��9�_5��4|��!�S����I�.>�81n���X�/��S��6թ����'�+V�� 7���x
�JGaRUɩ�g�/��+��F���l��1* �CG�^W/2̀N��$��;Y�O}�*@:�Ʒ�!Kg�,�����}�?�p���R���T=�?����}��5j�M�*���!�o�(���@�jo�	_}YX��c@�${X�i��Y�j�p�H���men����ύ�1��"[���ncl&7�QZ�l�ݰy'�n��4cPʳk�%��,�zwe2�R�sq��Tv[O�@��+wX��$Adn��d}L$���]:� ��s��sl���@��9���J�S!z�l�l�oVx`]�~JD�.~rӽ�K\�'~	���td\���_#䄧�xЛ�z4C�$���^��*?嵑�l���2����q3�9����r�}[����C�ll��WS4�M�Ґ������dC�Ǵ��Į"�K������o35/�U���*��Y�-��3ꊆf��|�'z�e{����t�l�?� �x�>�_��y��)h�%�Ř�EE�1���ѭ �ڟ�iɩ�.�x��'��4;d�E]��7�#�|�9�$���3ObR��=�|_� ��m��s|#a�2=��o�o�FB���r'P����@�q�_�iI��q�T,��RdZ�Ar�c~c�ғ���N��q^�b�!���bs��0R�|0�v&�H��L��It�іh�E a������[-�l�@n���wW�x���"�uX�����y�L�و�H憡u�� ow}�rk���n�=^΃��� ���l���T���ӿ#j0bY���6G��"��Y��Z���R�L˞7�^���N�� #��*3�LA�ת�P�gy
�s;DS��P0�j�Ƃě�:w�����)����)���a�pp��<~:?(%h����,iu/)&�:���ɤ���5��sJI��k�]�1�U�fu�`a4D<c��b�]��^�k�*�SF{ێ�ɱ�j�E���'`�����C�������N�԰�DX_�l[x�/j�.��QTF��עq��%�<�r2ټ��'�͒LǶ�����=k����EeV��h�'�n-���;�C�UQk���$�\BF$c�<o�.�w��PdD����oM���_���?����OUP���҉�Y0	u�hAL~'�
#J�*-+�%�p�u/�C塠�TYV�C���l��<��O�BKKJ~���s/\,�_|�a�����+x��N@O�}UR�&� �F�
l��D����iV�VL?�/�=��T���~�}��-A[����?��Rv��^M�`z������)�؈j޻uPdѴ�8�I�|��=T�����0��E��u��>wU�\�\�D���q���ij�~���9�f�#T�|&����I�F�jT��~=�	`j|N�1�L�0�}�_ԑ��J�hS����B� �@m��f5$�����p���0S^#n��n��3c9E��%�����M����r�cט��Z
E밁xjĮQ�E8'kC�y����S6��+e�ۃs�Ni	3j�DBq��jX��6�1�-�+1���V�w�i%̓+��G��,}
�ӨvqSuF�`uHP1�hgŝ�u�)qj�pmI�&�x�W�w�L�n�)!��l:�|�
�#;Ҟ�>��>7�J�hA�`
��n�,a�9K�P!:��f��^�I�Y������̼��9���h�R�g�]ᡙ�����4Y���~�u߻L���A�"0%�g܍�V͋UZ+q����3�H��q_��,Z��1�G'�Qˀ~d�t������v�q��l��s �w�9@��9�gB�Rǟ�uL�,��pr�ʡ ��<79]Z%��/�8x�RցX������TT��v��vo��W��p0+�{a|�*�թB����<+��4�
�ۿ��r��i8()�SH���f���g	�2�д$6x��`_�6�h=�n�%���WsKD�}@�uS�ހ��:�p�5HɎl�j���m�n����E��o��K��@��-�(�}r�B_ؙ̝;�;o�5�A����B992 pUB)���k�4�J�Y���88x���&�@?޻Uk\9�6��Q��;��Z����I信��:�U\�w>\y;(��� ���0�Ȟ�x~��l1�Q�]* ��O�����[4v�������:�Ϟ�V*CD�� �}&D��:щ_�DlX�#�z��x�o�@��n� j�(^S��s�KT,H�@U��j��D���yow�7���}�쯶��X7��sM�iy
-��v�O����nV*�g����&x���#�����G��EU�%\��i�M�$dȦb����m3h&.#��ｅ!>�vs�psM�A���#khBu���dL�Hي��Kr^���7�@��o4U�e
�
w|A>�ḷφ<� yڌ8�����U���vUY�e���NJǵɜ�XWe0��qHn�\(��c4M��Z����Y�_:�h�XʓVh���8M�ǹh¾VgSit���/�AY��L�~��;>��t�$�]�8�������k�v��;�@����@�Z+g��B	�1�-�z�b�=Snю�S�.W3k=b�� U�9���F���/�$��G/�4�c��x=�ףs�甸�_=������\ص�_IӨD��,:<�c�ʙ��Ȥ��*��3��B.
�1�M?�<��lꖉCљ�ƽȲVnlq�,3��
*��oΙ;>T�cJ��nqL�?�u��Z��.�|����c{�)�U�f�,I�)[�D���A� Ы__�q����{��q�}�TzW}@��ʮ^�P�.g��M6'Q��x���}H�WXS{���;���i���)��vQ�����);7x�����}�)Fϟ�l�K�7��УĝT|��� �������	�ҙF��"�F׉�`�?Λ��L���|���{�n`�[�G��&�Ì�\^5j^�{�"��K��El�0MӸï�ך76L�!~�7Q�[�������,�7�����Q/���F��N�rj%l��tSc�����T� �b_f8XpJ�Ѧ~��Bh�p���^����E��H�A��������E�T�68f�..�M�*�h0�J�cD��i�'��܉���U@Dl�	�27��7�� 8�-�}����Y���"�r���@��!=�RݟM��l6��i]�������
�ɼ�㿫�i|�vU#��_��J\����h�������|�W,\�i��=�/�/��A���8qKnؑ�m�|�J8�L�6h�P-%��*�b{�:H�)Y����K�ã�P�c���#��&��Ԗ1K{^�7��x>1l�Ih�=�ڮ���Y$ŔI/��B�k&M���n(ؾ!��o��}U���}U�Pu��W�V�:�c"�?xb!{�G���Z'\�۬�s[h�(:Xy�[i����&�A O�(k��:B��#�~g��,�:�3�$�`Zv�R�aN�����=�d������O�@J�nO�H���=��]�nޱ�+e=��$"�W]��{z���v���e�bo?����l[�|Q��'�H�	+u�`��b���T5̇)-�Î�*�]�<ֹe��Զ�X�k���RZ��v.��7Ǖ��V�ac��)��4��R��}4(N���"�VT��~3��� Ls�6�m���,k�sZ
ލ,}\h{xx�M��DT�3�$���!$dQ�x���뀌��[Ȣ'nMUbO!<Q�P_sI
(x�YA|3ǽ�o��2O�B�4�^-!��=��g���	/��8?�%�.�p�RX�8*�����1xփ�e��k福����J���ėS�o���P����J6�z|]�8$@�?��� '�t�h�U[<�K�',�����Fr}�ـ����������O/��6�&tR�h�7���/�����a��Õ+���#$!l��3�)i���-W�
��y�2m�S �k\3�N�
-)��(<�5�������>�#�ebu�����Cy �+Qs�م�e)6���*�W=X������W�AN긗�W	3�3��b�3�������*��<��ʎ����& ��zq�`+e�ܓ	��t7j��3�TK�2���AjW&Lj�'��G�>��G~`]�C�OA�]
(�6��bГ�����5opV�ۊ똖 �W��?��F�l�CV��.K�����Q˚%��z1��_��M�ׅy��&��3�;O���չp +ёR��N�9輚N��uH���xV�n�kQ(苆SP�h����3���70��c��"h���I��q#�r`���vϹ���Í�:pK�ew��������k���:H�S>�HP�eE��*@���U
*�U�i:��(�À�6��9��������$s�1EI9����g�LS/�9�Dic+����?�D�V �|���SF7��X�	^Yaf�Hgq R��O�A`��? I�e4���y�^'��@������i8�����_E�QI���h���Q�Yr}�q�Z�p3ݣI��ӻn-R|�'���~�@�v��%�b���'�
���50�<T6`>��w��5ȰYÎ�h�$ٱ�Wi��`2�K?]��
���kA~	g�
���؉M]r��<��^=e�^M�� lP�|	���awf�I�c(�9�R�r�٥�)���%���	!��<Rr9	��X�Nڄ3����n�����H�@���o��o��K_Kf;��,!+,2��C���7�Κl���v�W�-�z��aqy���bYC��o�
�3�HfK�Az���MO}�xA�x��N��o� �q
]��叄����Z�9Sy_�xXX���nr�xR���]�k�ꤐA�V9���Y���ο�\µ^�zD�[t��Y2Uͯ��!�Ijܱ�k�o���:�K��'N���s1�����n��-`�N�4��]g!�p4��-5��.���}�_3ar��2*�oI2�$'���N*���Q57���� ~|Jl��D�W9Y����ޤ�oԏ�H�y�y�cNՊ����A��\/	m�ϦR����6;��<^P�2�����|U-��L�Z�!�.�P��O���Va��4��qW�L�Su���#�O�m�	wBʱ2,"�t�FXI1���GT=�k3�Q�>'�����
��n�-;Cv&<�6�X
���X2�%�#��s����c H苲��Y��������yOb�L��]ܮ��q����J'ŏE�ю/CDT�!�0ǆd��>�{�.����Zn�Ֆ<mH��xT�]^��Z0��%rU������>���	�0���׈7XA�o�N./�����|��5�Q�`�,�����4U�{��z�ͧ{�<�@bq:�r�c�1���J��C��ݤj� �����B3ѐ�� �)#V��V|�-�ë?�) ���X�?�0���U�*��$W�.P�g�Zy.���hP���6���+����XRsd�;��d̟���������ˑ,W3�#*5�<�<��d��/nť���A^T2B?��@�9��7w��c����� z���my��X�0�7Inl����"�C�x>���Xye��}1݂��{�3a�Ou������:�c7����$\�蟍��d��')"?�Tn�J�A�4���;v�7R+�J-�Ċ���tr=X����9TO�w������W�xd�^,� s-LD�JH�Cvmda�x�\��n/�M9����9�_R|��O�����0f��%�5XھP(��d��ev��޽��Q�H\��i��Ƹ�0����@�7��N.(�X�m�r��e]�&�z\��c��'��U�Q���)�Lm����K�i�TG?z�l�⣯P_
:��)v�R��Z��;�}g�ϻ���̳��>��8z|� u�Ӑ��+��'k�>!y���Uz.(w��8��_Ed��g?5�����%�ჵ��k�����F��Ft�ẁ�i������躺B�+Lȕ0`O:�F���߃�&@��l��I����⽗�n�����!fJ�e%=CH��!D5�5���
I�'ϝ������mH㻧��l]���M����Y�@o��e�o����������e5�g�4x�*�~RS�mKNuYB^�l���؜3E/��L�`�^[PP�1��7m�Уo^e{�Hi�'e�J�Z�/B��؎�V�W9i���
1~� Uy@gp�o���f���A�fO)�ltX[,�5�69g�9q��_���}(' ���1Eݍ������쟺����)�݁���tCj ���s[p����GE�)C���Z,�?��濍��.�ۅ��$����6]n � ��7n7�5O��)�c��0�pn�L��W�9-��Ps�[�������
j�3GBh�2�:��|YE�6���g��r���'Y6��ֱg�+�A�T���R�"�Oc?NLm������������
Y�n4�U� �>P0��[o��̽!N:1.JA"6,�?W�[s�(#a�Uc�sDB�nIK�ʏ���x���lr�p��Y{)��<,L7�F���x�B���(��Z��Rx�z#��H�K�s:�P��j�;��Tj̳=rZ.�I	�( �Kp�(�s���GV����!/4?%�K�4�������w/�E�7�1c��RvE���J�A�7�1N��߆қ�e83�o"���
O���]r�M��	nO<k�ڗwE���T<���*�$Q�T�8e�7�������8���]���]���q#�������.�$�x�ip��?Y1�G4f�����X�I��Cb�^%���#f���@-�z���`X���*O��ؕ�k��?,6]<���4Yx/�Ѡ��#�څ�������ʻw�bnbg��@y����\��	7s�-�����2s�ƴ��b�M͛��@1K��1�4x&20};�g0�t�&��PO/z�b<4�$�Q����b^rM��B��:�5KdS�|+���k�Z�9��2������Ie������^&�&�o?	�K�Fs|C��R��L)�#���7��?XP��T�ݚ��*=*�L���n{׻P����J�{t6�u�or�r08�e<Q{���yNZ��e�T�������O:P㕌14ކ}�� ���q�@3{�h�r^�>yJߞ�K�ݝ������k�@2U�̂=���Pc�2��c	��Dҗ����A���.^Zn	�D������'�bB1t�n��W��F ?21���Z��^i]�C�$��j���1���Y�8�S��>�c��2,&8�Ј#:n�I6.x_��A��wvm�I�F	��ŵ�<�l�]f��"�G�����B@��-i/I��\l�׃H����ĉXҜ�ɸ�M#6}g�Ed�kX�"���T��7��
>�3�h���M���1"�o\�F��s�?��6�lG-��ݳ��K|l$���)g:K���z\xS���2{����5l�8�^��(���9F_�`X�㯱������R`[p��)��9�k�uF�Y�Ϗl�=�Rs�W\"��o=
��!(����o�[�'� ��� �^5A%Uj_���<e���,q�u^GL��}��e���ʏ��[��鐝����i��6���0��"sE6r�ř	����U[��g�|�n��&!yOD����}~r����n�S�1<mMxhg��0hU��Y8�J��0
}� Mf O��z���;�A'��1zۺ�F�;Ĳ��eH�?�0~�:����n]��;�����$˟�dN:�*��S�uz�6��`�}��G�W�:��&e�_����/��f��^�2w�Y!_HzB!�!<��I�c�d W�c��$��xy��-�Ê�!~ �36u�'2�j)����p �D%��7*.����7`�Lx�T�1�8�^�°r�䍋ǡ{��gB`�C��h�C��CW����e��<����ba�j�9�	���a�?�O �Ek�r5���D_�@�1]D��@$P�r $&j3-�+�P�_�������A��y��O�ɚ>��fLv��Х%��z(l�� ]s��,ݓ��^�+%� �(+��:��\�tY���1+��q>��n`���\
9n��}"���a-�~��A����s-f?�(�L�'��)4n.��Dm;�溦s���f�bx]��	�~�aL]mڎ�#g>=Z<]̡pqC����K�;�{� ���	���K<��`>�K�&�0�r�Ԑ���L�e�v~���Tl�E���J�"D3����1~���瑻Q#�\��[2#�')�Zt�}۠wS*[��$4�܉0�ؒ5_E5�)�� ��3�,&I��d������|�%9K��D;� �4��]3S���a�����W~,� GxV@gY�H$R�d�-G����Rz)��̲+kB$ӮXS�������l�N��0���H�l���o|�,l��J��g�U�&��Ho�3����|I
HƑ�B�Y�3�0m�>�~$ ��z�I�h�1��Ì����cdz����5�\�gd��3� Ϣ��F�U�F��M�;��n���33X��7SQ�x��š5��q�)�H��w�1g�ki�M�#��f�0����[����Y��dY��:���'Ѱ<��]+͇Q�̽ #���~�7h�l %|�0@�U����1�h��Ҽ&�/f"�(j3i;��N���4��4�1j��wG$s�zI�Ú�F|���j8	� �n_�i8�3r�'�k�ɘ�� �N�Q1��}�l��Y��Z��擃�nY�P�a@����j��.��F��M<�:�E7w��Ú��4�Ӄ�˴��j��>��g���w搉l���J��(�/&�s��3q��><�klx�)�q�`���? oU�7�E�l��n�u��Ѿg�R��W��>3�>�D �v��6�ʹ�A���$qU�hE��ǳ�	.�W��<n�����G�(�ULJ�:�f'&b��W���?ne�J@�{�ފ�d�6X��a�c�0�5g2�6�K-&~b��u]&�r��>����uQ�2�!�w�?O��=[�B�t;���z��S�3��t?tk5�Iǟޚ�9��b�ST�Lۗ:��8Luƴo� X��]u[\����Ġ �p�4�eL������@�TW�t�O�D+I���c:k豔�#��<�:烱�a�ZO(��Ǩ7��\Ġ�;җ�Ϳ~g#���9VrS��Z.f�A�g��M&��Aǡ��ٽ{��^M\��*�5Q�c��0U�G���`�˛�0֖K?2�㿱g�L��~��_~����Q��i��<u伏�[��xK{iQI�I��������@N�΁Yd�¶,/���ױ6՞���s�ߞ��l�E��>�A̼�_�����Kj�լ߀IH��J���|������ ���̆t���	K�U�Hd2��C���?�g�ޭ)N��l3":��ll����1�;Pf�R�WuH!�|�U��m����T�;�l������V�1tH��,�� mEwy��<���$��D�=�i¬�u�	��[5t��Ǉ�v�ف���.�5h۩�!���g�!H��S�� �yl�2$�	I_s��i��p�K�Ff�I���4,*�����O&��O �c�'�Y|Y'@ 3^I�b�9ߤ�\����/mS�Ȉ�H�-	�|��2Hf
 ̾	)Qo�
��2���I��l�����qC�������r����c�^j)�]���Fw����DB��O� sO̍/�x/]�Q������~��y|"�����r4߼��[lQ��b����6}+�qKP1��0����lXi��,�ݗ���)@������"��61!ǘ�&���������7@����HA0穆�L�kXL�9ဴ�%Æ�%^$w�x��/ب�Xb�<������-	p�T[���~�F!{�)hS�|���sSҤ��V����,��k�V%�Ʌń��W�ۙ�r� ������Š�X՜Nt�~��OI��O@��-Ql���>5$�OM7��*aS�Q������PUE$d^�8�_F��:��#�E��K�q��]Β&L$������ɜ�
��+>�q�Y�U����v0Z�	��@��cչ
{a�c�d7@�a�`y����Ó\�H*���V&�g��[j���+���S���o��s�x��IB���|���3��c&^�A�r��\S�W�+�l���e�ViX�'>h��*��?mm=fG�cE�� 1(H"�Q�Sֱ0m�ҽс"W0�ҹ�όR�z���-�V\?����4{GjP3jľ[��$(4�D��])u����d��Ej�Vp��o���m���
2���5�NOQ+�=��-��J��.`���2G��	���������W*$���7+������WJdfέ���W�����Яv����1��m���^E���Ģq����sb�e��KL�(5ƌ�mL� ���Ѿ+�P�?��/;�k�UUpovǪ�J]kv>�'�� ��.]��4?Z���M�	�;s_��}M�\��gN*���#���Uq��>�o������Qa�p�g�6���Å���vJ�'mnNG>��{���*V �
��YI��M�k!�i:2��-s��;����`%�h��=���2�[����D�i�9E1�����tioMBQM��~Ξx�sYY^,�"�(L7�y��Ƿz�������������D��oF��oiu(���a��mG��Ō��w�фh;��'��,�[����l]؅�VF�$9x��N� ���y��xj�8��g^�f�ᱹ]]��\�0}SJ����.08f�?+Ɯivh�x���N\!���S�=$��c4��~D	ޝ\�;\�ŏ1O��zRQBк�����;7F��k���`�NRK6XS��^G�1��07H#�����d��9u,~E{Jo������h�+L�
��ռ��ѳ��Y1s��[�����+�h�D�S�[qV�B7�1;d��lV��h���l���r��Z��V�hS`wp��9L�qL��
��0�?6$� ;�����\�{z�Vc)���M[��.U�==���iM̊�����v��Ȗ9��i貯a<ae��9oˮ�8���՝8��0�(`6|��#�����y���c��%��1>x���p�9��!3���`|+����^���\��AF��5Z��]Q����Q�i4�A�Z2�i���f�r�3�]�����NM�@w61���?}s�>v����'bZA}��r\*]V��~�H�u��rN��B	���E���f/��(����	=����%8���T���W��۠U��AH�� ��ޕV�� - \ƽ�E�Y#ߡ�˄J]?����Y�&
3n��=���Ĳ���3K��@c�T�i�Fi�D�r.�z+C%R\ߑUpS�sQK���UePRRw��E���U�r�@s���,��h�0uXu�����g��f����8�LHB�C�ɜ��������ҿz�4K����Y��C����HX��0R�̚)h�����;�B �w`��8!m���`�a�+��F��$��9���e �zFǆ����L0���6a���6Zq�	�"sH\n�_z"p}3Ν���k�=��8w?�Z����	��7��9@�W�4�m����#��]����Lز�P���S�0	�k�w]4� �F�Y~ڿ;,�k�7Ý)4��sY����D�Ayk�<�D��~�"���TτM�;'o�NHK@ׅ������w�3їVJFh�?2 ����ՙy��T�G_#�5��#����Kp4>��ɠ��iM2pc]W�m3��Q�U��>S�%� LC�{�`]�/��0ңx#h�]�?�uY�T���3Gٝ�J3�0��AI�>)��)ǯ���1a�k�=��wR���r���Ę:��z�7��5�%9���d������g���Br���ݫ|�,1��J^�N�✮�W�/��5:��Ѻc���O�5$J�X�ask�������ƾ㼞PF͟@$L�.*����0]"�a(��ۣ&}�iX/��V�j�U��|���:����K��̧�	�0�_�i_2ZW.�t�Ox�e�f#ȞO���4ݾ�u�~�����Qj��ߋ���ۖdn������M�Jʖ���;Fw��k�s�?&��c��賤�uW?:E�u��y�
�!���(�?@6�tY3��z��k�'4i��*��K������\f���@\����8�Ɓ;T�m;�v�*T�� sC_�Z]�k��,v��4�}m�]��b��8L!�N��Wͣ��*T�"�}�b~��^�"��~1���N/v� _�20��ip�P�ʳɑ�'�SZ�w�>�)�H�.�����A?:���3�u�J��� Kc����1�5���bU�j����se�	�}g���Y^>�n�W�K"Y�0o4+iq=�ݲk���ک�k��ќ2?O�r9y��ζB ��J��p"�	��WH{X��R&=�Bݣ�rfb���	L�x��"1��C��;�1���)�H8�d���!c6�̂��mt��I�]����q��P�c�ƍ�:���$_�6�T������:5�.U�K�ݲv��?��G�YF<XȴQ�d�������U�0���覎��e�Q�o�f��Pgm�GXۀ+� =���G�-����]D�wC����H�_���~+3���/H��
�,w�~p�=�>��U��J��"���t�p�-3��HkB��˵x'�~E��!��r�H���Fa�pǬd����J8���#�G��-�y��6 ������p��^���0I�UM��N�M��hh�6�J�Ǹ��u�I\��ly�p?�q�%����ژw��&V��p<(��O��5�/W�`��,5On�v��ng��C���PU��Y� ��W�� xRzH�tQ�IC�D;��~�`���L�4R�Ұ�抎k�|���b���,d��V�TF�y:?���õ�4���e͙��fʢ;�Lj!�_���)8 ?�2iz�on�01�h䰇��q[!G{�T����gx�E�����/≢+|��,Ը��n�A�)�|���|�픘&�}𕿀>��iJ�L}��+!��Ql�����l���c��B�>��	�<0l�'!�j��+�T�*QFg>Lӛ�C.�+���tB�Jk�5)/��_t ϫ��6e	�ɞ�l��hx�Q��o#��Y�j�-9��2�I�(P��z
��`���pCâ�}��h1nS�[ f:��t����9���%[���矙�%�)���y�Ӷ���6�f�ݨ�%V�H��b&Ǌv0;Ҩ�c'\�;Q�zV�x�OK�R�:m��1r�(	�w�\���T�8�Mls�@`ZP���t<�{}J�J���|(]���< u���e�*gCHԠ0͑Wf����mf�"����;�MXw��5?��Z+�K�#���hO�h�+x��ERGA��eU8���l����Io�S-�ݾv>tI����@�o�n��Zd�6��VFD ��C���+��`Ū9q˖���v܇ANxr]�>w��	־*��h��hX?^�f�`�p��|��[g��X��b?�,�f9����xލ�_D��N(���I�r�P�^̇Iń�t7(���.���������b���.�1�^o�R�I˪([<d�v��G��|/��)�r?�_����T�A�Ax� �R�A>X�nO�:y���5pt��� RE��jz�c���	�;`5~��(1C�SA���D�(�Jn��ݶ��#����T8%E?A@���zU�Z�wDn��D)��k���b�m`7=.`~Ҡ�>�׽톛2�_2����j����C�&��l����Vio<��
��}�����Y��TԒ�g3����1�<��'��|��ĺ�z�FL�h�	�d&��/��k���xjմ!�9☗pE�����5���3uFO�����;�3DH��<]Q72v�#Ofc/�1噦 h�,�}�%!������/u������Ҍ3Ggd
'qR�5�;�Z�n��q���?�ܚK����A���q�\��M8��U�z-�kƨ�n�5 +2r�-wj��	s�dW��+���ρ	��	�v�c"A$"�*X��IB��L�۽���Z#�c�R�An���Z����N������\�3���d�8�E9�Y)*��N����~� �$K�c��qOϿ�q4?j�C,�������_�6�����Uc�L*\��R�g��]��0�:����H���������Cŷ��l���Gc7�v��I���`�w,�0���/!8�����3KK/l�Kҋ��l�T��~�j3r���4�r��~�:�