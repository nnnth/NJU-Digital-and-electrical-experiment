��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]�����JSD���aV��F!:�J�D,�$k�JXr�}"|m�z1��!� �*�^�ϼ���_��
}O{�����'�.#I�b�k��(]��e�, ��y��_SJk����Is@��;%��m�P�c4�u��3%�4t6@�M���0���w��Zk$�a�J���fq ��V�X'u�"־N����ŗ���F�,8u�>mRfʐ᳎��O�&�NMPFM�*�%"t�#��xx�g���y+�U�2�W\�n)��F�N����Q���O���0N�?��g���poK���������� ����x�a��!�T������Q�^"�j��TU]l ;�q�鱞�����;轊�xN�eƙ.�s���������f��C�����F	��M�b����[9ѳ����$��}S򰏔(=t8�f�E������܋�I�7�P!��\<�C�+�F�Ch�?�k²��)�K,Q�	���������b����G��RF笠�UM�Z{��Q��/-]\�'�6k9'�s�������x�Ol{�|��9)�;�5g�-~9	��g���33ϩ?P�i��N��%ѷ���c�b��;�H:����hߠ|�Z��Jࠔ6�P���J��;'#�>�r�z]BWIgB�'R�*.��p���)�\�dx�I�?�1�Y-*��J
�ͱǷ��U}�pHgW�;@�9�F}����j���@�=@�~_��!������㦊�P�#��h�DR����o֍]��)������{�	๟nQ�����l�[� ���~�H\�F�����?� ��e�.f�(���{�Ip"B�`.*��I��9��9
���׫T01�q�%>f<�u=cd���M���ߙ��4�pPxK:�x��qE��J��д��d�l�A>�����fNd�r���>y�+�jźґ
ݨ�% �D��	�����,`#gZo�����kK�`z�%��ͫ�MM_>0/V4��`�����&�-��6Z����I �+3�ȗ%����%�O�:�RO!�Y^X�n�v�b�T��׉��ы��Xb���4^r�{�BB�$���G� >��D��e��Uq:/��mT	D�:C�g�R�#m�j��1h����z�9tu��6�Yʯ�*N[:�;�
��j�T���kkQ�M�A�MBQ�ֈ��1��G�Է\��z�g=Og莻b����[�\d?��+��5��Ņ���R]�	Eb�z�%cR����G�-1u� ��|N�p�]����A����a�M�_0�p����yzX���ü�Qє��%�O�E��@�D���,:]dܨ��;��x�;��]n��m��ΦZ���b�q�W�����'� y~�݀�$� TA��R4S��+�|�Wyz{��D�s�Y�O-6���/��$�d�7�}%���`P�b�(�RG���I�j^ʒS���Y�H�Q��w�tq����K��qIzD�2����T�h��\{�!����
^�_������	bm���&uvd����)�	w�5��M�zPl�B�|�JlU���5�ݢd~��	{�9�u�B k����X':�
�[wϓ�#�R��r�?ߦj�2S�q)��
T���G�k�g��ŗx�.�J���9\�c{(ϡ����^�s�,W�%>r���w]K,��#C��?.��X��5��:����˪,�� ���NG�.(�����=5>=��k��_�.�r�(�ގk':Qb��D�`PS�X�`A�(z�'T�皝@r�f��������jd����A����y$O��Hϼ�.��(��ԝ��6,7=0ub�:��K�|@4G�Z�"��֏b*���>����&��թ��v�w[�1 Zo�m�.Mh]r�f���2f-w�=}�+ڍG̠i\�nl�:���]���_\b6C�ﹼ��NC<��&�jp֫��y���<K�+4��p���M��T��X�afQ�ph�m�)M�Pf