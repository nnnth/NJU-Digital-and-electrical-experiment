��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��c����"3�t��%.S��T.K��8m0�Vy�[���
�����)rǮ�7w����اޗ�͖�_��D�-Q���
��	���DoI�4�{m�����NUc��0��ѓh��ǯ�5**xb��ŝ@����)Z���t�ߡ��y�!I��ulz�[�I�q�)�_�O��j�{�m@=��<WcZ��[��*C����^�����p�����.X��z�'�G����)�~n�1a`���靺��y��w��ȒW�T�1}�W#7b�~����8^��=J�����{�/i��5%Jg'!�rw���g�wu �P+}n���a�;�9N�I��ۚT�]M� �,$�шI�0Gz��)e5c�����R��E|�X���#R �ղQQ�����t�]˴æJL���1�o�x���D ^!���} s���ӣ$�E*F�~����a�k�{�v#���Ԭ� `�i¼�v�d��c�+��B'ir�7�ٞ�w! �zr���`"y5H�İ�G��&��f+&��'�Q�f��M���)ttm�$��NC�Q'�O�)�1Z�ˢEI�H�\!ߞ�g ҭtEuD��$$�ж��!���M{H�2��B�F��=־��#���V�~gI�3�},<�ѡ�=u�]�l��Gʩ�)��ͨ�`�%�y����\o����(E# �� ��g�B�U�?�����a�C���
y��I�sC�K �)��a�&Nx�P����*������5�C�`���B+��d�����u۠o[o��?�5R���^��@�+V�=i��7ڝ������,�Z��M����f��qF�t�<j�%U����T����#B���oj�Zil^��+F�
M.���>�y�ȝ����w$�s`�4{�JD�=���.�"rV38�
O�R���5�=�o���!C��Et�K�|΅����H�����
t��R���Go��e�DS����h�(�u��ufQ��n\��݄@��/UV�P��L��')����ɟ���m-G��M�
�-?P�)r�Z�m�x��N��j�Ő�������C��_�U=*��	H߸ʶ��e���Q���Nf�1;�u�{�Kq!V�ز���B��S���S�Ѓ�.'���6|�g5l|�WJ9��`! �"^Z�����6O3�-��x��u���~�q�4l#��%�d�O�.G������:NF}��򿕛�w�fꋘ��B���+��^��[����� e�ݢ4�==�/>K?����E��d4�w&���]�(�B5���ɞL3t��|:�a!���� �#*�>�s�ʎ����W�V����h�3\9�@nyR)v���L�.A��� �<�$	��% ~Pf�<�(X�r�>X���k�X�̡\h��ݖ�[G#6���H���;�����E/�4��!�O��D nK�n�wU��^��vJ)��/���$hW�,d��ȯ�p
�$�𛠬2E��h��׬[<���-')h�����[���w;*O����W�Iĸ�c�g�RKD�����vB�'��F� �I����=�Fu
f�3�A� ��H�(�!�fE���2z���~�|l0��A|M*&]�Tu݂�]h�V�;�x�K�=��F׍��]����}	�:2|��Q�B�=v	�Lm�H
,�M[Q/�2#��s�n�z!��`AXEb�a݄���GX\����4��H��%@C�֜���
�(���ܫ�2���b���)i����C�h�DU23���FV�<�w�R��L=��{D�i+�u��O�{iG�
���`W�ؒ�}O>RBEi&�4���
m)��	�/�j�픟L����n!!�b+��K�F�^���0v��7�N�x�v�ݠ�%F�XX|��"�.�є>ec�E����$^�$G�D� �}�&�y6�e߮<�mY���/��K'����Ko/͙��"(J���n�$�&���o��Uq�jnc���y�7���Ih����%��⟍�m�~�Å"������=�]ʯ���-R����P3�t�5H��I�6�|��(��"&5���s�P��TM˰+��Q?��@�[p2�E=7xi�}��p:;�ӭbj�%�&�j�_mۈ�f]A��o�������~�q�5��Άa�� ��",�=�NŤ �绡�N|��+�S��Z��!�6ͳG���ç�Y*��șX�ԱP�IJ��A�-�%��P��D��&�u����gK��+���C��L7�3��$���zu\Yܰ��o�{�[V��Ìg^|�o*�|��\�ySI�������N��Y�L5�ɒ%�Ӵ&����ϩ.�dWegO "J����];a��J��q7gk@��ܦ��luj�4[<xv����v�rl"�����]���#�Y�� ��w��0+?����?��G߼�I*�i��"�n^�:�͋�o���F
nSqn渠�p���@�`���h�h�Y��l�[����^�mf_
��gy(����R1�+�	����1쮐o,��X��ߖW8�$��Cv��F��UNV���f15e�6��7��UyJ��q������.�X2��<)y��ƅ0�;�wf3��������r��.&T��\r�k=���E�,B�5/���_�~o��r�gez���xW_����]&a�L��#�Y��t[�Y�r�6�*g]m'�ȟ���A�@�j�t�t��u=�k�|_f1aq��k�)-a�#F_���3P�>X�-��9������i<1�4>H��g{������o1������_L/��mC,��p�g�c@A�BRq���#[:�=7��t\�Tw�	VH��t��f����[4lb�}	���m27��0��(����*/�6�Ia���0��]R�[�U�݀���d�y
�8`��|��;�By�wK纗`�x�g^B��t���f�1w��nh�VN(e��(t/��s:E!lE:Z[�9&(�G��|vT�p��\�l�	�Ի��~DlW���8�n��m�h�6L��9��UsI���������Rx������p���WH�;0���x�"E��P�y�G#	�0edl����j���QN���;�D�ǯ��%,��W{��M@��Q�*ԥ��,�~4�D�DUh���
�����+22��>c���ub�}�0�Ţ��˄�aC
�d�ܳh����k��!����}�D�C]��Gi���?S$����?�nT"�^]9Z;����(�܄�@+d_�t�>9눋4P�:S>۔��@��=�5�G�;�����f��)Տܩ�J,�E��O��u�i��&<h��TS(�A�D�^�D�Vr��Os���Ae`�y��zmBd�09B�/��l�$�r�y�~��g���&Y@X�!*��6�::�Mӽ��L�&n����~<�T�ޒ��v?�Z6ɗ�\!���Y��x�Єu��ޚQRcWr#�j��W��q6�"vIl���ѧ�;��"N" $Α["�fe�b����^K���������~�O��'���}��x$®�V�l{�_Ư*��H��5)��e��W2]�d�48J�Ԁ{J��
����#���º`���� �+�R>p�W�@�+�1���R��F9v��ƶ��X̖>反�=R���Kߑ�QMKd~ [l4�S��L�[5x[���+�a<�\咸��-8O1Gχ�l�b^=����J�\�����r\X!І������d��)�0�O�V��;��|l(��l_�Ln|��0��+5�6�Ž�.c:�����E�<ƿ�,��2F':s�vx�Q��z4<����{��Pbvo+�Y��[(X�(�]��2��l����o7�&�Zg�H����@��\c�ڜ����S*哗.h�	Bp�5^(�Q� ��8]�����*�Z��_�rB��l\N���H͒�B �?�䫶d�Y�8^�U�#���S�Y�[�'�<��A�I!I��`n�OjOb���4�kZ��d��ry	�s:DMDb�B����7�ߊ��o;�Ղo��ʟ��cP�a�U��i�Y��^��B^ԡ�G,��ڰ�&��P�VR2+(PU#��-��Q��%2w��fA*� }7���2Ŷ|*PZ�XCR+Hhk[$�4�N������%�[�U.n
U�@vNH��@Jw�5�/�>�r�!qT�|B��;:G�	5f� �$V�v�IV]�����)����N���?�؊@"�B���}۠���J{���v#xT��Q״��3쬙*U�(�����V�z��iT'�.��|����A���,@�Nwcz�b�vh��\� �Ԑ��ΰ�L\xԀ1��a{l�VG7e�a�y/�C/Xȼ�RLR��p�?��
�^��<�>�j�	����1� c8�����F�6	�d�x��R���0�}%ȋ^P�Vǉ�okk�F'k�	v{^�px������oa\�Tz����AB�}���'�>3��^o0��2!J�&~4����P��,fY����A~L��n/�H��M��+���g�
�4Ҡo=�l�i�~��NR^�{�6���*�nM!�I|��w�������aL��۳T�Mi*�P�܇ilO����PLO��&=`_�����p�"MqS��J=�9r��"�fK%c��\Z�\�2Y>Wu=	YN_��U�q#�� �ޝR��ѩ�C^F'�9cK�[�ۺۚ�;��(���ZJ�>m��E?�Uw2�Q��)L�����5Tb�����[i3��ޒ�����Y{�x�?n���М��y�=I���Y��Fڤ��ם�y~�
�D����Rb��ˑӷL���཰�;�u��53�?$k���-̠�m�$�V�Y�A�8��)s8'��C䱤��L�}d��2��$�3vƖ����m4� ���?S ��<�a����A`��x$�_ocv|�^��=��9������9 
kH��M,�_��)#Ѯe�v?T���zF�;�K���h�ER,Z�f��}�ٌiC]եv��!�)��yG�;���%�/R��%�yv�Z��W�Z�dF��Q8�����Xe^�� ���EZ�lդ>��4�����b�s���{�ub�VF]P��吪g�39���#$�{��ބ|���0���x�t`Aў��םw	ͷ}p�sJ��~��x��x��r|���,���"�]�t�E�r|��!��R��VB�QQ�w-�ȿ�߯�F���Y�^�3�ѱa��i�����?��]��A���T!�jD�<�m�51��&j4H+�����<	���S)�=0�����LC�h7Jکn���s����u�Uc�'A7�/�픿�HY����{�9W��w煄T��f����V��l�����f�NmQ��y�e�^��0�A��,�iH6:4�;枈0�-������e���6|�~<��"�I��j��]lh���+o�΂��δ��;"�	ׁ�y�Vp#��� ����j]�Vb�Β� k.�Zި��K�����Dʔ�k�I롾��||��-PشG�X<y4`+�K���=\r�Y*����hO�Ȓam�mͶ��h��%+Vm��)���'���q��u��ي?�q�Ts���r�{0��R�����y�]���zfz���<��gܬ(�L=���R�!o����A�tߍ뾅MMq���5�O��-�WItF�Y�b�B�]M('Ò�?�J���ҍ�_
m���b�ҍV{`��L�mfU��ŀ�\�jC+`˒g뼾�o��T��$����Bů����ݏ�릎%b]Y��9i�5ؾ��0�� 1�'��&���m�`�~�	�̘S�K8�hlDg�W��0dU>�x�kh�@�{��9���H5j��S�@抡� d�b���r���L����� ��i^���{_i��>1�W�dO[�
JC�me�Yk�vU;��߬@9�B�q����h�����g�VR��A�#�2`+��\n�ml��Vop\Gg
�i�A�x]"�0_�S�,�h���2�Gfu�-��g �%v��/=iOQٚ猫��Ϥ���AE�-���f#��4Q�A�CC��C��b��`����v_)'<!��m6��י	鰩�6��Q���WK��"�,��Z^z����|����}�����W�,��Zx�%R�X�EAEd>��5Cf��/�?��v�!�#v^.무Jnk����e3��j��}���u،֥Δ�G_�'J��BpN�3����w�mje��g�:e�F�`�u\���G��7�D����޳�ݠ�W(����'�4���Duqii��K�w9�&�*��������aq�\��Pc�f>֎[B&W�Z7����a~W���
2���F�Ҵ�l�J���5�f���#��YD�p7�5�Ydt���x@`|d ,�%�>���]��m�%��ƣ�o)�ГX�K8:�i���X�Bʴ��ĭܪ�JΚtiܓ;��a����~��j=�Iu+��\#��_W��gq<�~�c%�7���k�1R�<�� �UHqJX����K:�<��s�?��-1V�" r&�\�A�~M1�0�m��vxzܮ�6�4�]��!Bʻ�!�7e�C�sSD��2��P�ӄ�9E�܌���?�߁�9�c�,�G٧]=����'(/n7�6Z�f�7�������7ua!P�D��F�[�J>�@�䍫P? Y��CA��AmK�Eޮ�u�{)�	� ��?�ێ�f���;46�%���Y���K}/�'e������K�����ъ(�~5�EV>���C������r���CAO������4����%	��a���/��z��
T^^}6�/��Jp~qE�A�=m��#3��-�n���hS��"h'�dR��赾G�&�*��r���D��N�������&��Ҝ��w�4(�!��ťAΝ����D�|֝�Dy:4��>�2�&wM�-�H�%�_��T�� F]��=�胨]H�5h#e �b�]@1�)|^X��
��I��QcB2�����3�)W�X+�m�0�ʸm���p���]l.,�f���������T{��rer0|��S��R��<�x�;Mɥkt�>�X���j��zu����:NI��&�֞��9�=vb�]�	V-�ޝYy9A�Έ����`s"�=%����}"KD0�QGx�5��p��?㝷U��<d2�0�b,��Ƣ+�cOu1[����gT�Ug��X�Իt�3:�,	F/�x1��a�-�Ny��W�ED��զH��		�w���H� I(|�w ���@C��nE��{߶�P�=W|�[=���y#to�0����k�g��'į�y�x�پrޡ�l^�~���5y�$,�ug�G��1�K�>�*�q==E�Vck�eK�Q����.O���3o7����ؐ��v��˰�?���M��j� r�[�~�`����j���؉3%&�9���<���~|Ґ��
�o���s@�#aJr?�H1��h�]敜��0���8�]fB�.�Nt��/\�BS�;��(�Fb% s�r&�~a�=ZK�;�/��(��	!�Ḻ����/�J\0>s�V�~��m���MQQG�����o}�த��1�~]��á.�1�@
#0�=h�[�:)���;����i�N8i:2��sK�b��b�8�* 7�y�7����X_�N^�0�Y�ih���H� 7��(r����|���4�B-�w��4 F�7�3��%w9����
��q�?�dD;�x7���z�Y<B���ZT��\��],�>$mJ��Ó�W�%�r#S;T��j�3����+��"9�Oj<��A��փ�=���u���o��-�"6"X^Ʃ���@4����}�\���O+me�X�k�
�J�QM�>}�����d �X/F�V��f�z��ȶ&baz~2���z{�&�*�]�;N�g�؇ѻ���L�(�<ۑ2c�@&�J�\`i�gr�L���H.�����_��x1J����,@��^~���h��[��՝�28u����Nv�*ս�-W���!+������� 耔���������Ş!��5-4s֗�:�����El�Ls9�B���[_Ԧ�=q[�� �`��FƙOy��-A��YVoa�IvR�Qc���/ى�n��٧���|�����R�,�3H��j�����+Kv@������v+�'��@���kqf�B����r�#j��l#h1��j����(�
�:+1��b;R�yk;R������Ŧ��%acN�Nrӽ�>���_�8��)s	���]��C�$ژ�_Gd�b�?��l;���V��em�έ�~�d��R�!�V���
6�aqHU���n�/K~R�[.(�,� !Q^j݅g.�p:�oɨgQ�
��2;��>pk��/�0�����r��MJ��}i\�Wx?�v����[�}ő
7�����p����t������f�mx�s溏�8��Ja�y�Ol�;���sB�2�_w=n��_[e�����E�uV�q�����d�����vџ�d`�h�m�>��+/�e��9I��-;?x�� ��YU�)3buc��ֹ\!�ӑ���ۭEc-_n��a�E���¡�&J�b�dBb��%l[��rٹn�\/�M� �y*N�J���¬��}$�s𣻞HHl��Z_���0>_U�p$K�	���6�?ԝ�� �xv|���vޞT�/Ow���2(:ȿ�z�x^���a}I�E^�S'^��.��ds�!A�NvY3�g�
��@'yGr����ќ0t��M�܇d�
̮���ʊ'&Q�Y@ ���nmH�~l��]7��'��N;�Z9�K�n=�he8��$�W���-�8NgP�ʚ��;MԂ�o�����|�t��`����=7�a��(Dg�Ck���*����B��a�~Ϫ�0M�p�b���r�`htl�K�.ٷ�h��\�(D�����#��V�5���mb���~1��<�rE�n�44!�*Yt��?	[.���Q:�5�&����Etwdw������w�O������l-�,ET���uU�5��ggKH�3�O����vP���|r3A4�pX��ͯ��Q�U�P�H�"�p�>����_��JgW�w�&���j?��x�D�/)���,�.M1vFJ�^#�="n`���:IL��bA��p3��L����Aq���~D�sE_%�d�;���(ð�J����4��SR���~:��1\bX�Q�5lc5^����,�#��#�k���W-Y+�-��m�.��Ĭk�Rjj��2_4�|���n�	%f.��7����4�㤵L�L��ϝK3_R�$l���=q0�؀��_�ě�׫�����d��C���ݐ���X1s�_�E1�ѧ����5U� �Q���B��؆J�e2�;��a����ۯZ�arg� ˘':ث+��2l���*�	��@�IT=���xB�&��K.Ҿ|���ֺ(�ԫ$Q���i�]J=d�6%�/j���f�~X��Լ�T�y�N﯎Rz��fsန5�}pT�{Y]?����N�Y� �;%�Y(��d��LC�D��1�ުG�^�����mA�
�ǚEė�GWKaxae�M�Y<�	"�giW.�����JۥJ�"p�g鏥�*��N��Nq��ܨ�-:�5VJ"3��r�*eX��<_�]��o����0���oU<������U��
C2������G�T[V��.���G�Fh��>Y��1�K���G3����(�~��-$6��:F�+�f۰(�� �á��-�@U�|���.]7L:N��Ǟ[�	s�\�BB�΋���O�)��3ȯm�����v��)#�3j�$L��e��e��Bs�F��]�`��ɳ���q~�-��a�S"{+_���)nʗXpܭ����zl5b��z�6�0H���I�[E��v�`�����Dr�����˧f?���Z�C����i�s4�
|'�Y	��SU@³�_�l�����/�F�)���K�ش�u/�[ЀT$��0hT��fg�Q���MO��F���?��!�∼��:���zȋ۹>A\�k� +�~�2I�3�+q��yo�.;�t��gb�u��(Ќ-)Z��L��1Yq�v�2C� ���>��ѩ4h"{*	3`�X����vIJHM���� #&q��h�Ua��Ŷ���؎{�$�E�o#Z	�^��w\���0ȕ[��<o ��ظ׸�dr�L�|7�D����t�P�3�Sjx�Z����c�z�01J��1��.j\�5p�@D�auATd���D�9rw�W��+�ُ��}��(���{r������Y�������\�%h���\u���hǕ�H�֯�8�%���T�O�����w����0�⣥h���r�6��������\8Dj�2�֪0DP(h�8�G`(����S++�����
z�6�J�[]2I8�e`�3��9�k�Y��EV�H�����^.}���d̐*�ÂI�%7W���kB���=���g�bf�����-N��O�8�7�#y�c ^j��k��55Lf�Y�D1�5�a��K���ɕ������%4���lb]�[gsT8I�u֭�p�e�b�^��-�]er��$�M�VG��q\�l��{�Ov�$�$j�!�+gK�z���3e+ǽ	aI؃uoV�f�_��0ė�B�@���y\�aMh�����x�)|8���;� ���Y�g�����.�I��R�T��;�e�0�[t�����0Լ&B�����e��[t�Yl{ڱ$	A���W�v�;Rn>���3��!W�$Q�)��d����D�k�DV���%����l|�!�\�Э/i�^A��X8�5$��J!hS=��3�������hɭs�xk���\�b�E��d*[<� AWo�dbֱ�s��<rŴ��'F�;^9q+��o�}�_�>��.	���?<iXܢ����ί��cID�a_��]�[����{{��VʈY)�);���@�9�,�n�� 3m,1�XȹYw8���I�x��7J����8��N"5jcꆘzS��P�7`���D_+�QW���8{�w��o�k>�#�Iiy�q��xb0�^��]��{��7B� Ηt��߶hY8r��0����y����1gOBs�0Z�6�����!	��ξ�t�n=�K�ږ��l�������Ff�H�/.���jh�[HUD4������W����Œ�I v�rj����~�ǅ"hY�tϦ�!J�ۈ4Dyg>Z�RI��LĦ=�U2_�����&�B����/��z����#9�Ɲ��7i6��v��ª;|���Y�ۜ�K�j�n�.h�`��pؕ#x����l<E�8�����\�O@��<4%-]8������5on%����rΫT*��)������ۧ���g��a>��{e@�M��kx�^"ж��oW`R%Qf��%�E�=~(��Gߞ��J����d
�d%y�O�.֏��&d4�!�'�cB���l��`l4�KU[�o�0,(�5JR�zkA�s�`��>�`Ɔ{��(�8sP�Q���;�9�u��]"H!<�9��������ZӒ��8�ƥ�ڞ�����"��Z�/7�c��U��E�Lw��Z�{��X�a(�},�l)��l#��%��Vi%~�E�e���~}���~���_5$���l<Lui8I͆-����JP�
���zͤn�����R�{����ۯ)=*8	 ���o=k�������*0#���q-/��g���y�;ʟ���h/�����Z,-�}o����c �ëy��IX�1� o���h2�mߢ��М�L4�/1���菻}������;�떸j��f�LMZ�S��񟉙FqΫ��걔��y�`�&݄3sX;guL�+����Z����G�sy��򴾂��%9~۪Ǵ{5�_��z�z�v�I�!Q�����Q���4�u][�i�Y��>��0�J#  /ǵS�<`Q����Zű��h���Ka:G��]��!z+ 6._1N_;؅OEs��cт����5��t��Ǥ�&A0
���Z�4/� R���eX79��y8���2wm�}���� �F�1(��:R��h�p�Rǣ���B	�'u:t}��Y��5r�1u���"v�s�� �l¡���
{'R��$Q�
�pdӭdF�ą!�/Qwt�{����!4�[f���i1��8|{��>,֘e8F�\�8�c"����'���,�lR�1Td����Y�a�����U�3И��ot�����o��A�n��������5C`����y�[��?�	E��;�Quh�v��ef=a�Ԣ���jS�	:Rӷ2��gN(�:~�d�k�z}#�8���ǯ��ݫa��S�/�Zq�'� {�Y�F�/�:�Oy����f*�����(H{�i�=0�߲\��i�h�UD��	�N��aH� �Gǭ��=Y�
��d�<���w����Ձ�[�Bผ��o����7�b����i/B�	��˙Nk��w�2wA�S+�Ŕ��vpk2���	��������a�e,[�c	Ҩ�!�&�;�ͣp�5��c���
z	"9y��Sq�*��[��-��%	O �](
���VE﫺9mv�]O�j�v ��e��~�_F��z�?'#��Y?_��:<k�i����~��0:q��|���t���`�?�@f� f&Aʖ��oII�Oh����»
���R�g-v�Zņ�ih:D�|�Y���]�g�;����X��&Iһq��S��t��zoU�\s��ZNrd'�;�O�N���LA-=Ÿ���q���+�]	\B�.��O��&s� ܰK ������݈֤�M���N&���d�4�34r���;c%�TLI)}�g2�Z����� W��|
7�`<�g!%)��AV�L��)����m�ܬ�7"�/��<��W� �1��.b [z���y�(;^BG�@�Y�l&T��4�y�hH�0�0�1�\.�NyS�N?�Y�;���Ԥ�<�b p0-⦙'`im�@!W(�dpF${�S�U|���F�Օ^q���^.�f�RI�6S��w�0ѻ�+�6فŏ="�ڔ9�3�E��=FC:�L�_2��Ma����I"�Ʀ�p�-�ȉM���u#���Ȩ�C>�����Ş,�@��S� ��H)�ҏ��D~�O+���,?�l�O��.�$�x[�$#@�%?�ǵ�c�\|ĹD)���V�Y\�8�#��`�ۈk��	�7ښ����h7ǃ~ġ�RIU���'�ߚt_�nR��N�d�r�����s���J,�	�	��Vӟ&jT�Þ@�wc}�=�J��0$�r��f�gϦ@�_Y����E��rE,���6��?'�뭪��>&�K�������p���[��@������䞎���{�Nv6X��:�7	ߕ���U�Z>H�����̕��̛5���ɼ��Cp/P��o���hs���X;���Τ��1ǰT�D���
�r/u��-����TԑMpM߈B��9 ���mc[S�k�Zdc/�u���
DS�i��7�����Jq=�����YE����B�d����HMU?c�h !��M��-qq�t�;���L����1!*%�-v-�̛E^��P�E�U��m�&�5D�WT.ƞ��/�J:�ϗ���lC_m��q�֯�d^2�����rYZ����*��	4��`9IB��)��H>��}X%\]�rۂ*�lk�z�{f6�D��A7D� ���ޘ���l3�dU������.ͷ�~��>b����A]b(Z5|cb��H3�?��}s��0A��UX�7�W~�S�s¯\`�ǘ���>_���;�*O�vp�j�B��`LZ�%:ɀVܛmaj�j&�������wuGI�1�Z.rmUH����|�`�Lx���g�u�4����3�z�5��~m;���3��Y19I:[п5<XL�a�*!�
�ʛ#�Z�ġQZ�i%�+�!�Q��xD����C�?(�+;��bi�K���Lʊ�-{Z �;��ΟNhr�DaI��z���9�8=.Wr�&���8J@X% ���|m*C�^��ڔ@��:�:,��2a�$�؃���j.�T���+nZ�Af���-�J+*d~�F������i��E�80�����X{:�cr�Y�uқ��,�ƌ�0�<:l=3���K�U;��7�&@9M�䜹 �7�(�*����Q�
�7�/h��:�i�E!ǁq��*�e=t���z��Q5|��/15kNX磪��چ!w��ĩ�s��,<J3���È�MZ���?N#�l���g�h��i�@*���|����F�q
���Q��ܿ�:u�E͟�S+
*S�psKw��VJ1,�����"Y��ڼ�K\=����Q�L��k�x9�t�3y<�r�$;s�ğ=������a@z�Tv�eV��D���;�3��.����c�c����t���v_��u�2zM����p5IM{��]��6��0V-�<�xO�OI�N�/
b��QZ�k
'��]�oV-�Ogr�_z��0��+�M9���Δ:�_��ɜw�V���z��[�l����B����g�帑�<�3~ [���SH���:��4�FV��g`l�l�AZBE.	\�%���5��wc�\bgO��U�N������p9X�{�ho`�ApD�9-Q	�M�GDx�
��ĸ���$q*S�����Z� hoK�!������^� !	b)�M�ƣѬ���iZXC)tn��`������V�[�A;�����Ru��	�vի���18�b���$a�4��������Zv�DSz�a�s�Fd�'��8�A2U���f������NH�E*�u6�E����IS���YK�����ͺ���uOh��`if
^��i�Ȕ�~G�f(�(�z���4Nk���5��-���҈^IA��x4�6Q��|cQ��@h��Z�B�+&TS�8��b�Z�A'�n���}�H_����di���o}W�����R�>3�M�l���1s�<F��;�U����^M:|�ZY�H�1Z���p�~��<��4��Y���ɠhP�ʼ'SM�qP�ȧ��P��|PF��[}��p�#^����3�	�`ǰ��uC��뉥��6���]W�roz�3����<6)*^4�\��!�MⱮE�'�O#�����v��3��f�zˤ����ǧ0�zW��:�δ�!�d`��t�־�e׬<��֌�n�%?k��12#Kd ��,��o�����
8^�N$�kEN�[��S��U�*�]\f3����H��'�]X}8����7im+]�=߶d�������v�@�>9Yg-�s�dɵ�kϚ�E��pNy�A!��8���4=1��l��S�8˓��Z�I�н��\��;����6�0�ۃ�aP_���JY%M*����>�T63��Ai9�w���N�Oc�I���t�+)�]l<x�'�}�U\N���.C�788�Γ��߹n��O�X.�7V��x`*H�M�E딁��(ԧj�R���	}�����;������%���;�p.o�$�5�* �:��H����;��H5I�L'dUX�^��`h�,a&��݅)��iPw���X��%h��c��ߢ`"��x�.��B<nw��eU�'�e�.|U	���6SB������E��(s�T�$�MJ��)��^6ŀT��k/�K"�nl�;{%�;��|��7cI�R��sb˂�9}@-<G�jt39��pL'S��@�0�r1k|�N�X������\(sX>C�1�����E���zP�²��i�Bn�D�m��AI�N\�� �	%�۶DUO�
��{]��3�9?5oa|.	��������b	ƍ��=��f�Le����%}a�U�{���di`�N���T�l�I�1�%GZ��.`h~婈����|�ȨR��p+�X�\RA�1[>�3��\_$�E:5M}Cd���!��@��J�黡�1e�rTx(qQ�z�W/\�X��&A�C��-���N�A(&~1�0����v���
mr�\�.���TK���:Q�U��Rz�uWj�ި&~��,qu����oТ��X�`�15����;�٧4�9l���;�,�'q��r��#9�����w��ʠ�EE���\��X|��q��,N4Z�.�N��?��:P�h�y�0�D[���cƠ��:wP��nQw��k�O��}<���4?���М\�ۭ�/E=��_�vY���VY���\�����::�)ns��LC�
�?k<��?�U���yG'W��`f��)R����l]+1�+i�r�Hn9��k6�"��{�J$�#,��kX�����H�pyq�<2���G��$-_��y��&&#��E�g!)R="g���e<g��d��Kx�\Ŕ�7P�(�	|}B�L�ɒ=�y����L���_@�M?>ַXhsC'�����,�
�]<��-������ώ��n�$#C��t�R��<�x�
=='�o��}�N�CϦ?h#���>��-,����K��N�� z�� h1k���z��I��\a}(xԸ�g���*U�&��?��O��?�?`]a��S.���׹�	���{�vَ��fz�mj�Y3�j�^�� ME�p��a��"�yr�d:i��&D����:ti���ɩ��v<ʃ�l�Ӊ��&z���X�G�	��[��h΃i�M4-+�]_`��5A���"~!����3�+��E��\�L!1�g���t�"Ha@/��~j�I�q�e�i4��Yp@}߃��r?:�:A(�����Dɦ�	0a*O�-�-��]%+��
�Y��a�~�kd3�����2K&~ų� u��~�l����'�Xa�A���fQ�UP���j2�1�/(��yG�]��^hF)��	H�V��s�}��y,�9�6//�5��y� ������y��~�F.�)նE�;Fw�0���繧�/A�#<.�i�T)��T�|k�/ޠhgq�B&��E�M�{qy}��ܑ2���z$P�?��K��-��_�64y�ø�*%fy��u�K���􀷜�1.TV���8z�@��%�z���.(I��0�+s)�W�j��'1Ң3���W@)�˱����Y��/�`s�&4��Qjg���Tj�OS��]�ċ�xx$��� �y�8����aB�Ԓ7=y��	��R�͢����>fJ��x���&Ľ������N�Ǒ�Ƒ�����\Q��F�!�IWC�ZrџMJB���fm�d�1��5&��d���+m.��q12��%�-C�t8�}I�W�W�V�h�33���N���g^T�8.I85��?w�?O� A^J��0J_������@�m���#���Ux�E���b��L$�����Ŋ?dԆ^SH�P4�F
�:5n�L�'�?�[�&o+������t�R@���ET�eƀ��\$�Z!19���p,�U�KW?�[A��u��[M����U��=A�l|�;B�����S�i��9L�k�D�ޣJ����/��cg��<
���ҳ,o�_�Dy�����KaU��� ��1!��k��F�n���4����ш�&�fEx͡�V"���Dw0|+ZN���бHX'�ye�m>��5�XQ�L�M������k���v��P�k[4���11�N:���8�=-�u���:X�TQ�ryw���10a�v���Ra�lP����!Q�7 ���<���\\����y �{��͞:h+a���<���\� �v�,���6� ������K������hlة���N9@�2���R�jz��ۯ�deDS%6<R%r˒`��T���Q�6�^hP���L�7���eGsH�E��B
�
0�m���}Ϝ當��\[��g���
#�޾·VnT�.��,Q0b6�O8�✊�Nh\?�]�q�b�9�%i�{�F�ʅ�y��Vu����ɼh]ί:6��9�NVFc�2�������O]E��r(SU+�ݫ���CwšBu֨BR�3�K��#����� ���H�wQ��^�mf?�|(p��}�:�'�\I���n��{��:�j�ᄰ���_U-|^"8w�T���H��0�V���ب�0 9���B�Yl�m�?��'�OQ&�������D�<�hb݋��~w4��NX�Q����1�UC��d�E0�����[������o�a��U�$��(�ŎA"S�u�e�>���?�A��eS������7�K�����(�RBC���A�������Z�^ȑ++&�P*F�TL+�^�v�Я�-?�$t��0�j�)Jk�%.,\�(@�3������+-ы�$]��@�����ʰz�k�n������Ɔy6R�������!e�"�B����?��,�T��ū�~� u�f�o�w��f�י�yS��8l���1�!v�P�ۧ֟(x3�4�'S��f8|o���nLl��RuP���jf���+�W�z��f�>+:f(H8�� �*���9,3AЧ��I8I����	@�.nY"F�"��ډN�[���Rf�'��2[��
Ȍy��K���d
$F�/,�<���I�N�?�]0j��\����?��(����>�5�kf���$�Ɠ+���]���L}�9�%3����ٛ`�By'ۓՕx) �,���Y�}d�7 !ù��=mE��	��	N8���:�!�Vw�]!���/��M?��6C�	rN��������%&��	.;��a�+��f�N@q�,���ѻ��qS@��p��sނ��^����rK���'"[R!p�ę��u�h�{�?ο�H?]�ދ���
�݁�P�v���_O]��CҀ%��c 5wMp�b;,�WB�����ZM�ݚ�坬��if�?Q����T�z�ɄD@rn��9���CtbR�"�zp ,�6�0���/�7�+\I�?�l�gk��hd�P�F^�����^ksJ�:_�
Й�TX�bt���\Z��j�2���oo�C�!=u\(<�x�0�z�~1�:V�����1���s���R�3�ܑQ�`ћ5K�5�4ׅ�Q��������&��{�s���'�bJ8{]���u, n��kՊ}�|l9�C��1��5\W!��
����Ll��ŔmD#w>��Q��7^����a|AԦ^��a�|rPL����E���Q�E�/�^F��贽}D�(���gzb.&£�s�`w�w�9�̓���Lo�����LF*�#�&��������$�a"xe�,$鑤�31�^�q�����i�gs����G\�i��.<l��#���+/(6��.A�����ۜן�]����d6����V��lן|����/67%�t@=)�Ʊ�R6��g�Zt7��{s�Q�1�V��{�{���*�O�y˾��d�o	I�
�n�(�n���Cfy1�x��}�(��j�,��;G�\YL�Ӑ�
6�����R��FS1�mP(�����0�>�b�6�g�3\��N�� ����!hm#o�mѺ�>���u̹!]��R�Y8v
����˽��+�P��l�)9!�[C�y�Ɯ�� h��������/BJe��9�F��� G�{�F�x�9�'
(ִ�����B����X���/dz��dZ�.UŁS��t�R�"���>��&��Q>F��vθ%�vD����<B�VP,_���-��^cL�Jw�I��͓CN�"�W����>���m�-
����h��^��ƃk��r��3y���9�Q���É;�b�h���������1���[�jTG�|�vt���=
�=*��v��1��)<�p��Jxl\���t�*w�l�|������G�[g87�Dnk�I����ZFa3�u�,r9���֛'�:j�w ���h�����Z2=��6uQ � ����Y�h�(���Mxc꠷��<��������F�`)��Q$��w�W���%�ξ�&���&��8��(ۨ!�$s�i	ȫ�JIG�2���YBo5�}٧(����^�2���O��<��2���m�����\g���j���� ?��n�,Cbo�8㣐���ށ)���[	�g����+�~),�Тk��
�q9��)��	�tð'�"�C]+�z8�c�wBL{Up��i��:H��jyd��&�K��H,W�j���H�ܯ#�+�ʐ���`�x&�Q03�����ճ��c�ڪ��-U��_��	�vI��	�����Iz<=f�C�8�|�s������py�GPcMmp�T�֭l���!�����<ܚ	:�0I����2g3⭲��\�	"�����bpZ����p$�,�s�psR�E�4�@a��L��/�\"7Ӆ����Tj��.6KRƨ ���:�vURpX�o��d�B���UUB� ɵoI��w$��'�
Qs��I����?��A���8FS:�[眅���3�Ɛ�ב����K.�:y	(���M�ο����m:�/e]QNΥTQ�ۂ�+ux��6'ss6x@5��.�Z�5��;�u���,p}&d���"0�VnN�B߬���ԕJ��a~8ǽi`$�[� J��J��0��f:�A�Ye�E�S���"�Р��z��#�����S�9:�u���M(�?"A�P��ҟp�8���jBEv1�����S W( ��fj#��?�cޠ<�C@A�>V?c븤��è�;�я8��;#bR�9 d��,9��"�tK�7.�4��	�{oo����9��v�p���K廯��I^j���Q6>�Ǜ\k�o�\��wPB斤-��i���e��gL���5iH5��Xz@��u�t6g`B1��a�<�����	�*e�~U�A��\x����,:�� V!c� {������+2Q�gd/�,p���6Q�,�7M`����|q��G����J��?���ڟ5�������?<iJ�z�^X*���sf]� �c��,�q'.O��`@���:rB�Ù�yr��.z��P��\�V��\��[��7��x��*q��Af:N��ߝЂ3k}��b(R�&�Gs�'bS�o]B^7'�3g��,Y+��}!�%�T���Z��,���0�}�X��~@qV���rML����L�C賈���-`S��"eiEߨ�C����ҍV�E��k��C�M-?R��%��.p=<�q������\d�����������d�^���-{#�T��l��� � �&����4WL�F��y�Byl��$A�產͉�jJ�{�8�A��(D���ZF<]B����WtZ�5�Ga֞�fV٩Ttg7�m	�c�k���'!ש��s�c�Vk$D�a�P=�
�=]��b �&)b�A[�_�� ������{/��b�X�[@���>%N7+��yu�>}��n߆LQ�H�E
*zz��eΧ���bU��h�o����9 �]�}��UZ���T䯅�!a���?���A@��,�+㡘i��[z>Ecb;�ĩЅ>)A �\-�Q��Zh���N�-B��~[��G��W���xq'E�n%u�%D��0�N�oUD
��'��Xl�w�L��D���3r�qe���C�#��V$�	��kY�<���@?����ZFAa�#)��2�h����� ��p3;]ʌ�ꎃ��uR1g�\���1	6h߯L��}G+L��4�i�s�(:�tZ�3P>kR͠U�z�@Z&T�	
1���VhP{e�͊���n�tWʱ���4ρy��%wj>	8f����,��H?��M����q$�K"����C�MwOU�GkDu��/L4m�;�ʛ�UC�����Js~��(b��RRS
��w[�~M��#d�NC�E�͇�&�a���,����)aE-Q<{�ܕ���-�!2��NeR	�xm�'u�&�3��4�9�Q�}J��������󑫣�-@�F�v�E/ƹe����:��A�U��U���KH�g�0�xТ�Z���'l��n�gӫx2�T��d�U�S�
;�#8�I�$�^��Ƚ]a�;�f?h=�2���V0`�����v�K\�q<�D/��H���~ش�#�U�������x�G!����ʬLO��xi����ǫk�<{�����Y--R�r� ��,b�]h�|"]Mn��&!7嵴*��*���Sa�G�x�;�kW�T�`.���tѫK�\�����|t��N70e����"�����5�
��8���%v�E�y��>���M��/֗���Yb��.��I×��;[q�^Yt�t{N�`��q�.P<l~㛤dhkpxHFH������J)�(*i/z�x"ǰ���?�	�֥ �4�_�3I��q���=��o�
�� s��А�iJ3㍣��1^=�q��OW�SL��F���I�o�R�;��� �W�k�@�>N5A<�Ǐ�DP��6���vl/:��L斧=#~b������׮JT�9Ӭ��V&�ʧk�uy�aX�T�e�>�n�zW�~��dmѠ �rA���Sy��vj/�U�S���8"i	ūA9���`�g']��.x�v�����w*��52'���Sq��-���Yϊ
p��V��[��V��b��T�|x~aWT�v3`� ��j���:}��8ֿ���N�9�+���ɡϏ֬��!�������w��5۵ �\�ۊ}�v���DrR���b�r<O�J��1�	�OmtR ��m����(�L��d}�'������9E�l���g�k2�w���!B{y(+G�q���j�5vuK�!S���@��:�%�G*"B��ԫ/Ζ�G�� c␃�Ǳ#¸{��ٲ�y@4+Ȗ} F?��YN}_7���B֊sx��aF��?W,+8���d��hk1 з�qyL���ܫ��md�ֽk4�5]MQ㏱�X#�kF���H����x����Z#r�]$��H�f������:���?V����^���U��~U�j������I�/ED��SB�U#�&���Ir��";�O��Ĕ`z`�p ������+����7�/{�aN�6����EV]1�3�<�زq�
�h\`����jԒ�ˀ����'�J(d�d:�(�hH�3o� �K%�ӗ���2i���'�I	�C�xc"B�����lڌ������Ll_�^j�w�1X<�{ӓj�����}��~�A@�Aho�k��:��V�?5�����S/#!
s�代4"�y��1�b�3ZɮA����fj�i�[?�JUT@��TC#A��j�_��c�*�(H�zĒ��R��&-��l�|��fs/��1O/	��G��ue�\1�W�^��[���:�@%l���ܠ��`�r�c1��&l-�]��?\�5+�ٔ}�d��?�lgz(�F����Z�<ӦI�4�]�4����+j?o�(4dnu�$j<2{ޮrT��  ^G��#k����g�)mRRu��|_QN�B�H�c|n��~ͦy��~/�_=���p���a�ٿ�NfX��4җ�dxB��2�>���A���;0L�.5�s3f��ĥ��Ie�˫<}��mQ\��{����T3� 6���d�l�ae"�ei3�}��൉ڞ���E3Ch��g&#;�����1\� ��a cd=\���+���rI*q�F*3�ѐ(���WY��?�)�T��ɥ�<!���hq����f�Ҁ�ґ�X��oo��/5�.��F�X���dA�}�k�.{Ho�d��i�k�Y6��}�uF��3�El�ͨ����$���� ���"���~h�N�q��D�9���gEp\��#����l)�Wi��/�rC�9�ԭ[�*�4>�ȗ�p��M���q!�?�Iky8��N�N	Y��X���Y��$�9egǂ��a��`�.P�-(0`)�=ccX ���յt���c��ưL�,;[�*O��a���wR����l$�g���#���0Iɼz�Z��f�2a��EM_�D�����l-�]mы��k�&�̎Qy��v��9%Y%a�B�F�+f�d�lևZw����a�'0��O�\�
s��X�\���\�β� ��Xe��)P�~��Cݱr}9���iM�N�b�D8�Sڗ+��!I�e��P��I�\/�kf_��LZ47��f�_�ƃ���྘W���[^{;l�c�B��P�{;2+�c-ul� L���pa��\�!��v  ��|
=]��G��/x��t�1��&(�֔��u�;�$T\�a������α�ū;���qr����ڢ<s������'����	������N�]�J^4G�3U:��*�VԊ@\���]�~��р^��eG�K���O�F�ZԺ{*g��^<�Hܲ���T�ֻ�Y�w�ʥl��#�	�+���85�ͼ��q�?�e2^�IV�0�_O��[�&qXV�� ���(�F��;�ULm�E㞋m"�-XH�61�ص��,u�]�Q�j�jb�Q/1�ב�����s&��u�A"ƅc�@���u�6���}Z��^�Q��M�<��QΌnh֮���2q���&�Z��D�ʀ<��٪�S$W�"��M�y�X�]����,���: V������i�<� ���B��B�Y���?�