��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o`���d��]�v�1d	���u�C�[?�ϗ 3��kNm��5�/,��JH�Rw��$e NMF�K��w�h�0H�ai����I��@	Kx�"�l)s�ŉkKz׷�
��[c��������l��u�_��Ss��"�7�����K�Y��F��-Wi�ؚ`4���P�P����ԻW�2�V�gO�z�*qn3��|ע�Z�e�g�������!��4ωG�7{},T�J���5��Ƒ�~���80�F�sH���U+i����:U��7X�R�lR�O�T�p��d�v�������@�y���>r���N�U��h�N�e&ٚ�j�����e����-y�{{���m|^��}N)���-�u	��F�_Nu��F��ʊ���Ns>z��=��)m�"v���a�@ZP�I��UP:r��i�_+�L���z:�.��rx��\��*�c���!5�{s�_8���{~,TL 3��Y
$����1����(�M�@�4���+��[��#r�.�v�&ZMI�U �x��Z���hX��$���ۂ#�_*��~�8�ѿ�'*�Pv�94��M��3�a�|���L[b�	cA|���.����^�r]C`�X����XAH�>mI7�H籺_��s��z|��㶰�e�*�6i�]�'�}�h��e�=���Ыk�8��A�99����w;�Q���y�I8K�J�Jf��Q��P���,�I)�<�c�غ��듪s5��ZR������*H$��L6�^��]WW)�7�i��>�PN{��=�am�Ӏ@?:�`�v	m3.ˤҪ).�aF�c��f��1J�B"J�u�Y��Z���N��ö&�W�Rd[R_ErjL�a�������b��>d{轓��}�_s�*ݽ��]��e�6��uL��>3G����e�%�ԮZ]��5��7�x�i�C����5:J�����.�E�
���>�L�,����
����A_�K���mw�+|���2�y@���<�����v9�®�9���:�:)��;�1��4La�����u��"d�YF�eR�jE�j4.^P�`8�p8����%ǂ�gTĕ�y`Dh;��[#_!Z�X9��Y�r}�����P��;�V�^�P�o<M��}"��h,�M�^N�`Þ3�F)G�2������6H����Ŋ�C�M}�q��Ia�2���D�)���U�w�U(*�H!d��9ț��#�OC��Eq�SrCk��'}��X{P!��\�b������[ф����^���8..�&��y�g6U�ḧ@_��L`^"zP#�t���)܏��Z��R�t���3|Qɫ�x�amf�f��Ns�[��R�}i�0�{馛 4�o%�[x��F����R���N��롘߲�`<x"2��A���M"�u�ˉ2��Г�oo�|(����ި���:���`	��Y�.��].���s��9���2���
Uu�b\W���T6�"ק���7[W�_�E���ȍ�;��09�ޗ<�4�3���S�ϱ�8]��ֿxr<e���`m-7�L�彩RG(|�M0���gDjw~�ES��@�&��[���)}`ǥ��}/�a�AM�mq3@U^O��("��j�\>�Ԁ�&���$s�chܱK���jbj57�:����qC�p�Σ\3�l:AD���u ���m�4  ((#�RYI���;��mu����JgF�lmO^�X�I���mĨ����@ՙ5{���OQ�`��"��2�ɢ����+�l)D�2��m[6|˖ܷ31�\3���$��p�����-�^}��9��=��hN����+YlҭY%8�`U}(��1{u����͂ ��9������X��(F�1d��4�8���r��+VȒ�_:��G��_�{�:��"��T�?M�W(�h�נ̜�)���Ʌ�/ �},�l���:	��(#��FB�K�p�n���Ζ
����(>L��P�X h	�QX��pE�;쾏(��V(O3Y8+�c��@<`!vy��}�0�Qs�Z��Ih*9�+}��ϣVe�-��Ս�zm^4�17�ܞ8p �ᄇ�u�d�\8$�<={����՟� �n�;��/��J��S���T������ {u�����g'�s���&Uq�ǹ�8�2�����Җ�g7��Z���(V��T��^(�x��^���pq��L����ϭ��H\
g�c̰_�%��0�uH���/�}bG�6�7�2�-W S�o�w۱��z)h=8� ݨ-*���� ��s@��5�ܫ���ձ0|�7��U���/ma�r�A�̔�
�_�cBՋb�@�vhO���.B�/qb<�;�a��=���D1׺l&��Fj�2���:�ŜL�_v�^�9�5*�X�AD����H��27�!{QtΙ�ULR��mF��ݽ�rG2�:�R�/�"��G�������*3�"��Vi�|\	�6����We�Z�8�c�& q�*5t�����.�jj� �=�3w[5�L�z�H>.-Ă�o%n[���dJ3�Ç��w�O����m2��3q����]�l�Xw���u$����vǪ}ua�#�'s�r��k5��y������F��&X�F�M'��½]乞rGf�Å�A�E�z���k�Tb���+��Jk��kM=�1�����ME���u�=�%�W�$QEʎ�[�'/Cޙ��A��B�t�d�_�u�$�A���У��� ��GDq���RT6:�묫��}�'��P41XՖܺ]m�t��u�T�&cM
 = �Ag:��f��Q�&5.3@�)0��f�T3 o-֍��ۧ��a+��y�?e0���Oa\���d�t5�]& X=�s�h,:2����͜���ДE��P�b�Y���\z��ocT��@�pd��W��@a�^騮ţ��O@�q��_70�����6<D�t���ޑ�۴��ᇇGe���>c<���I5��������R$·�
Gr8�K�<�0��6m�u��{�:QZ��%�P��E� v��@�*{f%-� �x�=$�#������� @�pܪ�-<��H�7>�	桾�1�EP	��Đ��dVB�oNvHGO{����1N�X�@��"ٵ�����`��w�p4�LpEW޳ӹ���6�������i�*��k!S[-�(�ƃ9_���%�i����|؞�/�n��:��m�>�!U�u�5�mA��yq<����{+m8	�@,��T2[������ԗ%�R�y`��;'k�:�X��TVS}i�"��!�!|��Gi���ʶ%	�����qp���h�F�E�
̌������%����9$k���+%�E0Sӟ	�5�)�.�t������$D�	�����f1wrh�Bu-�3%�C+��+�W�����}�aA-��5�cΓF�y�E�bZm���n B�l¥l�W��s���� luth�3�I�K(�=��ˏh������[�2����<��'�n��/��m:�:`ǼY�Qմ�����nf���6�`@Zk�ESV��9pS]�:���� Ζ���Z��R���@T ��Lv�+���|E�3��&Rwvu#�:ϙ���]n�rW�����>'�al+ſ�h MI��f���b�@�~P�7�p*R`�I󂲹9�S�g�C�e�����\#�\�����
�ri]Y|�����u�_�^Y���x�g���9�k^hр�����sB\��:�<��?���u�e��*�g�r6�	i�ۄ�Tɝ��_$Au���[G��,�AZ���K�n�ςIUyo���`74���^j��[��JvF�Q�/}e��*��pM�x�{��g�0	 �S�m�?�*ĺ<�����e�J�r��Ț�����7und��RT����Vœ|]A �1L�9��g+�w�Ϻc��K����L
��]�z�üK����H+k"�iAg

k�.���  ^��{/�����s7���<�A?:׳�X�|��N�3��,��˓�~S��<Gץ��+�p�H-1m
#3�B��I��:@-L�NXC�������D�t�
��kzWn;y�)��;�>�ZX<Vge���77�Ead��I��+`�G���eq���8W�B2�M��<(����'EŀvO{#�G,��m�1D�"�X�
�ކ$�3��p�f�3���
�XO$�J>&�Y�U �r.f���p/*l�/�k�Ⱥ~������B�c�﷿��Ȋ|�Rds�����L�^�\��"P���o^�l���R��A��:�}��C���9S�0<5z�H*
Ms��=
����we�[����6<9LOR����x��h-��=PΧ0&�?ՠjeÆ=]�p݊۳�0{��aH �Ӂ�>�zK���n�N�<02NS�'����&��T�W��<��T��mm;�Ks��'�!�9#S����
g��}h�w9N���+�L�QחD��i�^��{�m�fu?%��9�W���g@��~�h��I,�"�\+	o��3b1X��!	{�Q��\c�4`WaYY��t��O��*�U
`[�%��7 �@�a�V��C�א�sm-�V5+owl/�LÚ�gI��1���o]������͕1G��sS��x�[��p�V��K"c�a�㣛m�=eoI4��i�}� Jw����%=
�M��O��/4 �}�P�ᝫ���iq���a��c��iJ�t88M�������z�`�+ߠ���=� �r!��e�Q����*��\\f����{��L�"8^��\���}��3�U"Rڝ���0%�ۈ,�V��@2Y�d�A���9�:ǩÌ��ʒ�ߑ{���e�|6�N�x�%Y��裢�y��2-,����`k��C��(�9~É�a�0�j��[����B0rw�� ��f������E�,��p�8�o	ſ�nJ��f��Ga���h��L���S����1e!\�BE�&�܉e��O&�ȝ�J6k����z�S5��GI���A�a���Ga? �Ss���]R��aRfɍw�c
�6bǆ��~�������*�����*y�l����i�@-O�2i�S��m�s��b>�5=`4G	y�����dn�S��-T��^�/�7��W�|�GQ��l�|�?�8r}T�j�k���
�5�N�@�䋜g��.,�	56},�z]JO�����ݠ��t�Jo��k�l�e.�	~�!Xy8������><���D\�|�q�Ζ�(�۪�[gH���(�ɳdB��|���}��|�x"x2��O6`�g|r�a.hd�Q���D�Į:��t.�C��A"���}]���'躮���"6�R�`~�m��+�MX�	&N��FSQ�hk��/� ��dł�ɗ��D�ډ�%,�����O<���7�eսϏk��0���ɣ"�_�)�cE�����_�4��:t)�*3)���԰nx�6k�[����%���m6��@��{R�On�+i��&\���񜉊�øG{f���B?'����S�(FZDw��I����(��bG����vܭ<�qtگ2�}�T�J��8*�0Ȁ$��B��D���һ&[)���ƺ]��	��I����fTTu;�k��̇�(�9�OX�l��r6RS�A�N�����H��V��ۓ2�f}_��*�$Ōtsx�pI���N5�4$��#L��u���FI��\��4��Yjx��krS���k�K-����Y�����+��*�$��s�Y�WR���ꬔ��F1 �sZ}%}�����)�cг��!
Q~C�վ�;1|���dvo�D��Mm�p
h�n��kvgW�c���	�oݍ��H������^wr��c 6��53g������?1�a�
��'>3f���z�o�?8a��\�U�ב���~�i>��i�ī�2����=��w���������*'�I��Gj�Ŷc����qD��2�c���{���.K������_�"�OS���`��(E���E��>ʉ7;��ے�&_U��I�������/'.�4T���/W�n��x����˵ݏ�L>ܬX�Z�?Wg���	��<�,����S��/DL�&��0�>|85Ė]����`Z1�>�1������B�; �8l�w6v#0�u<If�5���mY�k�_BV⸷��s�>X����m�rq$�"��y<��v*��,�.��Λ�L��.u*T�ɏv��`c%e�:<�o^LeD��Z�'��_e��$]�v����x����T%���B��B�x��k3��'�N�՛c-�U�ak���+B�n˷d���[��/�bA�#���5��e��\�H)	*��#5��1q��UE��0�F��Q'`��m��*��Ӑ�2��^1�h��wvbљ 
���K���ٖ'���������xn`�������@�]�C��-" }׃��V8aI��/�U�n����!`�;���9�ԡ���� O��4�9�@@�i��`���1����ʛ�]�"�g)4?�<���b�ʀs��ͳ��K6�&����5�U[���#mQ��"�m4aIn5�,i����$j��Jp�M7�.�z�e��b�D�'J�+�3�Z�����:�ܼH�Tg�����~��y�A�H���@�A���idb@H^��Բ��ֱg�A�;��%<�Vc}�F�'�m���,� J���I�8�������>�Mg��c�� �HOXI���� ��=����#:􃊚9	�]����={F��s-�a;����,8�Є�! ���0�'>�F���7���0��4��_�m��ݚrǂ\�~Fxv7�	�<G����0w�@}���5���Aޑ�]y�<$i���5p�T�|n�8\B���7�Sz=���V�f�r^٩|g�:*��L�{�I�wD�ԅ��F�㩬�)��ۍ���@��/��Gm��|��і��� �t��
!�sW��ᆝ<&R��ݾ|�.M)�]1��<��2c2b��3�[��p��c��z��\�S���_�L�� ��l��D|�[���Q��
�̲�G�N:��Sx�s�c	�/9(<=�\d<9��>��A�9D,��U�h�h��,���hw�t=�?3��勈�$s��RǢ�̆�s��L �l�k���'J���k���;~N?ܠt��ڂ2����8�ڑT{ x>|��	��:p�Z�}�x �B��d���uXq	N�r;��e2��b�gq�eD�@�5!-���4�Um s�>JvV<m��I��%��т̊eS봆��F<�
�δ�q��Rݣ���x���dj#���_�|�+պ�m�l9��-�
��������^�ZyF������y�*@C���oS�sKYU䯒�¾�Ì�,5ojA�ua#��.'�"���N�y
��4���y�*����'�L��� _{���P�s��N}�)�4�I��©�c,qoxY(qA��<����}o5+���R�k90�9��t��l�;	�Ϝ���բ��l[�j�)%I��qq��[]8�|< v��a��q�� ��O~6ӔxX�-�̈�J�r�# �ô�C;�G���/w�����%(SS
ҫ&����UOܭw���@���d�Hn�딙'�7G��_e�-�3Ow�,�/���ĄA%�V��¾gBxɻ�-�g%B�4����L萰�:�X�j@z����vAC@߀�	lߺ����DO4��mw�� ���/�ݻ�j��VB΢�5���G�dRI�������&�`��LϞb�w��]-�>��6HfA$�A��^p*�1�kk�^��@�d����}J"�{��t��L����%�ty	``�=�`��v�D�2����Q4����\��f~�v�u'��,�	���9�0������	��D�3�v�H2fA��!&��6IF�qP��is�}*��&AW
��P��ΰ��YL퀊lqLԯm���RH��d5u�D�fW�3U�.�H9[�^P��
���K3㐩3>��q�A���ΎY$yK:E�t������!n9(�r_â;�|��hD��U�C��s��6�F��&�O�,��w5�]�ES ���]ktT���Ʈ���Um3�G
��cF.�$�%M<����4o(hY�z%4CԌxZ0\xaZ�>%}GZ����\"a��OoB��I�m�|t�.x�bR����K�Y�����\\�a�E�wSK�M�NRQ���+/��O�?�2]]I^���=0����!����µ("�*�M��"��1$MtO���]�s��W��a"�]���^ݧ�4]����T���mw��"Vc ?K]�ա�H�2�15ˏ�F��+O�>��հgß�H�5�[Z��|��𳳩Y�Z=gZeS�e�#Mg|��:C����}�� �T�ѭ[��k���W�_!��Dȹ����=HT\a��6���>�!3�EŘ�����}��9�/��m}�Y������O�[3gr��n�'�� �jT0��%��v�϶��Q���켶]b�Ybe�v<pyRo�e�K-�&� d?~}Q�,�C*�����}�ή�Ͷir�6oP�$����Fs���G�a�#Ĩ)��z�9�������V�c�ٯJ��\�s������ ��_CW��AxU'�+�8�y�NU�d]��Y��J�Tw�/)3D�~�k!W���M���Y֫���3���v/���v.{��+L!�D;�k�\�e�L��'������+e��4����
�#���N!V��V3��}E�\x�/6�M�Q�b�Z�4|VL�e��PF*�]��,M��2�ɞB��N#;ㅪ��%!�}t�� �*��̻��0yyG�Zt�>�{H�� <���
Ϥ���.(괕����*���P���f�|1��/������	�z�(�8x!7e!�Gz�yő
�w�u����4��Q
��öa�ԣ�����E��ֿl����`1>'��+-����Na�UN�o8F��6ݻ�a0���z�cR��]D�>�S�;�j�/�O��U$'��|l�%�Kt�G6�:��A~?�a������^����`*ӄC������̌y�&���>�%'!�|Gf��Y��&1V�w���]0�.^���R�-�<�C|�O�c����c+��mi$(�P��׉0�X+-L��ѫǤ�g�Ld��M���,��{��qm��U��ʶ[	���f��K��o�_$��h@ݲ�?!X�в��㠗;���i�%--�����3#�t��Q4��M�PE�B���^��;�;N#�!0�eˇ��%2���DBJo;�`���ǆM8d뾵�;���tV���������W#1��$1���r3j�it�=V/����}��o&X�:�,i��Y�	�A�+k0��w�J�[���Rm%�/O���?���P�r��R�ȢzN_����'9F�}����ݝ�@�^��m��^���5�,�%���^cnǖ .3k�	�Iw��<���u�'B �����o�5�I���[ +#��̘�bu�~~���x�͘�e��7�bL /G�(�iz72U�HJhv��ի��'�lz�0��Lb�Y�l�[��5�P�/����ǯ���A���[��g��f�I���*�~�%KD>���Fְ�X*���I ��n�M-� Cw[��"Dm摥ޒ��n)�=�Hz��l�`*�v"/��PQɐ{��K���*ǲ�#4�X�H�3�p�F�.pҲ��ߙ�3��W��	;�z���;��vh19+��|K������&��v��3@_ٹ3�J l_���&]?��Y� �¯�����h�`Tr4����E�ا�<�+߯A|�"/�=��;Cwp]ZW6Šo��`�11�ޟ���|��o3g�Gf���-�c	�>�$����>��Z,�<�m�_S�_TmY헩!c��EV�r&���Ϊf�$=d�0cc0��ǈ�q$0��z��S�G��h�
<.= �R��4R�?��52oX���O.�!�Dy>��J�T=MFu����h^[�l���h�ֈ��з���\�p��w�W��oӝ���1B�P�۾�1���-�@�+� vсO,,0 ���@��Y|/3�`��CJ&���D|�h	�+\n��}X-����b�%�y2 VG�Լ��'@VlD��\��˩��槄e�Α��8ܭ�(%w�\8"|����8 PY�õ'��u]�U��]�$�����1��nn���T.Eڏoڏׯ��&3�2��LCB���O����/Y���-���j���$��Ѐ����
:?���9}�l'ڸ��ErJ��ѷ<�e�!�3ҹN�����+/�#q��?�K��+����?ko1k���k�L�cY:�� ����zm��o���?\�J�R8 ���Md���1��2���x̜n1���[V��Dl��q�L|/���䒽6Xn��\ɹ[�%oI.��Cg�b�\�z}w�z@o��'XE�'�:�,�v� U|�9xm��6֡�G����'^����S��L�M���:�]
���C���9RK�i~���v�'��zmh�����ᄞ@I[	f�k�M��D��5'��Bv��8����RmVVZ���P@$� /"�z�W�����Q=�����j�-���ކ�g�ReK{�	�����z��ߕk���R���::�`��
�����U���ŀ͢��-;X$�e�i�1xu�����^"�Ooa��Z�gǵ�� @�#�X���^
7J���?�T\�[���\ H@��������^S͜q�k$C�y�ޓ�!M�>��3v��tZ�W뷿|qQǆ�s�IJ8��ű�_]��/u�@�%��D���C��Q�3�i,��1u�N�1��Iz`]��!j0ߪ �Ŋ�Q��'�v�)��3������]
��cf������wj��8�`��E>���8�x
F���ʬ��{v��3�;��9�r���)�'jt�����oz'��N<@��ſ;�XX/<R�f�ֿQ��m���u�����y��ꇖ�S+�<�g�ۍ%�����ur�Uw�6#�0��*�U3i"�K����_�fע񹷯���C-t��OSU9�A!�p&�Ck�Ї[n�>��:��S
a}�$7}�|���LF��?�}qs_HF)�B�P�ɂ��nS���NGN�c1�N�'�:+�N��4X��G�5L�Ǩ�>~f\½y�ZT�ë�6�=����uTK��3cT�n�'[�Z�4�ϒ�uӼZ��ө��V��k�R&�<�E����6f��s<2�W�r�����Wҍ��Ý���!y�