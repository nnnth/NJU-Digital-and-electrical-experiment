��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��oڀ��ՙ��3!����d �,9|�;��z��.q���{ڧ��U71��}y��|���Q����w��HTfZ�<�� �v.H���G��"��z'gi��p�d�FA���4w����|��*g�ߍU�i&ߍ�j�|�im[��eV�pa��*Lp���dmv���j-5=~X��$� u�\s�����N�)!	�*|C&;�騸��tx	�h��xE"j�Uf ��s��p��!;
��=7�r�fϵ���
-��g�-A��#�o7}8�[�;���Ա9v��~��DB\��#�ӗ�/m�$�݉�WS�ux�S���^��T? ?D�	�MJ�׎�d>�#�8j� �� {%Ր{ۋ��_/�q����Ď$�+CR��;�^�I䧳I�ԍ��d.��B��R�qT���^����!o�Tʟ~�<#7kTݟw/�Gy+&`�k<Q�����y�J�P���w��Ӽ�����̼�w��D�!s�R3��0@�T�9� �eM��f43�^�1՘�Z;�rD�簽<��J@(H��\�dM�sv���r�;
��$l!�*A�7���z�4=��|2�?������B7�:ֽ�1@����=Z�Qg@�=9�����p?�v��ʄ��e���%86���嶒�e�D$gS}A�t���}sG���m�.�{���}+�x��U�G� r ��ﷶ4�o�0:�~ñ�֙���1Ā���Ǎ�~͖7�'m"	 ;�ᩑS�,D	��qG/�%����b����85ɋB���4[��(_�A.��=��\{*Dk���Th��G��0Q%#��O5w{.,)��g=�yf1L^%����`ǂ�R���b2G%{o����X�����%YQ����[�7Q�fh)l�� t�Բէ���HU�!7�������B�7��_�w?�M �O텿���F�2Yɤ,�u�+E�����݌����[=l��&�6N��m�ƟbI�m�����7|YG�&8"�5��׿/+�����E���Ǘ�y�B�Ȉ�	9�@�H��c{�cV��<r�(���)�_��O�ORߦ�
տ)��+3x9�H{v"5�,�B�Z��K�dl�5��8`�uj��'>v��j�ypM��]F�6!��Wk�IYa�� ��Fȸ���'��褃�g�H��W�v���}�([��$P���8�����2&�T�q�N�;`����v e�19V�<�k�3:��~?z�2,�l=�OF��)�~yj��<�M$�\ӵN��w�
&�)�H�6��m^:�Uv��\����&�fF�v ��1�I�r�w)����4j�ԣE���v#��1䒴�S�s����{��FCⓜ�L��kw��"�ٰ�$@�u�EeK|��rP�gqt���E^�%�x�5}�2�Ma7VJk��ۀȳ �Ky�{��$fgvg�}m�%����ŝj�
�U�5|�DyXo$��R͜'.NO���U���eD�(�<R`N��w矉o��>���CQ���g��pf㡻܊ژT����3�l�5����7�&�(�t钮�J6$���W1
�վa�>��m[�S��d���hkqfշ�3I��)���osќEj��Af`M6[����ЎS/�zn�lƆ$9��!�qR@���ޅߒ��-�� K;5|���O_�zM:��F�YJ���r-UN�^���O���	U) +�s�V�bLE�{	ܤ%�ڎ�$�W�r�%��Md��/�YθH�5�|�<�����L�m�Tb���x�Qu��udə�I�E��S�rJ2����/]�:1������szea�e��9�S�L3O(�,{M��yh��X9��1�i+6�����-�>l����P�J������>kT&���1�M7��e���0'l*3NV������9])����i�W�� L���c�u��O�A&���	i�[uc�{����N^�*����n�yd���m<�X7�wj��DCߠ�0�����z�?X�`��(/B����$�g�v�aI�`�Aפ��
�s^�����ST��m�d��ěc�
�D<e5x���l���T���+�!��A�?kP��1[���:��E'��-�_,m���ش�떐��!���ജ�6�G��4�zq[�"=���n��=�#&����pI���\2�@���s���\L�P7~�.�5���*��s]����P��g�H*��T�r��NUآ���$�{̋�����ΐ���e[�j�WE;9�h1��%�"��� 6�8t����>J�VQ����ƺ�ֲW�Y]���q3V�=|��-�L����(��:��Y�Z<���<����X*R�2�tKc��A���v�J�!��T���scE����ڬ-�o�+PLeS%�F��u�S75l��z�WH�9ܫ+G=���{��O���}%$j�*�9&�����Lc�+X;�?E�j�����& �-cՉI�
� ^��h�ㅁ�)%�q9ͣy)�u�n�s$ywxeC z��_(�_X���/�n�xy[�3Db� ���Wet���֫6�	cWD�:�C�c�{�l� ��[�i��Lh���HS~m썝���8?����J�<�ɶ�je/[��C�/�ۣh��;������;��i��B������5�vc>�;�ݘ�-Yc"�|�93����y#��<�(���!��]@��j�V����={8�o�=��ă���DXL%����*'AFl�9����	7&�	���R�A֨W6��soC���y�MK��P����̳]��
��OH�8��*$�����޲hއ�R�Z�0�Z�q����hK��9�s�d=rJG�L�+:�߬�����Q�Ƙ�s�kqw;���Od�����3K��1�	�T�m����_�;�0��w�R��g�tRΚ��"�do�g���l��c�'�y÷�X�o[���
�.��b��m�8�x��{��i&��!�)�L��Cc.glW�����un�ZN���~�׹����8�P��(t���A~�J�N�T�V���%sʲW �K��o�ى���W/��H���WXjo��1��,��)kb~	y�%�?�gz��Cޖ6)d�I��q���93�ap�QD��6���q�`�M�btP_m�nŎ{\�S��L(���kF$0И�%2ҋiW��N�l�i��_gbF	�v�ˁ���3H9�Mγ��r�:J�%��3�t:L�ȜKsQ_�5�=�\��;��SX^ȹK���[���2qJb� ��@�S&���A[�O�����e�z�)z�7��|1rN�o��b0�p��A%�H���8��ϭS�t���v!���ʍ�N~��k�ԙ�X���o�Ld�.�).�6\�Eg�t��3;��gLdٔ@F'��O,�q*����Ƌ���!ꩦO�o.("��v�K	��>�^�����i3�4Q~,�L}�=�A;��E$���d;}��R��k��
��`���0_RXn �-;g���SZ����>Ul�.�wQ.�b�6��{ф4tg�Y����m�JғVD�����`7��9x1���}h|� �=2�IY�y�1	���vS^G��H �
/�`#D�t��EOR�|@��h!�'����)ݧ4V&T�϶������I_�v�S1���%
��K\֚�/�Y�`u����u�T���BH�D~��Q��,��%���B633��d|������T�������=��zz�،��#�tW���iN�/��Yu�ܗ�-lE�Y��̵]�Z��'F���Ý�����eM���TD4[��H�+��A����� ��+����ר�U���xw���S�e��˯��3�"ե���Ź�22�q��-&ët=��M)'��x�-uh� �����Y�����{���`���ppk\/:��?��������qG.� ���L��C�@��)D���X�M�
��!~��s�|��y�{b�ԙ�-�"�F2�6<��������8s�Pm~��䒕�˿�T����"��O������!x�[/c#���d"�k+�ˢ�LK���#�E�i�޸Wf[.D�%)[�Z9�����h'�s�.r���� E����&4�n��6�������y��RZG�(�q���3�b�)��H�nS�3F��Xʃ1�[���u���9S-\Ħ�'t�~�����t ;Q�hH~�wT} �x� <�,H�i�U&ǶbE�C�>����/N,�"��BNKѺ��M
���h,3��Ź}^]c��R�:�)=М�˕T����Y�� �Q�(�u�r}�ĴV�A4�~��Tl��,{��X�gs9�gO�#��V�ŗʄR�^�]ʍ���pk��ը7sb����c�9mf��-�~��2���D�h����yh�*�Ż1y�".�d���y�&к.���ڦL�*�5d9�A��Zy��No��$�0s �"�	�x�I>�)�0����f��}��p8q������q ���
M��'cy5?���N��� 28�]c��mƞl�P���b���T`�|���8�LF���(�K��T��-��n�\�tw*y�>P���.���nR,�Ө\���������)�r< f�z���gE4�Ȟ�A����"��o������,���c��T\8����un/��j��m��(h5 ka�fL'��h����L?|2�VX�W)�	oT��WT~��k%���uאi%���Ͳ�L��H�蝣%�Ee���J���&������y!�O6!W�<�m��uBC��a �I��Ǻ>�AE=XZZ�˾n�+���%��,Tv+����SP	74K����%�wg1df�mƕ�,j{��ychެ���n[��q�e�U>�@�ַ���T�+%���:�:=�BѭXT�kOw
Y={-�\�.N�\�K� ù�ݙ��a��r��݋T� �|�fR�r�f(y��O��7ڤ�Aw�S�<��m��yd�n6Fex������F���>,vԵ�V��/�:oo���x����/�ư���kD37��O3�y������V5Ӑ�e������jS�6��N� o�1y��NZMc�R�sp�#����W�MX
7sk���9,����|mM��K��e�m+b�����hF،�O�T���_�Fx�#����Єx?�z�ēa��iΫ�W���Ơ)iթ����֋o8O�9���'O�H��:5�-���ly�A��+;�{'���%�����n=�;\�ܯf���y*��\� V�̈*�؄���fqʖ��~٤���,WPS�k0��q��"�Y����I�k����nٶ�\'�k!�=�k��(�a ��'ߕl��D�D�������ϣT��ڽ_�x/��u.x�4[P�ܣ<OM�m�n�)�x�~ǌ��I���o��n��j�(�C�����=����k����z��K#P�[,��;Qٝy��@��e���8�Mɪa���E`J^����]LVZ������=�K#U¿��Ŏ���z߁="o@xꀠ���]����K�i6�ݪ��r�p��\��8�7�0�gY���}5ziừQB-��Sc���u��R�]��Pw����K���(�O�W�����2�xRgo���wi�5;��T<;�s`Zt�,��1W���qb�s3�>ݓ$���J𵾻��oϓ�~�!�0��{��_Ƌ�xŌ�}J��M��͖�Ҧe��EHo9^�_��:�XOi�_�K����u;��7D
Q|�CM�sUb�1y��^�#��F/��VD6��E�9�]#
�*���o�Y�ۉ�8�����\'{O��d(��J�x�o�A׬�"0B2�IM!�҂c���%��f)�gz�@f9�L�S���Id�PN	_��6�-`~�vω��A�5.!j�}���62Ѷ�s�����d÷7"dW�t4�2<�{���WD-/)s5J�4�f9J
�$[�AwQ�O����Ptv@
�y
����Y�"F��������/�`.#F�X�lȧ7�E�67��vTK$���B���G��]Ɨ�!0X��뤄��%#�N�H=&�ݴ'��@
�����E,h�r�k�6EZm��~:j:(��
+Н���&X����i�ֵ��l���0Z�2ҤN)����֜��;~
OG���{���Wg�ޠ<5m���rX�w$��5�炈}b�/���=�\ې�/ 9��<�+������K��"�L�U� ����C.t��زF%䣞I�eI�A��I�IR. ˓��"�F�]}��oo�7(:_��'�7������=��G���>�!�_���ҚF�鈊Q%b��oc��J��-q��м=����g$��C�(�$@.z^���97�Q�O��U�<�lr��1̩e�ْ�ۡf��H�%��ٝK��Mp'i��ƙH���Ї�{�q�C��'�Pu��X��l��/�y	-F�:�gGH��I}1��2�nL����<{ >`*9l�yT܌��,=r�=����y��=j(�����W=Ը�ym��h�;�g�&?�� &��Ԣ������[$ƻ��ԏ��y��sq6�/bn��ڦ�W�C�u�1��e�פ߸�k�'�,���,F��2��B��9��S%;E�c=D/	���!�<�{��$��OZb�8,"�
��=#����/]�Jr"�vW��e�@�
��k��d�?�a��5W��j�
���P"�'�� ��H�rWy��m�ȃֻ��t+��C�Y��$&
�3����#��=��̹�L�n�
����[��d�e�Pd��ڡd
M/���4;�Z�c߉<wu�!����R�"��+9�~�Hh. �6y��W�,;d3�!sv������Qɮƨ�yw �q�&��Q�t��S�6�n�LT� �L�	S�� p/���!�/�a�m��վ�v(�JW�X���g���jSesV��s�eC�^wUF�+�H��h5W�ӟ�J��0v�H&=�a��@Y7.y�@��ͭ�𡱅S�G�%��ŧ[���,������\��Łm� ���2>c��4XbY�,�	��D�[bҨ��r��{``���tX���P\-�xM���+Ҹ;_�8X�._�����SF�X�F� Y�j�Z[�&����򠒋^��8m�"�+�d�)�2(?���FWh�?e�25W��En*�萎h��u'���*�JH�s�:�U]ɭ
�y�!zhE�k4?E�o=<dW�>@��� ژ��SZ\��[K˖p��gn�8�o1�>��Az��{wb(o��?2Pt�H�p�j��O� b��zdj���SG�vZx!�gd�q��]Z���
���I�d��	�%mn�#��pE��U)]��a�,T���-m͹�f�cW1�<�q&�f>}�ebǏ u�d�xA�`��<=j�t���O��D:�Zri��6o0ܛ�N�Z.u��2�e��n�'wn7���}�~�wD|2?���/�Q��]��J"h�Ց8 ���h��E�[�HN&o��9�dp
"��-���.1\"�C1t���9�7W����O��˴��J%�y�φ
��C�!�6�qW��ǁ�QY	��n�]��n�h�o������{.�!_?	,����e��d�bi� ��W\�L��	����Z/��M���g98R��J�c�pF� �y�wS�>;�e��om���>�!�R��F�¾���a���<�����< H�H)̼7�%k�aT�NN�`��ؿ;a��_�p�k�����N�����!���<��C�S���Q5�N�p��%7���RQ����Æ J�z�f�A��hQ��.>�~l��Z�'��"��gr��+�`��
�OrG<�d�Aw_8���ȃ���@�_;�C���I�$�+`o�}�H�hE�^x���UQ--�����hqr]�Pq?E��	gp�8CT�̉�Z��K�:�;��"N�~�`�)� _J�j� ��\����0�N�
��>U��o�%я���B���Z�����ol6W�x��]&�P�'�9����Oה�H�X�\����.�F��(�wR�:��Wk�~��j��¯D����H�^QF�P��	�y<]�9�*-c�	A�*�˽F#����Ɣv���|'�kY�|;AS��A7��YJ�`u�4CTT����2��R+h�t	Y8*��}ɚ����SN��2���@WxT��%��ǿ�����x4��ID��P Ɯ��w5[�kq�tX��{�G:��ӎ�[K�%�b�ʱN�~:�w��	'�)gD�̈#��G��hMmӜ�g�k�c)=r۾5O�Cti��~�$s���A��h����?�6No�O\ԯ�h�-�o9#�����M���_"g��Ɇ�c4�,e�EǍyx���\>^��M�6[��[2��"�%��͘��׫�2��^����� 8�B�^�BK�X�զR�1^g��x��}�O�֫��c��@��ǓϏ�Z�~]mQC��
TT���E6~B���G�%u�Hp�zk+`*�O�4��>�Y��#l�:��	�7�D���)�%0�-ǣ7��:�w�����4��=�� �kG����!'�Q4��׫o����K�d	��b���E����}���s�PI�9_aP�u��ďOFl��p�/��~�><������$�´��X����xP�X�ɸc<�_�r��4Z�mz7G'�P��K�s��T�#�w�R{m��}���£ ��pZ�n��=R=ӎS���_�j��@��ػ�Ș
�=��Ƴ�r�ϗ�f��G��F���+4�tH���-��f-��z��-	%�\�]MO��_�%���Mz�ݻ��ְȹ�3�+��$��3�rSq��y�c���nO�.}�N��[yW}nĒ��9�~07R�-�r��E�~�P�䅝^](�,n�>iC\��V�X���F��Β�Y��n'�Y�M��ڻ�2Nޢ�vbN=l7���W��)��8��D�g�F��lòQ��v�Y\���p�'�_lư:k�����\-�1j��.�_��������O����|�.�׊����� ��g�E�<q�Bqg���+��������A�ױ�|�ͥ��>�;AP}���h����;�ҭt�Y�C}�Y6.�	\QgA>Fq)��$��2�f��y�J6���˵Q�H̦�Zn��}�6���n�Dg�����
Ђ��bm�oY��1B��ֵnLI�*T^<Phb����M,y&�#��L"�MzÄ��MJ�_���+~�.�z��<���+��  vvT�?y��^0\h9��>��Vve��fX��L���֘к�S�U��W�f�k��/��O��(��Fs\��"N,q� X�׷vR$�Utn\;pV#ӎK��m����>>�W��
ǉ�(��q�X&���i���,$<ƅ����Q�ڏ#y���"�l�\�`�%n�xur�b��'��|�~���!����D��8���q�#!@���cӭ�xQ�ܝ�����Y9˃�����Ö���d&G�0ʹP�Iy((st93wq	�A���d^�S�Ny�r)��"�M5�\�>�-MK�O��?5�'���	� ߦ���D~��LR�9����fz�Tk�Sq)3��"9K���B1��<���Ê�>�T%;�hc0�Ʃ�*�28�n����
�����Rw	���K�v���xi�?iM�c��陮e�md$��t�1���dP��=[�".�q� F/�R�������~!mry�G��o�.m�D��q��FVd<��� ��|�����Mn�ŭ�� R����]V�!i���\��
f�|�i�m���tr
y��C\�b
4�(��$�m��-3�$�pFˠ�����DD�i���0����c�p=�G���v<������fj�x����/]��Bͽ�b^L�@�_�,�c�.2B�	Έ�xT.��Iu�������[��*���A����b�Ɗi2���	^�8�#��z"k)[���:<g�i��v���q����lڏ��N_�؉lҀ��:�f>�p�9vg�Aօ��4�Z�~�џ�7��o�~�`�hP&�ap���S���b����bG�}#Aʫ�v#�G%�K<_������� $��ʛ�{�o�E�R�N_�H~%{���ɓ!ˌn/,~�X��?��i�>,�s�.�?��!���j;<�܇�f&��h:��N«��\��|���w��{#�6�0�*D��:8�C�P�Qj#S�@�����I�t�ԭB`�1o?�]M�o������J@��b?`�ܨ'�*��9��>� �Y�@�êK�bϝ]�%/:
Mw����@�&&��5OE@��Q��#:F��B�A�?e����*׶fǊ�h �R��~;5i�{[֯gIP�{o�FA/A����D�)�F�:#�*gP�:����~����V�b�.�~j� ��n�v�ہ}V0L�ɧvu�-r<!�4��&�N!�m�!���l	���&��$[�D��JM�W�dЦ���$���ri���Ke��n[2�m/qv���=4��'8�\"o��Z�U�qI�lpu�I�T93�qR�&�z�2ֆ1�k����~м�l��	~/����.j'�X�Ɩ���7_wsQ%���n
���o����S�����.!8�<���Ѕ�$u���jˍ�\��.�<o�'`�� kZ���:����@R���[����w$��h�R�!�[�{�Mj��q�W��U��a��e�<��丞x4�(��lB�G�g��l䚗�������B��3@g���^���R�|�e�R�mԖ��ڜf{M�יU�Wr��
b�[Wo���D&�,��>��i�e1�H����H/�ޥMv��@֐�?�:k�|��xb�Y��\�V-��򃗡'�$��	�ȵ�k^�g��n���h��̝�@�1|��aϨxǥ������. GƳI�����u��Q��_²�5��/C&�~9JT����5��L���3܉�%��-��Zu�
η����K���q��/��!�6|2�v�e������p�2����������2Ѐ3���E3p���jZ�i�!ҏϜ�b�AK��؊Gh{QPo�����h��X�,��SF;ht;�-X�'�(�.�7��L��"���z�F�Z�{ .m6��/-W����P���K'Ŝ~z}2>{NXI��$��#���L"�yb��~����8@�;���\O-mP�]wA��H�,Đ��6v����K�����;/x�K_~�����ZV�7+��������d����S��h�>Z:�9~Ac�����`�"Bl�r��q�y��V��Yh��wR�E(�_����E��"�3�_#�'���e3�*�/��~[
f��2�q��_�`�|��V���1�O�Yюn��Z�Z ��i�覞��9�ٓA	�<D�6Y#�|�j��E�i!�cj�cxã�Zc�Nn6���奰	6ܚ1l�6l.�ގ	�4�1ɥ����ꗓY}f�[,��!,�E^Z�@rҗ�~f�
BO��p�W#:�)W���Q.�6<���&�.� �� "��;�e�dY�ق���U�3@E�Cݰ\A#雟\Y&-2�o�ъ�}�B8�^r�\�:x�K����v�s�cR��R��	���SR�����ч��xq�S8L�&9i��7��oOp��H�ψWH�a�����Z���A/�u˴_�{��>+��I�X�޿�@�f&}�p`�Zb��ݸ��yK&�p��A�iux�n�b�<�t'�����gU�������3j GoS���Q���[��0��U�៴Ą{O]�h?/o���T/EMG	 �O��7
����$���dy�~I�ѯ `�#�, �|$�H�I��&(�C�2̬� <��6��ŴVh���}Q�n9�i�o��5c��8�- ���"����V�ә�J����-bet�E��28��2�-�l�9�va�K�����OXf�?P:3J���j��d�v>�9Y��B�z]rx�IUy]��Qh��1�����o�yrS+W�b��R����g���.�^���3R�>�ۋ�ܼ����r����pfJ��6��~N��1�8������~�̎�RD�#��8�1���E���Eo]X�.�<ŗ�A�����Q	e:#�Y�$�I�%�i�Б:z���Q�7�D�y�H�RHs���!����a����fi�O��ŗA�f,�4�nY.7��Vo5ʁ�Ē�Ǿ��X]mS�g�;k��?W�]�uF|�XRlR�\4L��Ɩ�X�V�/#�$��N�Bq�kVn}�I9��R_�7�OGw��ض!�Q|�9�� [��gp���4Z���"i�wƐ&�5�n��W��ϡS�Z
�m�!u��{	�l>V��u�����"�BB��L^���(��$l/���Nn���DZ��&r�!w�il�w��UC^f����YP �cr=�汾|n����9�"�<�E���@ �h��!`R/�k���.�����z�T-qi����q>8��e���
.s��X5�Ϡp����y��4��B��"��2�|ɪ�NK+����n�4���)����Ѯ��qr_�l_� q\Z;�f�z���/��O������{8��a�T1�?|���`bԫ�󜭎u]"E��V O�Ԑ����\��$�F�W����q��q�����l���T	n���l��c���z Dq�Pi�aV���#�G���c_̮ۜ��L����=jh�h�ߖ��;�R�K^n�jza�.�R0�Sp�P�5㰬�\�v�2>����%W�����$de�ث䜧�ܘԤ��[�ɭ�_'�.���eéڜ��j�L�z�qn�}�AUh�&�C��IB��߯5F�1�]ei�"�!�"ʫ��\Kr���@xL���-���x<�o��K�� �pKTf.O\.��5�g��}hlO'��q��5fġ�d��I�ì� !_�$lm u7��������!N��#�ˆG����f)��=��n2��6��t�.G#���G�O�.q��c}���;/pS�n�J��6M �G\�<�>,[S�3�ŖWӅ�"â��3�լ��"�n|��7#��/�k^�o�����uB2���ֽ�롓�P�n����Y*룀ռ��sUav��o��������� �)�4�7�_e�j���5y��J�����>�>ߋ�2&]&_ƿ�b�
�l1�nFB�G�,��g�Y��g�?�k�L�H�.�k��ȕ�����#���*/L��'���~H�8��ɨl�Il���� �yI�iJ
�*l�k��W�e�����x4�Z;�V�
�^�hqq�}H���$��P`�7�Ϸ��� $�9�t�VT�Q���j��@�e�/�}R���o��kL��tO��/�(�Zˈ��;��29�=���4)�0��{�9 cn"���Z����^���K���j6*j���%���V�)��I?ҷ#�yz���H�:`*�F����6����$x-�啌���V�.u~�ET,�+���W���`��*V�������2���%� �1��3���=�����R �����Y��`�}b�/˵�,w�Fa�}�lU�wJ?J�cmw+�uϴ�~��Bƹ�^�	G�ˁ_LRB'7 ��G�ւ鹒"��iq�9H�.� ت^!��v�@r) ( Qyن���}y�5����Q�֣V��AZS�������D�ё���0lI�����@��;>�������Y��k%�s.���퓖Ӆ����"�"���ܤ�F~B.j�Ŕ�&���� Z��]u�]�Y`(��ˌ�u|/�%a'����X��M��6���P�~6׈��0���U��_N�j�H~Z �O���o�' �_��V�3�� (��8�d��o�֊ǣ�F(��?ڔ���^��٬��IЮ
5�ƗM�Z�Q	��N�"�#��,l꤇h��/�G_Y�����!�N�
����F�HO�+N�YO�fY���� ;}��j|�k����{���HP�R�_ݰ�I8��h�%@ip�l�f�U�VGW��Q�o^[��+������iD%u޵��"p3���&��(��dj��{����ԉ?�F��nǟ�R��]�ه���|if��j��0V�9uE������3d.����Hw:˒�w'�A��/�\f�V$�8Hk0q�c�A�0�<�z�gX0a��L�۞)�O�ZE�O"mB*=�&�R�=��&���u�����m�,S��-G��O/ ��Mg�%�҃&�X���mU�zӶ��ʼ�Mo�k�5_����&á3�ǜ���Z����e0��ϑ��J��n��9q�xd��잜r��/1/
3rk���`��^���Z�w��������遒�����&<f�����^|�7X��\�3h�����3�u�rJ��%�)=٨~~�i3�5ޝҡQ���̝���t#{nn�WT���{&y� ����^+��F���a׍���
�	�FQs�wу�Y��"$f���k���/ ɰ�B�#SiM{�	L��s:���8�p(R���I(�E�ya���l���<_5Oy�赵��d��Y�a2o	�72�5�V���[:�j�!�U��Եa��m�a<\Шm����O5������wzg{�����ȉ�f��� צ@��B�͚*ش��г��>��c�Y�ʛd�K��.����7�y���酳��D�X�b�p��d����Ot�W�;ug ����:�Z�D�>�u��C��k�Q��>W���I���cv,�SL����5�s�\>��+zH�~L��~�qC��u���WG�s)�(P�0l����*V���۩�Ԑ'���*"���R"������0�����Z�I1���Cy���t?�I<,N�C�����hkp1[X,Z�;u����4g��Д����n��\C���u*N�������ϝQS_f ��S����u�Ay�R�s���7���rB�v�<0����Hh��e�<	�^\��/mz���G��_�j��t%��;,��%�T;)��q���?�U�a����)za9쮯&�3��H��@[�A�;�w�A��w�8=�9�a������|p��}3���J2P�DG�4~ԠD�&�ӝ�|1�2�;�7�A�=����D~��~���si ��9e��q
�*�a�ˬ$|��,π:�v~?�����쨘�?z�� �����g�q�����Qx��[�K�Ĳ����_75���=u]����W0 q �3g�&�"�r�ȡ�)f�����Ҩ�3��M�Q��7�����i-�.~�i���U�2�Z��ٝb�~�����X��+�Y⭼ֳ߲�S�����5�K����Y,܃E���É���_K�7��@y���toʻ*�g��=3C@�oؼ�g"��`GB{�_ ����`��D4�i� ���{���#چ�����ME���H�� ����:.�9gOUw���e	5v�V��?`��檬-�l������C|e6�2�׌���-��a(��2�<���X�8�ڜ�sɧ���e؏���-�zZ������@���T�.]�q)�V�y��vB�{%���޴^ƖG�
�AΗ�Ad�C�7���iM�ɚ�7��Hr�,�{��8&0�۸���՚��_��O\����R7O{�@^�*�V�p&�$qάem:��q�A�8?SD�~+2&������_FώK�/K_�̴�P(��=U�k�tD�����g8��);���,@��7����������٪��:�������++�ΠQ@z��=����5C7��f��$(����L�PC�x�y����p��O�.���LI�0,��?@�>L�%���o��-W���%G��wo2G�¤�A�W�����lۢ��Im`nX;��i��X��P	���x�[~�R?��j%?Π�&_�y3YI��o��$z>z���ݽ� �Ҏ�~�
�=X��G�����퐭ARE��P9S@ݽ�+�?@A��Nb����eu���Z�>�9��!zU��Uq�՚�H���A�'v/�1M�����r�#�c>k~�Cl���0 y�J�%?+W����3�<��\͈�Q&o����,�J����ʲ`�/&��T�7������-����U; ��Igz�'���2㣁��t�Qv�E�:����z�3�W��i�,������9�*S���A�����A��V�.�jz,\�x�W���x&��,��U�Py�A��5ƿ7��8v]���2t7&��JEmUcA������#4R�&�&D��f��H�s�J?���$:YR1#N�[�B/+�TT>�kp�x���P��|#��CP�á��������'\�`rΒ�&��É��A:���O�bq������ Xh�\��w2~���1����Jeӑѭ���\_����GK6�}�/��
1�����}�KK�T�����1�42�b>�z	Go�y[@L�fF�>�����RÄS���_��6�n1�&��A��ғ�4w�b:dc2��wX�
�wY�q�z���4�����Z��V�3j ��z�� ��u؆��#/����TXDi$�}�ȠM5�/C�6��܂)Ʌ�TΕ��|�'z3faIX4�a�)�������9�:�``�߀א� �G��LC��i@$<������5DS��]$��1�R/FIpZ$w�&Y�P��Cݱt�r>䛟7�ȹnSA��1�x�$�2a���?ȴ�ₗ�iqiy��(
V�ԆF�X�_�&i��bi��wl��t?"�������\��z�H�F�9�s�5�8�en|�v���L��8!	�^��L񊣲Q�i1R@$�aޑ�糡�����v��>�d��^.��[c�Ɉ�|'��ny�L]����C��?~��$���9�,-�"��$/ls�������%[�'���ar(!�� !��LI7x$��	�MNҐE�d�«1^�<�B�pD�3EC�=���s�>> �J5�Q+5rf%���,$~%t)�N�:�ɱWDG2��X���ٽ�j�b��z����_'�!U̡�.����T6��+�1е�9���"<x1ݡ�\-�z��/��V]��F�ƽ�p����ZAũ�α#�A©�_���X�J"�c�L[�/
P&����3�����Q��a]�^b��_�)��ˈ�ςq��&�^�l{1�o�t�������{���F/��tl�9�L���,�s�2?+RF3��)��j����(����!X$�A���,1N9�}%TO�c�͘@y��J��r�ؑV�_^��Q�ǀ+�t��1�#V(�>_HZr��rI!�*B��x��f;�$Kq��(֠�*��X�R�Šޘ����=��@z�N�(C.��ϕ�?I�����Yщ/��rp�)tĚ1x]ɭ�����"�Cb�)[ȁn�5\{��S�$�����+�w� �T$�BgA�R׀j���q�U�U�'�����owD�����DX�@Y�1_)朐I���80��b�����]J~��Q������<'��Zf6�ϑ}���<���{��{l���xy�j�EVhsI��q�$J�x0� t�#p>�'Ѥ��E�l�_�v��+Z[Y��8�H������c���6����F_LX����SL��T@~�44zm#J>r�V�����6��w���p>�>J�գ󊙕�ub ''?O�<���fl�$��ӷ@��I�e�������%D�[xX
��D�`渽^�a*^�Cv,Ø���S}�34�Y����W��{�	�ŢrRM�QHw{�'��Q9�G�4!Ӭ�I��zJ� �;3i�.�%��")#�~~�*0Dc��Bъ�����2W^�\��
����g!�6t���pb�j1�ʰ�>^�W��u�Nt������v���0.��68!Nka�uxR؋���$'�zxkR��L�d�� �aA��{q���<�o�V ���0'%4����b]����x�����&aV��^�ū'w��;���\��Z�ɠJ�ڳ'�;����J�O�ݞR$Ž�'�O�a���puC�b|.m�T1<d�2C������s�f\�C@�}�]�h*�\eM9^�⍌]����C`z�NH��v"fb�T�޾�:amy�X�}С��g����5��Q��������~�0i(�k��U�f��B�k�u�<nj���W�&�[����Ĥ"������j�p�ؼ��o9x�J�`�NB�,�Yq�6�܄���G��3T�ޟ��������
�����U൹�������w��l��h�Z�ʣ=�|f����|�+T��|�h���A)�r7��"o�+�aݍ�p|��^�'8�o�ql_{\���M�R�dQ��+�A�`��p�BN�rK�b�&�u@���mT�3�h�9��I���6m*I�5��NΌ�G�:�i�OU�*� �H�\*�z�R+$nε�8�Ej���~JE@"(7�y�B�s�Y���H��H�3�-��zf�F���{�3o�ӝCc�MK�:�bSE?&��x�/�5S,U�ؓ��y�
��aTx�O��&���ت�� r�ں̠E-���$sf�6�>c��
Vl1�����wy[7��5�+ȹ�e�rEƢ ������R��'^�����x39��9o]3
����j��넾c!�2�W���(�9��
��莶`���eT�+��)5s��]�a#8�bIA`x�ז-�������|��X&��D�	0���u� �F.�gmn��ה� �2��Di�_ϯ��N~��}��@�7�E��]��mؿD�#s��;xXp�&:��;<};�K��z#�-�`y�*u!6^,�h���4��0�!�p�+�����yK9#c��ő��7+@�%�k/[�(vG���fkQ�g(C�dl�J�f�J5e
+���g���$-�.�,�Y�&�tB�/(��m�UY�ֆ�b
B��V�����N�K�|}�������n� ##�������~ES��oձ�wu0*�%0^b�E�h�����'��8��{F`�����} �
!]������г��l��3��ƪc���Fd����5x��EK��#����R`o�U�K:wC�O����&���>?�G��lH; <*����v$hn�����f";��:R�����"f��[�HH���@�>7�!�~�T�p.�D��]��+=�TC�U�KJ�1��s*�a�,��z�5�?�Be�ש�ߦ���¯J0DgFk�#��w�2"�Q�W��������xt.;��RV�O]^����ַMf@��&�|�>UG��+}'{�g"�Z���ڬ��(y��<#4
�{���LW#�̋I����d!�������D��۽w�����|KY��qx�T��d�&TO�n2�A$'z�.H���
��5������t���4A0u�=y��j�ꠣ����ʇ<��m��ӷp+c2�1Ej��țC��KrYEѠ����T���oĸzf1r��D����"�Ɏ�ڃ��D�5����I�ېg�č�F[�����3� խ�����X���3Y��֎��C����;xÖBQ����E(}0|�Y����hr�2���KS��=�V�p^��O��WTR8��*�f�}�<+���[�Tl�.���Y6ŧ��(�����􈉄��W�X�wY�E,�u���棃��rI�	?��S*�AG�'T�ظ߂wS;o�OKE�7�7Y8(��3RҢ��(X�l68����V�_���{Po���=	�A�Q}C���2K��O"8q���X�f�̧��sP�'��g�HX��n����]1�AHY���8����)��M�4�{�'���aC���j]��8S-�?��:o��o1L���쵼D"��xPOރBƕXR��ۥ�x���M��-���/Nw�#՘Ȃ�Syl>e�ɼh�\"AQv$��V>_՜ڶ���p⡰^'��*mͺ��2i35OE��� �6�Y�&��Y�� ϕm��d�F�[�n� 
h�������LT�b^�j��ӎ�?u�;�"9a�yy�?<�$�?��kMk���ax�f�`�b�)Gb���KZ�=�n��uWf04u����U���%fk����iʏ��Jk"�����vɹ��{f���ý� R
����uHq,��^�~H��Z���C3��}.`Rh�����mbHh��[�լ��5�f��Q^~,�G�>D����,?��+�թ*"�k��F�{8��ګ�no�yrf���e����s p�a1�Q�)���6\@�'	�8�^��]|��Œ P~�s%w�:�j0.�#� i�A��|{��o���r�/}��+�Yb@Z�z�=��6��lL��ɑb9�N̲no�J�2gD��y�Ff���v�#��\�����J���Ȕi�fZ�g��&)��^ɓ�{*Nlwm�u�Г��.N�Q㖡N+-|��C�t� W| θ�
ӧ�R6���b'�P�<���7�=��~5�lK�U�M�X�|��-�4�g�bx�e�_�'�[�.��vʳ��AA�]kO!���(<�Qj����d��4�(2�o6��r��r�[��P-E���1	�������Ғ�r�z��DC`MP����8~:��ĳ�|
�X�����>�*iI��w�t�
wA3vâ�5*B���"�K��I̖qj�^>��������Tо])
�l������P���$����'�8Ho��h�+��K��|��FqI��!P��$s��Ǔ����`��ef��Q���kM�.�W�7�k.�'�kĩt��ֹdw]��$���k4z�{�� ��g�?�;����[h��$�ݓ�3�B6Se�M�rE����za�������kӗ�G�Y��,���ߧxY�ܳ$�����J��^sl����K��թx�~-C)0�R���.����p1�d��le�����t�9:��ln�V3�g2�%��)Ȼ�?��Q�ꫝh�g��;�V�H+a�w�n����g.�X��k��<Ѯ;�V��ض���7���C�!��ώ�ݬy��ݦn�d��ݭ���]��>��� o�u�3�w~��!�I��_��_��e !p��W�q�I�wH����!w�XNe��~QPgr[) *�W��J$�]���緔��#��S๿\���k��a���
+�6�{*Z0&������.go�'����Yw���"*��
yv�紖n���K�ՕZ���%��d=躶�0ң8
<���b���G�%ŔG�Ф�����֧,�&���v�L�K��;(ݞV�NU�r�By����tPJ�2B�5U����jձ0oq�TK���;;[�M�2Yi3�N��K�JnGM��c�q�<�p�Y�Յ���_�<-v,au4�X���L�)?&�B�1�>6�ŀ�ei���Լ྄�W!��)��BW�?~ ����Qn|gO����ʛ<���|��(��[T�ؕy4?�dk���[�����&y��Ui���}~��W�c�e�}}V��u{�<�V�U�DE[��#B��C�/�9�<5�,:>}8'����1Y����������q���xK#�u6�Q��x���;�����!5���!r�"q�
g�����ñ�h\���(�ߵx�Y��#7�w�_��A��~�Gy�w���3!(혘!��!���o����s2M��n�#��m�l"v}���)Q����i+uc��҈����F�_�6���;r��^O��'�������l%@\49Hx�\������:x�L���E�ȟ������kOK��U��Rwc��[�U҉�RƊ$���-�UO?h<4�#�R��o`�Y�7�b�'��Э�ܙ���YO5�K"���IV�5��FtZ����OC��wz���b�)n����?�s."������M��WA�֩�)hsV*�	|vnCKskv
�06s���^V�C��āݧ�����=iz1�H&�y] P�?� ���"��E��!U��u[7��I�����7F��_̂�2���4-��T�m��}��#_u����(Cą[o��!�覕��f��q�_e�G�)m�O�@��(�����M��kBK�a2�J}�u&��~�<�+U�#���)Љ�)�o&k: �j�F����\h�e�w�ɡ�h�>W��I&���h$C��j=u�&��/�}�Þ���5/G#s���>��73{��|�Cޞ��X�[�b����b�7� h�����{i��C%TP9x5&�/q);�_��	�`���������wnǢ(���^�i�����ˋ�ݨy!�������'z�n�	�`-Rϛ�@���{�����F��X �<W�$dv�ĉ?&,3H�ǊI�򶰽����*�A~^f}l��j��\r��.ζQ4�/�>�G�Cq,�Nk#M�s\u�Dv���|&]���]�p�]�Ojѭ�Iw��4��y-�X�X�r�a"���ޣ;�V��S�q~�]�joOG����=@�3����)��x�^C��d�|�6���P�r�X����UU\_7=�M�l"�AR{y���(<���_X�P�"�T[Wwмk~Z���1�[_��▀���an'��(-]C$묤J?�V? ����Z�$*ǌ�{61� ���ȹ�`.��6��(uޱ���`�~�,�,��� �{�]��}�3@�mvO��Q쐳}nA�
Qx)�@^d6C.���X���y!8�����"��l�	@�oJK��d���Z/��ݎ�#{r�*���}B���bvC��ْ�9�w!.}(���Y����\�XYOb�y�
�p�HK��;mcZ*L��b��7${ӳ��9���V̋K�WK��+(2]1��I{������53S[����5 �M�������~��Pש�SE���FV��[G
b����78Cr�ϟx�[����$���5U?���+�`$�����.�{����Y���J�j�TM�K��?�mNH��+�����H��\1�{F���}=֕�s���״��몀�5��-1����ݞ@�놷��xJ��Ut�RQGޜ+����ed"+q�r���H�}��ע.W����nM�����v�ŠUp ��#�YAz�}FٜJҮ��q��8��B�c�P��Q�a1Nǋ^��?��ՙfX�M�d|���~��%ݱ�8j�fB��h�zK�����_K�De�w����2yJz��]�A
���K�0gt�YˑTzt��>S䵬P��rh�l�AX���W��[|�WP��?;%i��Y�'Ee��o|�zU]rE���c�X/�tB^_<"&�
��z�v)�%�D{PO���80�B#�N���� �}����5��Gj��gP��&(�`IW�s�����p���JH����i��$1��ĉ-L$d&٫*R�#�*�>��Rg�(�9���<���b@�a�`ͬ�6�r����S������8P����ڒ/�W�[v;�N�NIl��ͣ!��_^M�G�I�|���'����s�dd4}ZU�7!2�]q 5���Ģ+����?�ax�Т���[�����r�xi���d�JdL��>��
�
�ff0"�U�it�yh$�QW��񦈮�+H9r=Q� /g��AGk���9\|�~Mmq��+��p
�0��:ԣ��M�Ra�����e$,g�9V>�e〉Gccϑ
�՞�28�Z!�]�-V�F1�2�2i����ȦϚ=����%�����s�����ʇ�e6W��u	�Ta�@��MSLF�u�
�}��qa��c��d���k5i��{���:f҃�v3���[���}"~y����%o�0sOj�Lu���D)���v�?�r��N��Ѐд����7]�A��>��?�0�T^(�2��m�ec�{'ʇ�U���Oq����z����E��5}ũu��.!��x��ڋ^��� H�� ��T�/L '{)jc3��3���ݹ��>��8��u�-�Nޥ-AH�뢉Q<T�x|��0�~��S)�+�LU���i�
�u�ڿ�v�9���*+���њ�w��maUrmB��Wq��)(���p�ag�����?N��<Cz�5�ǤW���9��Ϙ�i<;(��@���Ż;��Oc�"u,�}/�����gX7K]>{��4Ro$���T�}VX2̾�5Jx��2N�=���o��Ь�'0$��6N�
�m$y=?d��5M��� �*IVzoEg{Qt LB��?��ۨ@=�D;Ir$�m��͘x����pvh�'�W��	t�m���nP4nOWc@�y�zˀ	����M��"��z�YW%K����)�VH� ���?����RvP,A= ڵte��*U�.$���.[b�}w�$I�9n���b�6R+]	�x�D�ޭ��ʣȷq[����W��c��褈�e%^.'�����$d""p"��u�Z��o�G�����H�@�U�i޿0��r�}6�\����~�|�$���^O$�#�F2y��vJ��7 h
���J	I<����q�:3��7���p����$��}���q$��\���<�ՌΧ{��[cp���S7BTM�~��l�8
��U$�!����8�g#о�'+�o.y��� `�P�`A�̷�`��r�_��S�6�d��'�*�岮�����"�A��Rb f*i"�����H�h�u�����Y�K*�O��[b�z^�g#���"3����lb�9�� uHs��Ĺ�0���8Q}e�V�R�~�jTij�=���+�}W�Ǟ�pѻ�����mTɌV���k��yv2��F�y݉.m�μ{�:�RB��VUY�q�����'-��q]�]�JB3����X���[���i&��}���^hɚ�'����JUx��`hra��������*7G�}�[G'p��V1������D�:��6#�����Ar�4/��11�	���C��4�?H+��i���)LqOM�o�=kK����z�Zl�n8U�ifgA!P>�`��)>W�����R�(Ʒ��$݊�[z�EOx�9'z5*�S6u�'_�����A%7�Ą���ti�V_���c�ݐ�xn�[�{��#�Sf�A�)��v�?�)87FVl.�\���DJB���g���.�̢�����=e����L����!� w���E�hT�a*dXl#	�m�zl���c�#3��8��w@���T\�����cC�H��x�a�3������DϞfW^�������v�P-/X4��7=�*�h,f(bΈ6�=�Z�'9r��Br�������C�H2�S1X���׃0�h�8�4-�<?�5�=yPm�?���o��=R���7"��+SKN(�ɇ&�U�����(��h{$�rg ��?U#�X��������u*t6�<�/C�
OvB3ea�P��ާ��}�0'=�A�8��!^hZ|$�R4��ޡ��4���0TMv�Ab��-�/m��?���PC��4~h�gqJi�T&���K��"G(m��Q$��aI��/��k�O� gj��0���(�I*e���-�B�]�!K������i�ׇ��G�����y1��c���4���#4���mh�W�Q%�
�»��' 6ߟ'o:��k��J}Y�+����� $���;N���ٟO���tE�O�E�5R?�2�ʶ�����(a^���9�Qs�<$���r{иd+�U��T�wH�bD���ƅ{f~�Č["׆��7�n˙Ϩ��r$J�@�1`�- p9�	{��A��n�yL�t���okQ���i���xGSZ���#�t�J�>�N"�GCɹ�UY����r�&����!�1�*v�}È��>o#��̙�t���R�@EXV�ׅN�]o�7��J�u�o_sL�ێXX�x`�fK��f^k�e �mŨo��i�:��o��~��Yɰ��H`͡�FKM�4$L���k��ޑ��:�����x�T�h�N,���.���"��?�ݏݹ2a[�ytM�������g���@���/�`V%��P)�tU]	�5у�,��<��O��d����:75G��[\-�a���P�jh���7��mI�mx��<��1k�A8s��>�Ң����!?�7U)T�AP�g&H�x��=���HkV}<�� ���� t�]Ʈ��;F~�Fɭ��52����"-<�l�(�������wr/�k���bޞ��&�ލ���~�ElrEo�L?�خ�B�H& @P%��F�D��q�j)x��B}R]*>Z��$B��!�sn��!N����f�RL��x�	f>��WG�r\�W�����=�Ʀ�J^���m~����pT6,Ꭴ����l)D �Ug�4�!q���r�_����FF��T��_�:;0U�`�]���x*
�n�/߅�9���t󏶝�	��>)� ��d}�c�~ �.X�9:�H7��"��n�o�G�P�@m�c��[퓓����=H5h�	�p��;]i��X���4��~�.Z�y�b��ұ1�񟵅�23ä��M	.�� �b����Cd�o���9�w �p�ٚ���ZJHjO���?`8fKE1X&�UCP��Ѻa��U`�ؿW�G���6���TbT�C��l}������d� ��.YI�-\	5M�A6�tZV'���.��*�H5
�6�0:�b�h��6B땇���j����	���-��G���u��G|� �=w�+�&�[�N7��
�m��0(���Ǩ�U��̫M
ՏN���,�ֽ���N�ٵ:o�=Y��2i�����+y�h��KĚL��]W�p)��Et��(P��0�t���S_m
v�w�'Ey����BfA�
� �׀��k�K4ܽܜ?�9A��$��uPs���K s9���C_�VLY�I����L��1Tχ�����õ�������]�U��F�Cc��0�|�.�Wr�w�|�����I)0�G�O��4�-1�N�w���x�MKOq����2a<K����G�fFAm�y2&�o\w)�����#J�����yb`*S��%�i���{����O�_��ؑz��G�W���x��*ς�����B��Y��o�1��w 3���#W�1�����G	������k��V��3���\�=� ���k�OL�{�����i^>���(���[_�.j���Ӓ(gF���c���~���C[�����u�x��^u��_��al;�$�_��Q��y	F�Wq���{�P-��L>Bti����?k��ڼ�F~i�e:�Va��e�|r"&ʗH�[j�\�_y�.�	�\��te�Yz�B��Pqu4�?ω��B�a;��)�y�:��`�)�&	CVaiV)�%�`�ĵ�\�B�;UMf��ԄX�h-��;�^Ρ����t̩�E��bZ��fMIWۗ}���r����ت��'&�t�S�10Q�x����>Ϫ��Blde�o9	�q}����Ԧ�F�Fa���R�! �.y�1�Z��P0�@�)i� E�I;���~rEC�k�(@R���1�سq�A��뫢��Z��/,��0
�-�P>�H��*��9�I_Pw��mL�*��2��P �U,��:$L4�8��c�	
�������am�A�ד�{��������`�C�9���k��G�]/�I��eB�#<�A�=	zvCp���Z�������*<Ѱ��{M�.Q`)��A�Z ��vw�����Ά�Z��Ħ��&�'��@Qe�d�IE�'ogCO,Yj�	�?�8a���L�&/�ݢ]��pm
Q�B~�����GP?r:���s�r�b`�p��Qp�ȼ ��Nmod9فU��k��}`3.���qp&�����=Ǯ5c��E�����WJ�A���5�BM7-uK���C���R�v���2�Q<2�AL��lyd�*K8�O)�� BG���؉�}�m��e	�M�Ne��A��H�tRІ~��y@wh��;�����,��r��lÀ������"��{,aFpv�U�[�ٵVbv��6���V�0d���mc�r�ʛ��('��%M�_�Π汊\�5a�G+b��%?���_f-�YRC���(�KCR"��I��+��4����m��^w�b�qx�Ӊ#Tlĩ�{$uQr���D�<w�Z������ �Tg%>�#7�<➃e� Ɔ�t�/�i�
�������3���/^)�����|G�w��*�L!���� e��W�^8�KPfh.<A����MS��u��y�r���	��Z��PG�U0���F����pF��P?>{l��#�t���h�_C�;X�o�l�İ�����Z���v�(��l�I���/�R���+ ����zI�8&c��@/ӂ�bpŏI��C8��	�\�M7#���9Jy�T p��E���n)r4��u�P�V��19���ÜZ=�q��w�.<{-�\ [C&i6��x�_ �I
'�����t� -7N-q+�+vf���ZC=���ևp^F����̠�ӝ�^RiYFJؼQ���p��	?��גE���^��[�L���Вl���F�wT�DA�c����+�#[�*��~������b0�0���ĸ�|�Y�Q�kO�t��i�q����a�BԐ�u��Ү:��#�W�n�ͽ�69��#SNd��& 
���J=�-�PqY�����B�v�O�����.~d�U����q~lX�#��c�D\&!Z���y�M~΁/T�F��0�e��@H7���qH��`�~�gD����z�'M�}��R��ٿY�;��y&�q
���������g�^�-�h�a�9�AhCtۜ����o������!}-�<�%��H_��)96uV�(�o�=����R'�4�.��=0�N5�A��pR�^ }�x�4����u������'*n�G{�|�"#B+T�%���T���T�r�[���A������^��bt��m�P��x^!�����wm�Z�_�|���p?6�D�{�5�1]�e�Xj��> �̿��������K2R��^��4�ibt5e�J�1��s^�Df��9ޟo�V�vf��S����'��B���A�W�ip�a��Q��	�����G�8�f^HI$�ԉa�0'P��t>��� �����T\8��˸�����AI��/m���cv�h�k0���{hdb����N$O
h��C���`Ӄn�gLe6څ�y]�,=�,���,l`	7�ݑ�"R����Zh�h�h����l�����{ʘp�U��H���Bi$_?h1��`��@�;�U��˷�?�>�[oLJ9D��l�ӏH��(��r�Y=�LI�g�Ё������p�5>�Ի��;/8j��Ñi�co"���$�HH��C��T��U��߄`p��p���{
ԕp��Y��E���L[P�ꞇ("T�`�ֈ9�_�˔�B����!�ku�I����A5"���b�2�\����mU��#���9~[+���k>}�Zf 1��n�Ǹ\��o���	V�t,��c�$���i��U���6C�!46pzR�V� (`A�(���i2s���r<����N(z�}|��쒪��"��xp��XOUT�B��N��� ��H�]cUş
�"LQ����v����9�L�A�Nj�4,��q�L�i9n�I���_���_�q�:���'$ 89܎_m��Ұ����\�Bq���L�j=���m��a�/ۨT~@�"7{Dc��cr�S�:��\k�|�lH~��w�0�(�p��N�02ݩ��y�=	�>s�tqW�9Y�l_b���$b{T����&����ϳ~]j��0h@��O{R|�Ο�̙�����7�NA�j�N?���]��JzW��������ə�Z.{՝ᑎ
Ơ�:��
T��J��W����G�m�&�[#��U��~,�bԕ���&��=Z��^W��B��[�2�O��r�~�!�"��E�_1&�)!��=�*_��w7<!��T��&h�@�~4�i#��d���D^���/��CVo�Ԃw.��N��#�-hr�u�4N`�n�p�(�QC՚����ad�����oa.��1��=�r�Z(���,�@{�W+��L�J�/.G*����V����5Q�N�����ь/h�91<e��u6�
��+��U��r������?3�(�,�,�6�4�2�@L��&Jgҳ6u2�K֤ڗ�da�Mu<�R�V�@Y��I����}��tM�����W�4(��=9m�����Ӏ��
D����ͯ�WI~M�[��t2�K�M[���|h;�3��S��;/��ֶj^4��	ml-��g_}�5�k`�����xٿ7;6�Kt�6ٸwF6*�\�N��Ġ��z�^	M2;b��6�Y���x�����=N}Nr��o�x6�O�\���/����t�����k��7�����ءc1B��A�G� /��ȥ��:�μ��%v�͇5���zǏZ�2M�}I�.:"ߤML����h��tc��AE��G�~��~�
	#a�4�X��']��L<ln�:�g��&��o뢝����Qv$x�T�R��pz��ք��́�(~� ]��2h*nX��Ը�=kn͞m;���
E����5��\��m���GL��Vˈ�ϲ'��:Df �Ƹe�i9x�2��T�@�k�-!�������Wp����0m����.��gPV����T��X�׎�x��s�B���`;�hg�T&W8�e�^<�8��lM��ޱ��<���4{A
�ד~$��W�L�lYae�Y@-�Q�kv+�w��,d��_a�аᣢW��vYw��J
@A�/3�s�%���3�M
cP~�H��9x���%�7a��d�������}��[�Ɂf��D��Z
r�QPD�����W���^<�|��y��k���fP����</�Q�w侻A��5�c�T�3�Jɟ�D�j�|�5~������ V)�bV�}Z�3����rB�����:<�[�>s�G6S�`u�h�(���x��J*�9��5:���_A�#��i_lT���=:@���\&���M��#}[4�ړ��do=��)�� ,fJ�UŌ�����E��ܛ�aQ��RRu��#D�jx��w]W�F�r������W�H��c}`O&�y0��z���4~�)�4
[��߸5U��2P~��u(MEx���w9��L�νH�����-=�s}�נ:2�9w�:�~��Y��D"�U��K�W��Kօi�h�eK������k�S��${����ǶΠ��p�,�'���-�ْ��t�!�3��׭S��Ӛq���亳���4��$k�8�}m�����l�Y#R0#���7B�Վ��e�����9������c�;��1�w����#)2hʭ��m����=�?)C��+RaEp.�z����[���GZ8d�eP�@ګ;.K�6HFI���)��Uz���.�F�80�L4��}PE����J�xL9q�V1�z|VǆT�?`	�	S�f�Q~���C���u�3*D�1��q�~�>ə>�D6Z�=���X��9Л��Z��'lI��OPj��	�������u�����1�x�=�P���A!n҇��6��q���к�qX��e�kQ{�1Z��M4^� h�[GHݦ�J(�
>M�ȯ���8������� '�Q�U�Gphu�؈��[���.�H�h���X�/=|�ò�)�ZZ��?�U���Ǧ��� ��ޞ���6��k��7�հ���������v�eYQ�ʛ(�E �?��6�ɏ���$sp)�R	�;�B�U����vf�$_I��fy��������D��b5r��*hQ�N
���U�: �����7�߃b'@���Vr���q��9�Jz	&� T�PL?J��d��f!ۊ�S��p�,{�,'�6�:�U�q\������Q}�����{D<Q�h�ՠ��Ȅ���\���r���Zs��5�N��\�(����?.!��چL���@l�_ρI��:������x9IKǕ��Zb�V�d�ڏ����q���?̂#��x�4��-���`ɐYZ�o��U�R�r�(�-�"���Zt^e���o��.�)?E�@�i�P���O%{gAv������HW*mg�S�8���Ws�u׷HA�T`�{g�����m9*UX3��	m��rߵN��녡����kż�ܺ��[2|��l�����3�,8f|�x��>Uu��52[�2�Oe�R�m�ב�aM����i`��3e���ݜ7AB� ���x�����孉BQ��0�
Dl����3��OE�XX��V3/�,W���˫A@����h��D<�x�n�r��M�2�t�pgT:�g���{j�j��J7�<� DY��x?/�����v�����B�f�Q�F����]�-�<|����Ί�U�];��y��;�)��t��03�k�^}��Hd�	�l?)���K��hB  �u��~ts������G���V����ͪ%q�e-,�� ��b�l���5D��$3��rj'���:�����Z���G˚�g��\�-l��N��?��d��I��dC@}���a&��?k I52�-`۵6��u�:�?�+�Ezl��0ĕ��\��<F=���r%�f��H��&�?-�b�H`��؃��r�:`�j����h���F��D�������2�2R�A%�!�֚3S���nhB_I?~�i荔��\�z���ȴET��t���7>z�;<V���L�u4�w�J2G4.�?k�*)�pn����m\��'I�����a��Z��Q�f��T����%H4Ş��C�k-\�@�:y4ux�\w0��9�������[T�騭�{TH�����6�?1Mt��h��X�U�Rv����o�s��4j�j�:���}��0��w�~�EKj���n�R޲�`��� �Ls���ү��ɻ#�h2I�g�ma�*Ơ]nZ��y��hQ�f�&F�kh���]=S��8�2�3V�"�p�ܡE7��7X[ޮI� ������k��F�W��qv�N��ݮ�IP�V�n�#�b��/�c�I�B��Y�J�gN��O>�å��%K-״�J[/��JQ{����<L�G��0�j7�:�k�<�X�ipzS�����n����Xcp�|O)����P�;�`�rw@�c�"lq�]�0ɠl�Բ��HK��UT�f�0=vQ�n��##\�N�6y�O-q�	@���Ps�]��� M��v]�����XZ�*����W38d��o���k��񙜶)��{F,�}E@�h��o�s�G����0��G��:$��ː'�l���1�@�?,��ƾ����f�����W��A�@'�/�m�żmؗ�r��ʓʱ�M�&\�E�z}��mAX7�ً|�&1Ize�$2<j���N�=Y�3�k�#��e `6���v��?�9��¬�䂪�����{ߟk�ٕ����[R�Y��E�����e�21(iu�לox�\<��e�2'?��Ks����y���/�9�ga��j�r睘���%m�w���|���y��^pz���J8;��%�x��*0����.�+�
��P6����q`�����R���CԺ,�'���2���ϱ�?/�ΫK$�1��aσ�b�uY�`�%x��b/�n�>�B����¡����Q�eS-D���l�l��L�-�2�jc�4�����4�m#��'y�b����&�0 _<�Qg�~����Dƴe�,�F�%Aȹ2�0�n��E(G�p���]z�y/�  k��Y�}�k��/Hx���]��ky�:x2��)b��Μqy��E��5�M�n�$��ZC�xg%�������C�Sq�h�.FKH]F���~�2!@��r{\*����R��u��_0t�%\צ	�"�]Nw9�:VNw��ls�\Xr5ѭ�U{�i����t��̶�!n|�6�[<˥c� ��a7��"��H)9N�+�qx�BF���냙�BS}	q����/���Qx��p>xI��`ȆA��̩E�<]+8 ǱQ�v�Y����4�2�oK����'����\ڶ--�O�`$.�4|��ՅyaSsZ/���Y�GHW��oW��m���l�����|	Os�禤E�X��4�:v���X%V�آA,�P.�&���u�f�K2�J}Y������'NA�E�`��y��"D6���,��Ά�;����<9AU,%H%�v��H�[�W[�iD��L�a�z�ʿ��["jDgt�7-u��!���`���h��/7ZN遨o��;MM�Qܭ䅝#����O�R[[i�v��`�%U
q���:˰ݯ�a�!���+��I)�%�e�Q�%QU�ޤ��NlP����-�s�3��s���)?�I%��@c�|�x�F�Ga�-��|1a�̌K��"�
v���s�%�ؕ4���Ʊ��RD��2H;��`,5�� �|ðDY��_�_
G��4ϋx���������]2���T<?LIp��3��~O�%�c�r���!�?T^�Jk<��=��!i��Ǜܪ�J�O�6�,v���:`�*<!��:{��rȃ�$	���~@�"�Bԛ�y$��fO&ETT5-�BD�;��W8D�^�����A�f����M6x�)�ڠ�dA�]?�g���'a���+{;�]Ӛ}[`بZ}ki"k8�l`M��r�\^!�������C�r�{��E~I��Z�څ^�;i��)�dڇ,}�����!��P�O���ά�~$`Z�r�^�=:x��K���eO��J�֙��(�7M5TXz��RB/��H[,�f��[Ǆ�;}|�$���raUxL������XT�����'�,��!�+�<�;�����I۱-��X�N�Q�}�C|Q��n�*lT,s+�"3��F������}�YS��DuW�[�/t�/��Z簙�O�(6�z� 79X����^ώL����"
�dt��9�fd�8�x����@��<��PK	3��j-+(�K\�"S���A�*"��YX�����F�VG+�{�c�$,�V���U�u�,"���a)oP����c���W�^���ğM��� �*��z�[V�2B�}da��̜�	��X�}�M"��f"��à��>��e��ZY0�������ɺ3��d\M%�������G�l�0�m��-p�*Q=����6ǋ!Y�E�Jr_{F d��ʈ�K؞��F�,�&��/u�C�h2��H֥�U�m�JYz��Ns���S���O9H��zz�n�+�x`��M�ӂ�]RMs�>VF��X҂%��-��(�p|�&�#W�mɟsAo��i��J5�Q�Q�D-���H�Tn����Ҧc��3.���|vD�f�\�=�z�<���6�炅���\@Nr��p�����^��I1��@�E���� ��s!K���#I�5�FɿY�tw���u�jr��))���{���v�f#�a�w�r�F{M�Bf���U�A{>c������(���K5Z�IQ;}ܧu�q�½����%1���I�|4�p�!��Z��[[xh�P�3P��`h]������hu�S��ކ�@A�\(\9X��ۖ�	/ʴ��������u���F1�[���I���8x 3b�,5\�w���g��`��n�g�7�mƗ�[��ڣ�^p�)�\=y���gF�%�TԜD�@$o��㤼N���p���ECIެ��@�p�ĸUWhI���|��WQ��f\�? c\^y�^�mM�<���H�݀>���D<���כ}O���r��0̧�����ۀTH�/��!��x\�G۰�Y���W)��#{T��^jVBY#c;����l��O��~��ŝ�G���uZD1��?���o�7��W]�C����\/��@�yU���s�H�C��� QH.��S|N�֮�V�k���ApS0o�F,%��љ�@t�l���`�r�b��A������/!Krɝ��K��;��A��%�������ª������,�%zK����""Ⱦ������p�����C��A��^�^^'���PF
qoC�_�RMm�7�4�s�d�eEJu.�B���3��^j=���ni��a�S�
+P)>�����1kӜ�����}[�������r�	�ϖ{�XTN!0DMo6���w�S��An��c@vB�Ǯ�����Ο��䤦��A�n0	��5��Ct��]Y-^����%rh��4���H�߄KaC�2�4�� �=�����V/V�	���)�0�1d@Ы}c�n��Y�~�:�a��]Q2�0�S����|T�U�>�	���(����/�!$z��}`c�9�x?48Y��O�#�I���w�(-�DOҥ�ZC_E7�g>���%��^]�C��c"^��vy��8�R �4������p�Z/@�v��jn|	F$	/�6�)P�� ӹ�˿�Н1�s[�} 	��?���I�����̂u=��Ii������E��GR�&Nh*��_��+_��a"wz��T�O�8��b�V��a<�"��;0���W�h��mtmj[�g��[�Xgt�~�waߐ/��6F�=W�ˮ�z~+P��S�T|9#U����6����)/�6�G����^�����!i4��i�-����J4	w�挨�`��Ţx�a�#��I��6�_�	��=P�����ح�>w�d���Mp�1�Ղնdj7c!d%0����8*�#�W'�y��;[t=�8D���{�Ш�X�5w��������P�1�����m��p5�丯�����mv�tJ%�,��&\w�p �,K�spΝ�;�Z���
vL*)��?�LF����҉S+L���	%�/S�2���/���U ��a
�;��wN��|)�PϋF�<�3?��7F�ω�2�9䘒���~�iL�17�,,�+
�赓s���u)WO�c�'�}|�)��L+��<V�a��wX��V�������i��P@��)0����zGi��=�:��E&e���:V��B�F�/�Īz�i�ƵsQ�q��Ue\�~�Dh�X�l��琈�VGl�/�ާ�
<C����R��l����h���$M�"���lw1�y�PHHrP��rK�P��\W�ohv�o�"@��B������������?��2���[k�9���>?%F��X"~�-��M����oT�m���|\?�#��ػw�a�-�|��y�'���S/��x̔��޿\���)�7G�1w�ޯ4Z�*��4V]�MXS�6� u4�߹P-�� !W�l�f�<,��C�@����=��P�8��Mil'�_��Ng�$yH;�v+CN������N�F�h������aH}�&O��<����}hZ>�XpKz������\f���d�Th�$R��_o,qdX`Dl��$�y �<���05|�6ҠE��`vB����:)�)Z���	�F��Ih0��_j�v�"��d��6!���<
�z}�3���
�Q�( #�MAD��\���h�Ҋ�>*�Ƕ��N�`�<�=���N$��mpεp'e�kT�^������\��H�P		j���GPgҠ�Q���JXL��o��s�]8-|�3 7v���\?_)ã~�=ںfΞ��Z����kN�~+N�8�Cx�j�CO����K8�\�Ѩ/Hs{��T&�0�������^�n#C���S��5hp�s!��uR!�KR�#b|(�C�p�£�?s����b��w鈥&d��e����9\��RH�䤍^���j�ߜ�~�fY�[���M��M�h�SW�P��Va�9X���RX;H4�4��m�r>�W`G�[F�J*ȁ��hk��Hn8�1%|Y1�l����:O�1��
`NX���>��ۻ��S�¾�m+�yPV
���
_�K����e���]`j Y�q�)��?��a�Z������6{~��q��Z�8J
t+�m��6�Q��[6I�G4-���])�\*r����.p�$ ��� ķ��N���T ז�R����[��V+Ͻ��g]��y�wG�NZ7y+tX��#j�Aho�8��z�?������U�o0F�=��m��A�n0�&�`��y�B� /x� �,��̳Ķ����%rRbh'�H�&���Og��T��䶖DAC̸cކ.Gŏ��y&�_I�ϟ��m_�������y �������͂;���=į5���c60�`耵�Nf$0�#r���y��X�ƚ�$Nz;����dS��eh��|Y�"�J<��s���E��4|�!�<�<�2�X��Zۦ��PL��v<䬢	�x�r�6�z	�I�KW��[�3��k
��c���_9)~7����#b�9��KM	��������p6w��]hAMg��k��.كۣ���6k���$�bEԿ���}/����	���oM��v�c���HB���g�3�`��z+^ pL���*�X�(�l�\(27����-D{j%J�q@����]u���
����ڭ}M�y4�R�"��<C�a���TgP���W��g4�#	mҩ����e%P���	�����t:��|)�����Y�*}�kl��n�[sU������u��Klf����[iA�%r,��
(I&hE��ƲzTl���e\��{�q�8�c-�F���^��%Q�m٫�|fc�(�I�ĳ�̓:��82��NIj�#Ǣ��7H��-p[���=]̓-��7UD�����}�	���)����ix�ɷA{iݰ�)�86���h����@R3�=���!�i�MGeZ�̄C�I�_D��-��
g�$�!ঢ��'�!���ݡ���x�3� &������Zn�1��O��(
���k��������|�*_��%KZx��Wi�CI�@�ۻ.+��
���*2�!*m�=�ʾ�f� �Nf�����DY�N�1M�Ѯ��c�s@'F�F��Lޕ�O6���P�S�[F�{�ɵ9�DJ#��Y�86�7�� ��b��$�G�={;ȍ䳧Ӣ��9�Ԋ�A���oS׹RU�b�U18$wp\�G����0N��N35X��TQI*�=��~o������Vd��_:� �;W�5�Ek"/�G�NJ�V`Zi���!oY�Gx��"��<��Zgh�e�1"�V��f+�1�ͽ�t�e`Wð�o��!�6(=��a���`�V�B�?_fpō��e%�(���s�9���Ď|�+.o2'&���Kϔl�x��ޡ���`6ӄ4a���P���_m�;m����`���vwp�oB�##Mݑ�А��L>�`w�e�ej_6����6|��b�Dk�t�^';֤pC!�i�*q��a����X8�7�T�����l����W�H��(�H	W6�q���[05�n0�R�^�9kk�!!���髊���Z�Ɉ�iR|��BS1�t_���o�����WB����g�>d��u�p�S��%Q���:����*��R^�� ���d����l�E�[��XH�wI3j�<�lN�T����]�h��4}��Qj����P
>�|�,�{��KOU��bHX�*�,W��#�
�N�_͠�7�ĵ�y�v�{����<�.M�H��[9�i�'S���杻��9A��dפ(�Dh�.���7���j�+Qk
�M@*�{���dƨu���cԂ����{7@f8`ݱ^A:�_���%�㴽]�E.
p�~���n��k��E� 4*ގ��H�j&u�����$����H���xK���w�O�%̀@���6G��i0Y��f�W��rt8;L� ��b�b�M_�`��(w��?wo�ƌ�F6T��q�@Vfb����	�D�
ScF�g���_6��JVM����`�D��+���ix�Ɓ�	X2���˃�8#�E]_�S�X��{�{�t��'���A)3�4�#���x#��L���s0xr�M)֍K�n��g^�of/+�Ky�A��x���d˞\�b��.�����D�}��^y:��k����6*j*τ���L[���M��O��4L����G�p=w��y�?�������Mz(��L&�v�d�u�2�v��K����16�"9g�H�ݧ�( 4�}�"s��M��������E��L%q��<��߅���#���y�`K="v�d�����ѡ�DB���?��""��t����NZR�^�����o��%ޘye胵���}�K'�Ћ0�k���|9�5�E�e8:����Bކ⺋�P���A�-�g2���R�$��a�Ћ���K!RK���/�����y��e�C��$�BH&��"yOR���$���8�X�ʖ�r��;�3�@x�CO �m���)��;9���o6��w`�6N�^1���ӆ�s�$��b_ ����;�B%~~d%|��a�ؤ2FJ�1�.d"y��69߼�UҺ��������NP�`81~�yr`���L����Z���6lu��p׵��9YV�,��|�eNK��OIfd����9bpk��`�גM�)�TV=vr��2��s�A?��@l\3�،Y�M�<4>n������1v�B��Zb��+�@��6�C�t����&��J�Q!WP�d�5�p��wVW�����Q�7^�v���|�r�m�=�R��v���'�L�|�~��-(��o���ȣ�%�}��� ���[��x8^!��#<����&��y��r`~�ۻ߾��62�qM�NNd c�9�,}Wq��[���	A����MDpW
1�	G*di#�_�)z�͉p���/`6�q#�@	*?��0c���~P���Q�5���6�7�"E�m-�eg�{q7��;�V!�E�h،��|T�� ���g���Ś��� �.r֐L��)�[��+��?��p4��c����.tTA���%g]�]�|�K-`�r�]/��5��3a��u_���R+ږŇO��2,���h7�ʓJS�F$(�A(����6]��n�k�~5&�Ќ%l|���Z��>�%��Cj�j�Y���H����J� �~l��P����N����pF�yڍD�����y�~�0�ϐ�`�o��c�!�u\09H3Q�l�ӯ�����ś��Y4��z���i�D�X�����(�(�N+w6�N^�am�F$�w����{�T.�d�/��扣i~��{υ zY4�͎�I��[��ѯb�l�'sDr&�\e�]$piB�0룱����7޴��$KG0��P7p"۰��o~��j9=ت�0(����}�1|&��t�����A�NC�r�����0%r��N��K6e�&tu�?�s�Wֺ�H�����,s:Xm��.*��G݉�hv� �_?`ށ$��K;��.�>�ū9�,��̔�#���ӻa���Y�7��ّ=��RFū��@�d�|h6J�f>��%�-F��9�Rhٱ��ם_:P�s�H�U�Gp���IC�ͫ~h}�5ϰ9�l�j\	�[p�B�.�{�ڧa����Ab%l��h�g���k�Y���ָBWR�����1�Q��E#={�=K����e�_;�>Z�_���</Fc�c����v)��_��}b��yd��Ç/��\o{�쾎��Î����I<l�ھI��&g�Zȣr����ص��B����GA<{k��Ȭ��j��V��(m��s:��|�%2Y6��w=��o]ޚ8Z������֒�P�1H/`�<�p� ۗ��R=��cDD��PD�#�g�.�,j���myѓb��5�z�ʲ�%8'�����e3�ksi�����1�3jAkF��V_D�uJ	ē!дXux��B��=!��|�
�Q��Q�HϨ0�
E[�mY��E�KU�c�������rRN���Ѥ���F�,M��n\���}H�|��^�"'gI ]YY��f!��� �X��ZH�$6װz�M(�M�Ļ��9� �%@��7T�Eh�A2p%�Z�V[����n�N��'-��U�_�\�L���2�Og\��z���|t�$�o#�}�*}#��l��K�N�C�k��=\��׿o�l�r�I�Kg�j�(X�L��C�c�ߢ^�*py>�F-����jS�?zE��"a4�J ��(�;�Umr�nH��Йj3������ϾJ�+����yCg�i"�;���E�(�96�cS�$��N�cc�EP`�|� }�<U��Ȫ��5����M<,QT��V-�g�O�}�����`�)܀��/��ÿ�-s�%�;��ù�I�;�X�����D(�N���e��)��8:s"�\[2sKg���5��`z2�uD��O%j��N!]�QR$�/�"|rJn9t.͕��-�]�B c!ϛ�F�C&�H�v�$,�~����h;�*E�j���CM��T��^5�UB�T}�?{o*�c�[����une(�0���;��֚�[oer�mMe�>��x�4��?O�E�(c��b6O�4�_�i�h��8�D���"[T&���Pgk4�D-7h��K���f)v%�T>�����9HG�?ϯ���Ac=��&��_��|�0����^�V��6£;J�G6ytȧ�}F#jV��9����ndE�����<����q�b�U��]�(�R�.�h�-�vɢA�h�fe���x��a�q:�����L�%�V�w�����Ч��}C�
v��]�ې9�d��/����;�Y'�_.0�`�?-Ϯes�V���)�Yע_�]���xe��{����r�S��`��~T�Cɂ�����ۃ@N���������/Ǣ׀u&a�"�iS���`J-�K�l8�&=��qH#�J;�!*��=7X��P����7�Վ�����z{���T�sS?|O�	��^*�ra�����^��$�W���g�N���g��v�+z��ط'���N�Q
4� ɧ��[/-��o����a���Yv�2��h�ù��W���̤:��]���P�ǖ�@��>Q���
��|s�=&�����!�m93~(���2_�1���ÍR�_�q I}q��s�ϱM]!�窥�f���́o�<��k�����w&�sH���Ev�Ff��~T�0�5qr'�L=����!��ާ�Ќ��負���dꄓP3]�� 5�E'�>[�>/�]�);�v��Pl�^>�! ʛ!����F�'����� �}�QԎx�k�LGK^�n��� �N�#ox��J��I5z��<����W5m�*������eqg~���8��}��I�lX��{��r&�L�Y���F�s�D��ĴOx#��@�"��j��� I=��[O>7Q����ʛ듫���ޡT��m�2o9�!�J�k~+np�0
��LI%fBo�
�Fi`�i���
i��O�Ϭ��9 �p�N���� /�%�k{�㣨��V6��_`�;&���ZO;�,I��l6�Қ�N]n׀֦չ��R}�E������G��5�a!S�?ep�󯘗&�+]+����|~�{$�%L�K3�J�wb�o��O��6:c*Ҳ��KX���j*��X�߇U#�!�����J�"�]��gh�٩��y�(�f*B���t:�b�R@�����P��%�0�S�"�S��[���$?uq��YwXrLM|Xb�pC��
�cj 1���p�~�@���5]�*��[��jyrπ��x�i͞�d��y'^m�=��� S���{F�^�"�}���W"f;���y���KЍ��лa��^4�Y	)�`-�y9�55�愃�H��
���s�Q�p'�{�";�;~�g�k�@S8e!A��}Q��_Q(��C��䀙.B�;?R�ƀ�W��Ad�bf��(�Qr�<5g����u'����r�ȧ����Ɇ�u�:��7
?��>xE�����+f��r��_>Fb�iX&?l\ǘ2�_L�g��	v�h��1���ـa4TD��\�*��zeL��Z����FTz���<�Z2�U�!/D6����^EI�f2L��c3zA�:���R�N�?)���)&����95B#�m�;�HM� �Q;�U��Y���bl2p�в���8�t:!@�PL@�d�<0�,!O6�����8H�M�������Sظ��?ӠO�~�����{T��@Q������_h>>K?�[�t΢��C��� �s�qhw����_w`9G:�s+�p�K��u���u���%ϼhşSVM�_�P�Q��G2S�] }&ɉ���!>"t
����?�e[+���'"D����[��E	B���`����z�|�F��}h�7�*ڨ�}i8
��Q��:fe'���6�d�����&����{<Pk~����v�\"g���HT�8\�!ݞ'V�����^������l5�#T�3�t��#Y��ct$���	����g3����Deϸ6DK�=�V ��	AgI*vA��
��m��ￒ���R�¬h����,����˓/����!�ńF.����ǯ�3�)�]��r�r��P�~H�T~p�+��IY �۰��oD��f�iT���xj�T�'`q�,n(-)��x�s��PcS��$���8�I���v�����
/��"!C�1��YMktÙ[Qg�M��4��ꡩ՚�R�Z;n	��������-%m_9�s��S��̗]! [���%��n�v�^t�[tݞ'�n�����E�n'&��r(�����bO� �_��(	dN�+������M=X1u�2�[�p�<vA�����v����]�����>��@�)E&eg�V��yX�Rn�LPc��͖�`u&s}����Dҿ3|��	̜�J�̖à@ 0�!�C���N��x'�+H���������[�գe�в�BH�� ����F��WZ���A�C�pj1��2�M4$��%��x�<�5ߺ��}��E[a)j��
�6׷c�5SI��.Տ3R�����~Ҟ��#����^��B}C���$��y����D��i�0�OZ���w2���{��ܗ��~��km��Vr�Qsl���+L��n�%S���w��ps��C��X0SG�4�D�����|"�Wua�i�9[�^����	��U�M�_g-k,���E����U9�AU��$��
T��p�$]���6(ө�bA�\F�J�vT��%���V�GOF��������n�W����)8�U��B<3[�FOm7W�#��[?�Ch�߬]��)}��I]5_UY���f�>�@fs�w����|�ca����}[A��-?*���j#XC̼Uu�}�~�V�j�w��~/}���"�Փ$A&��	�:w�-��h�����I�E?�rWV5�2�F��@;�B*P�}�1>hou�U�k<�qj��x�b&R�:�<9O�h��Ws�������yi�Q�4ȯ13V$�ʮ���qs'�^}�m�P��v�:���w[����R�]W'��1�E54ma��g|����m�_i��l�F�gJi*��ϖ�d�f�&	���j��x����|Z�_�rul�ى#u=Q^��h�)8��eҙ��eB�������[�c�g���SI��	�Q���6�ƴ�{j&�l��	C��mݡFMl�HPI�/����\?LM'8�:�=PA"��%�\K+�U�E���2���gi���Zh����N�m��k0'1-vC@!ɠ@���W�m��&v�!�����伖��o�.��.�N�!�I����a鱓�")���jFLP�Y���ױ����o��� �G�ϴ5"B&�� ]�S����pwj����Ͷ���� ��&��ŗ���R�����?��e�sZ�h�f6���E�cT�V�ML˦,��.L\��|���HBG����n�Ɉ3��k��L&�-n�Ȼs���1:�{]��o���#�>����]�\]0Xȉ�^�9,��X��%*�[|lT��bP�����K?�� ]�-$�Ԡ�՘�=�dw��`���R��U^���[c�<*��t�O���ǲɚS�N>�������Ī�elJ�] 6@1���Z��I����8�`��O7�2����� T�1�����zl�@G���Ld�d���,�u�x:i2H��%�+F�p�K��]�%��MZ�Z����^�~���E�\cz~�g�NQ���駄�I��X����pH���1�e��w�J9\I^��$Pb?M���y�? G��,_�#�$Ӷ�k�ݔ"���(��$fe, ���Y��\��:]<��D$Du�����O�����>Y{M
e�jS̓Ɵ�p�`I�&xD<(W�"�2fYM��������?���'�L���4���Ô�ې�cQHqF:��6�Ԅ�(ԞB�&������=�J������bL1V7;<\�&�\�VM�v#����_�M�a�Os�j644�$�#�&���p�b�h�71^�%�E>@#���j�-���3�=;KH��9�0�'�4r��j��)��P�d�T_M��D�8�^`�<p���ʙ��y�-,���L��,c.O�%�O���8v/
����cBQq�Z4�;�8��I�eդʀ�M�ɐl5+����D�*���n�i��;2���_I�!�zO��y�|�H�8î)z+�ť���L6 ߠNǭ�F,�v<�K C�~�i����G"؟C^GY�#�Dy�r��%���Q�O�Q����P��<(m�w(���ª/����q� !��ξ�3�7�5����j重���abH	3���7'��
��{�2��5-i3����/45¥��vA]ګ����{�U6+.i��m���5��K)�)� �*�����H��9���ǽd3��	#�����������QȔ:��S�w� ��*�m$�j`��l$6g�7�� ��:��*��%��B��������s�%(�	��e���U��n��N7�ہ��m�U~��^5E��1y��T�:�������H{	�ѵ+�����?��8�CU�>yc��D�1G��iT�$~��eg��5�����މn�sbc|��+7D1���Rh�`�%�o��YtS;w�����p{�rZp��p~)XA�����ZY�jBp�t���"�^cQ�T�(�d��>��=Nf9��q�����~�Op��Z܀�j���X�u��qG�y�c��pT"�fzނP ��F�S��WB/h��a�1�	Y���&W�&Q�-�Z�}HDpr���'� �\�^m�SC7��aW31�����[���\���E&{]ZU��3m-m7��ԗ?��`�;�V���%�2":�&�]�~~���2���/��3oWs�OԱB�g�T��^,�aDѻǍ��t�5G�����p!0�Jgׄ�75���A:"��8��}�:�͋��8�?1{����05@6_�YK�ۦ�K�i��`o޿б�^ͺ? ��qM��[J�q=#Sr�X\�^�up0i,�Ս�_��Gݸ���9���qŖ<�E�}�p�@���V�&���A�8?��WH�t�M��9�^"�v5�yt�~���?�T�ٟ�=�._�����F�dU2�aD��푬Ja��p�<�Ќ��@��l�h@�N7�0���w�����.\Š8؟���@���u޺g��C���#�@� U�-4�d�d�d|�2�λ�>-������S8�^je�|nL����c��<w��=e��פ�����e�q�[ ~�G�]X`���>P ���/³���<,P?�fT�P'�И������,P~S��W#���M[�R/�1��K��]�8��p@uʃ`�Ӡn;�3��c���Yr�Mb��4�X8٪�ʹN� �� PǻA>�c��&����g@y��#g�vÀ!���3�׆�$l[�5p�h'�F ۠l̿���-� ca���m1�j2P)A��#hGb��9 ��5���g'(�CY��I�O��舥SC*���N흙�xV0���?�jh����i��LC,�j�i�j����Ëc=< �j�WI���˂'=�U��>O�;$��~���PW3�w͔���G���L}����;�b�o�`_/�'R?��9�A��/P�D���e�+0�s8�F�>S��*�5G��qR���S��m���Yw�'U�3c��aNos��4l���P5~�kS=S�j�;_'�u*��}.WTBn�m:d��=����}�kG����4(����I�-Z'� l2Z=����՞F�Q���N�#��[���?���m�� �Զ�"�� H���:�X����MYx>Gn��S8GA��"�݈�Y�n�Es`��@��Ě{b�f;(R~@"�Ni�Ю
2����0L,�t�G���2�֢d�zvl�ip5+�W��)?rU�i�N�M�[��	|A.K��i���qj�������Ӭ�����(u�ɤ�
�6}4L��R�'^Z�XV�U��/j`7��	w��*]�{��?V
�;gF����o�A��jf�v������0��te�iՄXc�0�&�`ؚBdz���ߺ]�5_�VQo��&�rPX^��k��K`�_���s��eS��E}��W���@�ι��2���R�61*X�P�E�%:UuF�RI�g �zn�\b�2� �V�U2ϩ���J ����;�cT ���@�G���s�J��-^Y
�ɟ�ZV���Qfr�um��e9��Ak˕����}�bk���U2�i��/W}�8f.gU>�ɯ�Ѵ���dwcҹ˼�VV���(�/knhR��7�V�����!��txŏ� ?�Ζ��t/�:i�HAן%�[A���>�!��9�^��m�.*k�落#ɔ�]��gW���&��5 j��*�2 � ��AȡP���)�����֤հ����Q��M��_M�	$'ܸ-];h���_%��I��Z���JO}	c�?u�86$`qp��/g��PƜZL�q1��e�Hl��0S4�ĶQ/j ��dvsF����}��$)�-�i�^�û#�T��!�b����y[��ѕ�s�J��kK����0�$��$�qk'��-�-�X��.G�+*�d�uɆ�?%͉֨q,qsͥp��څ�o��F>�m]Ffiu���8 �aFH.a���W>�xb�{9/�ޟ1��C�@�:~��k�'����Y����t}%s�&���h����'߮�8Re��u�dR{0b������d^	��ճ��@z�(�hh%�99u,�?k��叚_s�Z���� Ś$�(�7� T�ns��ae�H�;
i�4�"�k��῀���ETB��4_���^鏱g!���'�߭���g�Ʉ�����u��B�=�'!�Ϭ�Og�:o�x�4ӧ샢��q��Γ��͘9 >�xp���f�8�B�_"�J������+	�,hj� ����y��qk�������^��5]3
w�6�9�T�!���?~�1o�K?��T�m�V��Pq;�d~NՖ����r�M���n~S �0�K�?;�ɽ��t� 3�X��u��y��Ň�ɵ�]O5<��T�~�0ag�4WNF"�|�p��m�Ql{2�W�r�6H ��e4}�ʩB�2ìI��Y�L�t$��:pm�����s�ѓWN_ $w�R��t�Հ�Τn���-�=�=&h�L&�Mk�)	O5�U4Uz�qL:��--�<܃��e� ��ԀR�!^}��OD��qZ*h�_N_q��or�/��h�g���Պ�6	u����Y�LRړ��o�kH�q�ћj-��3u��L˴���{Hd���f��Y[O�	<h��㣄��(��Ş�E�+���hLI�3��NW_�H{dA��u�;aU1��&ͻ�߄�(B�*;��åw��W
�Y��G���
\m�#|�ٞ^��?ą_��6q%Ž���d��A�ѩq��~��M��V;�����A	=b��K�=b=ӿֱ�eQ�f�ǫK;���S|�opƗ�.��Ci�`�l�/59�h}�j��7��9D��x��f����J0[��v���ÜM7R|r�H��ެ��ؖ�`֑$�/�E���2��yC��
�����5�#���f�6Î�S�hI&'=�����I&�V�����*:�\hZ��)ŧ�k�N�x�������$"��)|^��@(y������|T$=�D�m��*��*������A��r����*&?쵁�2F� ���ܿ 価|e�2�?£=?�����U�v�W�
���I�?�r�uQ��<�t�$���i��7��ccr
*����S���%���Z�+��hA�a�I�3�D�%Ir��Cg�o�2�P��gm��nK�����8`����%��d׿[��,zB�
�O�^"�C%A�19��g�k�C,ˁq�N���p7��X3��垑&%v	i���Sa�w�w�yӪu���'�%���1�zO�?
���'J9 �>�H�r��'���V�"4��<���A �Z�}xiի^���'[i-��1x����;9��}EK��������D������"9"9�`l+��+��ө�'��;>�<ar��f� ������ޫ��Xg�7uO�4�ɔ!b�F[��3�5�eHF���#�`LEΙꂔ��~���dn0�JKzI6Bɳ� ������謜y��A�b�ʢ�ZJH�CL��Q�@�D��Õ0	f7���
S,����\���j%��iބ&�nM4��|�~nMU�G\u����=	�b�]�]t�������b�A����0L����,C�<�Y� �PtS��ul���E���e�d���l��NO�C�"��ʚ��>��~3ZjgZ�<έs����7S�< i���vʂ��~�=��ax9��`v�����)1&4k������%���ⶾ}|iE���3�����@L%3�ub̓v�d���d9���7bO���_��3��e]���JH)��F+�^Tc�ƿa�ɨ���2h�Q7��V0ݥ��[�aB��Ɖ�����'�W�,^��z$Psg~�l��N��|�\��R���7��0R�O� ��iD��0l���.KXd� �����:iݫ��¿��F�"bc5\\�?f�b�Ӻ.�|�.a���}6Y��Xu��#|n�'�L�V&�ms�# [<Y�����v����D�5
��MG���դ��^ӞAr}n���.U�:E�e��<*(� �s={ZJb�_d�
��%�6c���A<�KA�#ZїT&��8k9>�I�/L�W��g����'Xʆ�1�5�>�?�&01PZ���3�1=�L�^��`cC��KB�#f�:m/,��p��%&���K+Ƒ&���	���=�U'�#ac�#|;�����B��,Ȣ�[��r�mV��j�9���N[E}4�n�p�uSs����諻�I�� ����E�Qܦ(^ЙЋ�6�B כ)r�.*�%R
��ċw�\+�o���m)�.�Kr����@[ѐ��<�M�J�,�~�9�|�7Z�DZi-��~��<å"�Y���2��p�ڠ��%�˘�2��7�y�f(Lf����y��dk��t5�r���ʍ��k����g�)kcD\��ה�g�����ܻ���Za0�q�FQ�X�s�"o*��I��q�v���.))ű����F댦
����	YC9g\Ȣo��nǸ��mXQ����j��.|�h�yS����&F�|loyl�0F�=4S��Yu�:�,U�0�<Vt��D'��H����u2;�������=LDgx�_���#e�

�&g�0��Z
�\^R?DpN��� N3�=������-b���p���$&�����ut�����x*�>o�sS�����12�A�:Ѕ�;�V�~{}M!^i4�jM����+��r���[��HH x������LǮx\�<\�rT�&k�lZ���ܸ[��Z��14�>��1&�<B#Ra<�4ˆ�,�P-:}�,i�U�Ek�
�:�<�u"��:9y�彍���n;Z���}~,N�_�q�=f!����?��#-�ƶ}�R�)��s�#厰�Ҹ�X,BJ�]���12D�\����'��O~� v^TG�F�m _3KM�l'&�8p�b���Vj�ƌ���>�2� i�Z��`y�b*��/�x}S��%�o2����Ft�p��Lm�q0�҈9Ɔ�KpɅBN�!��y�xRc���8�c���a�:\|?�#i��A��?��Ew�w��t_Ax_1x�C�z��[߀"�E@��G��[�X�6���7F�`��l��A�O��7!e:l�Z|g��M��3�N�K������g�=������E�#����Q���N#�%>����-rm�XV^�P�+�Vફ�.�j��"%T���vf��_�"�K d��0a84�&�%"��^�Vx����RV�<O�tu��I�DZ���LTv��zz�&K�Z�G����<g��7j,^�\W�4&X�s�55-oS�����P�k����ZuW�����s��Z6�7��D�
���BL��1���� :������P�lޑ�/�KY}L�j:�z (���EѰt	Y}�u,���v�SŁVZ�����Ml�n:_�B����g��as*`3i��D5�d�/���FO��"��x��.;��^��?
..f��"B�̙s�C��U�{�8���нH��>�K��o���>�&"_�����=#���u�B�ڶ]�b1Ox�� �'"qS=3�\]Z��nB��2kbz�`�T��V�GI� �9`���'���������wM���ި+�Q���l�SC|^QP���ٳ&�kwKQ��IOSAi���̂��S?�c%8-�#ЏA��m+Ȼ���h�t1fp���h��C��=������ �x�D�TE��x?a�,�`����嶱�>�����ai��Pf� Z#!��C,e�<ΰ+{���"mu#@��p�:�����%�q_�}�vVJ Z�?�mh���k|������Vq-
�����J���������k��a(�#�����s�����N�<����&�_pQ�"�:���	#����&�[�����?��Z�|�eAji�a�C�;�ja�Ѵnn�Zk��X����Ð�'�>3w$ִ���iK�y�c�m�ط��5Vx���0��4��|`?�Kۯ
�vQ�ɡ_;Z��_�5�r��j}�׬Z�K$CX5ȳ jŝtz��c��Į�Bߣ5V�A{��ȱ�Hi���E0��N���hY&��?h��A��N��@	m����*�����rV�,���б�j�mpi��a�(�&����Ȳ�U�RBvm]��b�@����w&�bړ(OQ#����:hJc�z%�艜|�0ߌ�^���AoF��o����i�w+T��i�Rdō�w����1�Ӿcm�7Z�rII��_��3w�0y�%��Q7�����c{^ҷ������NM��^�����-;�v��=9��7�WD�_j���H�B��`D �WDA�|?�ʗT���:����hD��:��6L祺_lE�G��-�c􋼥�C�H, $��l8ٜ����B�z~��f���q�5��i-
롦����W����g%�?��\�$�slD8���v��3��Wâ"�5S@�}'>�YC�>��hu�U�z�|��<q�6��'���:��/x,{�{oo��^���*g��7��Q�CA܄I� ��E�s�O�fͶ�����M\L�&Q��].w���Pf��3�d�l��yRs(�a�Rj��WE@���j�:YhL���nD7Z���7�M%��C8��T��hkP
5s�`.|�4IM�K����):���" �_}�!,P�Q�Z0DΗT~��Y�,M7���Kz�ޭM�ב��v�ɲ���A?6����6�>@�I>��zKή��_�\��4(.��t�&��	��Kо5��u����71S����<���<�P.c�NK�+�V��}yE(�3�k�7����dH���96��@�'��JҸ�_A_��C���9�b3�Z�P��Q��K�&�(<C/p&��kI����@��8R����Q���^�+ϳ�	V p�to�i����n��tH�������Pz���c�����������H��w"���²��H��$�E��\	|���2>)� �a�:����7�:�bp�T, Ql[�$v���q��5���+��vbw�K�hq�pI?ٙ�BO�
��Y�ֻQ6;����c8�H̆��I��O�S��X/� �l(�Fh`��`	��[�,Y`l�8Vu$� :��l�O_-�D+~��'{�}�a���B�2 ��H=�N����c��[WKH����7 ���l�$���K��6ޭ��.��|̚bXU1�ј�h��j��k�����ٝ�QhF�,�aH��"�q����]�1���sA����+�ĩ�PW]��H��N0_N���	�i��Wj���Zy��x��5@i��?�Aa��Fz�u��t�D��~��?����frE2&������y}�V/��k?	~).VMe��PO(h�$ W�����;3�����<^�w�W��nv0���bLnd �����n�����ɷImρ3���ѓ8���g֜p��4!��2]/���䤫�ִz���\ve8qԮ'��$V^jb��
�=�,!Ur���#4xBʠ�e�:Q�YK��/�#S�iI_�/:��F�klo��L	�R�g"�o�C�&C��a�����g}܃8٪R�"�w��|��ڶF}V���\8�f���fԬ�;#%s>��6�jX��_*�p8űۓ�Ru͜ޔhN�|n���%�/1m�[~��W��[�H�4_C3�b�8���5J� Ro����J��]PSr��z:_�!��Ѿ�W�����6�ãZ�ڌ�{u��BCm�u�x��m'ҥ���qI���b1⫥(uI����恸_����������.���q�> ;|TR�Hi&���U��O,9Ž��9�������x��e=�s��Qᔏ���铠��o�Ow������_���D!-������H�g��������È?^�8���?������x��E���2$G�'j$����w��#��u�	-���@�"?�ތZ����u�E9����t�N�F
vJ����_��	��峢6�����P�xo�)��l���7����vS���!	�m�4I�#��=$(."��"�.
��~j@S���dz���7�\��5�������}'Z�%۵�ʀ�Ү+�G����n&*�bGb��%j��Qw���:%u+j�4-L6}!���u�BA?�P�#)R��4`�N�ߞ�#Ѳ���U0s��&G�̍�D���pV�T��!�Ú���j$�f�������i��Wl�����uwd7���j��^��t���K�n��!;����u3�7��fr��9�.�[��J�R^B�S���`��"\'��'N%=PШ�"5���Y�y���D�[a!+e�n��GNd��dBe���!��ݨ:������#e�-Nُ�y>=�j��.ggL������6?�(�N��Ǔ�J��sh�/CC�-'�c�ꪡpPV����N=�!�BgT�wr5��H'g���U._��ȩ�)�e����t`V��Y�eCA�V������x�]v���uS��6aO��[kvY�
Q�v����m�L��Nl�ރu��ر�1<���c��F�5¥j#�d�B�_S�����7�O��ff|�
��*���L ee��l�vT룺�-���[��s*�+�gX�9�S�FG�5�7'}k�\۵6v��<���7����� ����	h�x�C��sE �UVh��J���v����KLPL~�
NzD�ؠ�t&7�˶P1t�W��m��Q.6Dt�8�������Јt��,�4����6v}��4����J*�Ѽ�"�&�l0�o���Q��(D߶��Z='��]eիxZww���>��W�S�U.Ov�az	����C]�y� �������;h�z讐�bWq��{/L(������Q��Q�y_���ѕg����.S|5ՠj�����Ǜ�5��Z@=O�z�|m"��M�'�g�ڕI�q�25Y�g����.�������ꌂ��`�6�ǂL���Rz��D7��/��U>W��$t��s#��{�¾�wڤ����q
O4�}�<�q �����n`k���j��@�Ȼ�s���6%�t,��@�_Z�������"F���ܭQ�������VW<��}ye���C�.�'�H9łm9�&,��S�b�E�@"��&���L�9D�m��o4��i��f��f2/"F�&�/"U;�uak�l⤴�M1�b���:�"��&�rA-�Í?@ilD���=���@;]��l(��i㎬���9���yA�N!d́�����r_�&�����4�Q�����	{�F��z݌�^�t���������`ԫ�������6����\�F�_^�h�p��&z�����@,/)���M�����e_&��U�P�����hџeRd�# �;��t��>����Y��o���+AD���1���$�"Y=M�͑؏Т���y�!�ñ�3u�)nv%��T#4��W� �@��ٝIr�uJ�Gh��?Iam��@�wH������RI���}_-x%��M�g�[�d�5��R8H�-�ܗ�Ki��>�`��V�-C���J�ڗ�.y�j�]̧�3�������S��YA���yݘ'�F̉1�>��/�u��C���������R����5{�+E��]\��������d}��N#�&���8��b䭤K׌�L�yw6]�� �{o����n��Z5�̃�omҗ�Ϟ��ޘcY����ED=@�@�ȱ�����~�b"-�+@�&�㸢#o�rI�4��א����c��td%ir.PM.���V7�q����� AF�wC|\���^�X����Q�I;fM���_�I������<1B�����	K����H�;d��i|�q�v7@�l�6�Y���h��[ ���NA�H�5�W��\����ܧ�<�w��L��it]���5�8D՝��.\Q������|187����5i"eFpFI�q;�?2.-�]��X<�ȏZD�.�021�( ��u\76L3����:��K��y�׳}e%t��
l�j��R�J5��o���vf�"<S-X�0'ɮ��Do���,��&�.�,����pv��|)�d�Wt��1�o���N�����b�֭��-�����L������}ϩ�ɞ��!��lpfI�N(�J�1�/�?JQ ���ˬ�"Absc"�4j?��6e��!"�k�fy]�
��"�!�Sv":t���K�����ћݙ$#��a�ٟoQ+Z$�w���S=o�#m�^�R�&�sby>�.�&��
��5m�(V��49?�`J�@,�x����,L)*�$e�����4=��6�Kp�@�Rk�.��b�ps�<����<�*1��vW1O�K�:��قe�.��i`�	�^V��I�3F8���>�'*��D���yS�8v��4��k^&:�挕Ŭ�������Q��^A�ƼA2�"e�)3�
	v&\���{d�����q\��f�������Ҿ�l�P9�����!հd#��̿1����XS`2i��Kh����QeA��y<�$ M�7)�x`zz#7Y���)c.�Rc$|�1�>k0S��V�zu��HQpǾ��_|�L����B��K1>�� �����J&З^L��V�OŽ	�VPpȕ�Bc<@?�ռ���eQ,"\�S�6�p�M̆-(S��� ��w5^�C���¯�V�"�[0f���H,�/����\�&	>�b��pn0�� �U��̻�-ES�"�R*5���«+��vS�����u
`��ey��y��f���؍�+���m%�vh����	|�b�"A&�&	�b��?�N�����d���m�R�#YF��e�[���y8���f����D��I�,�H1*i]���1�W

J�nu�)�᭛��Y�3fՖ��,j��;X\6Po-�H���/Y#�bI1�������={M�+���q�����l<�Ʈ��~TD��}'�-�j%"(����V!q��e���b��Xӏw2�� u��c��?y�S[��1�fe�jӐ���|�ӌh�%������8��,���[k��h�:���.�)��9��t��)�_��,Qs���c3�:�����{��DO�����R	J�k]YTFt�|?����[e�䰩bM6�U��}���Dq���L�;!�Z�%��8j,nUb�7E'-�� �,���J��b$�*�[zjɎ�ۣ�i�`���z��#5VҩO��9�~Z��=����9^�Bn.^�>���,���fbVu�۷'^�`%�fU�Wj�����W���i>k�j>��;��aO�������m�͹��,�h9�s�@z��&���x�N�l��7�{��j��1�w��r4���@ڜE�1n�S/I!�fi�x����wO�``i.l��=0IT�4��M�9�)N�L2�m�g,�B�ٺ�_��Ϯ�k�r��$�CV�.io��o͈1��1vn�2B���Ϳ!<�댯�p8�#�~*k��xͣ-��Er���ѳ�z�Y�vF@=w�.��b��lX����y������l�¾qz'��7է�a�؎|��R��ɪ����d����v�C1��s����F�H��#���F%vp@x����RVn���x���J���q��iDU�
�՘�76�ܲ^ԓ�!�>���C�͓�Ӹ�W�	B��(��Q�	!g��c��N~�T��6�7 +�g���"����V�9��VQ�`z.-��PK5֢_�!䗟�t�,�V�-a�<p�F��/S�=�(�v1�P���k4!�p�)	�"s�]rO;�^(q:7�E��N��(�05t��(�i�;��%FF�i�9l6~�������2�eG�&{1�(,�!d��NT�1�ÑF��n�����¼��hۺ8#$��[#��/G��_J��!{J7���d�ۜOTZ���4���L�{��3ȕ����$o���	����c�[}x��-�?3<,��N�k�!�T�u��6�F��A��;��Xfנ_�O��\e��)��܇ZF{57�Y8���΄���Ӑn��n_��#���V���	�gm&���م�:v�snQPU�S0�@�I��	�?S��{�N�4*��i��8W~��� 
V�-�C|�\�U��)��^��|�ni�8""{e�,%R{���w�i�nUZ#��J�n�W�[[�0��W�O���@��������a���Z���4J�L��ۈ��HJ6��8mfoі�g�u�#�5}QT6 }:�?��G!S�4/o��3
�T�lĀzg�|�P�[ �KpK����dR$�'��^�j����G΋�� �t������^��X86mN���l�	b~��+T~{<gB�ؐ��#f�\c�.��3KI 6@�����dW1ʧ}���f��}-$n>�Q�N�K.ت����>WH��� қh"�#�-.��ݼ���p��a�K�Ŧ��}Z�P�wG��Ⴚ��e��#.�ux�fsFw]`x�������D�t�3w8�<�͌�*�o���._����~#�iܻ�dje�,��E�?tar�揠�n��F�����G/ڑ~��C#��Z�L�!�\P)i�d�!N������ �"��ʩ��.�m�H��LB#�җ�H.�l�\�ɖ��K�9��1��hl�=Ɍ�G��Ù��w�U�Q�&�2m	�/���z�m�s��A2
��_�[K
�ԍ��lF������(2�>��%����y���!��ќ:�mP�����w�����'-%/��:^bX�<S0�D'Jr��4���U���′��@~���g�v�������!������Y��	��SBT��~j�tԗ�p;�-#3��]a���j�n��6�>���G��B6�J��Z���ؗN�i��B�"G��XF���F�@`�AХ>���̉��F�������wf�2��7ԃ�u��,k�r����C��y4����=���o��c�ⰹ~�����&�T��Y�.��d�w4�-G�`$R72���S8�(�v��٠�L�Q2<*hXJ�4y�;B;���yi��x������nTݷ�Ŋj�C�x������555Yk3u�g��G3�d6�X����jJ�a�]B�"�+:s�Ga̩Uւ�F��n-;��y�������zp��K|A�6���0�Y���84B惙�\Z���ERt��h�h���o�Ӽ3�V�W1J���X������m!�z�碌>��9d�8B�| �����ͮ	N���m1�P�.�˸P���^�^��}�O������1��|�$�Mn�������O{�|4BbL�$ S�o��Յ�}*���3�$jT���@P6�8�A<�Q	�{l������V�IkзCC��Uw�o�kd��m� �VnZ\�;+� �w���� ��*��$X ^b;ߛ���n� �@U�.�QU��yd����-������,��B��􂆮㗹����%�Q'iB��/��D�=�vr���m�:�|*���!r[�i��9mN�u�δ�6�y(��q~���(٬Z�s%��?/M�npW (kh
үK���=���Rrˆ��/��	xo�u� O�T?%�0����Hg��+2��I��q+)�=������Z����n�4�p��"$䎻�n���Uꨨ��xu��A:b|��:��W�������>���E�p�[O��4'f\��m��:��Cf��ZW��qy*?���h��{��9t�j����}^�PR���
,��H���$w2L0㞲�y�밅����;?��6'�7�ȬZ�ܙ�&�Yp/���Xo23ITƥ��Ӣ}J��W�X��9���N0�J���]P�8�nī���/���կ��Op���'�p�v4nt��-r]�20K�?�?Ycؽ��rd[�g@EB3Y�7oNZĽ�!?i���o������,�$�B��3o�퍃�P��]�zUL��d>&�m��'��h�p8%o,�|c�7/��flnZ{x����O�G��#���!�%Ѽ�4��{ZT-�����4^�pNX��D���-���� z�pÒ�#!�律�3_Xr2����A���;/���3`W�bt�A6D�"�VB���6�`$Ą$�#��9��:�+ �"'El5;Zq�x��Ďa7�<q @<���n�D'feӆ}���ʓd��P��V˖�F�y�l�p����A�����aث�����_<)�d%T���k6�kgZ�?@h]}��T�9[�=B���K'�������P��z��q8�%����ho��k�4��A��gG���\T��_���8}�7R-#��"�p�z!�Qgq9�2<G��U^t��[V��m�3���`�NQs�����W��:�F����P��·��j�ur�\�s�ADzJ�1-������^�P��)�=���7->$9!�1�jd�λ�_+*��o'Ƥ�S>������B�e��d���IGWr��ѝGt�p\qt�������z��f�ˣ�I��� +?|Y@'o��Z���ĵp�?�ۏ�,�Xs�`�=��s��So������P����v�p��n�4�>:����hZ���Q0l�Zci��!��װ�Ṫ��-_w�tߵ@�����f�����5VGD"�Yș/��l�������}���E�ODV#�w$IY,-�׿��2)�=�
�D=(X5��0#�&Y�W'x�=�Z�df'k��m�e���Th�n��f ����������1b�ČJF;�E2�ߖ}�	���n�;#-�q��"J@߄n�}�R��u�吕+0_*�,5T�x2�لo�Aߌ �Ra������h9�v�����u����s�6.8���'��=Ɣp`���5)�ppN������Ip�TN�,�9�a�q���}R�Xn�+�?TP� e?m�]����r}a`�.�&7���ǣ@��:���z �� C�b�	������<�����o��H.�Xvo���.��W�/���R��R�}�sk��'S�ު�� ���"�M���-�`J&�,��!x���Y-�̤�-Ǻ��]P�����&$��FT��&O-�nq�Ο��g��#���ko(N��uh(��Xdw��gh;���5�G�u%���N*�E PL8�h~�8/�w� ��7S�t����6���9�׿��y��Zѫ��3f�#F�`:�h���3ZCW����,� ]�O�$1��eʴ��jmo�9v���ׯ{���ʱJ2�d�����YL�'诚k�@�+��v�=�Ul�ޭ�IӸ�L�"cw	C�PU�K�Uy�a�uH��U��샲Z�V��C�gcq������EXY'���[��A=ܖO]@�8Nߗ1V?ť��`��b!���NF��3��P���D�bn͞���(�J��YY#̉[�h f� ����e</f��K֋��>�5}�>�w��S֝p�
"a��E��G/.��4X�����J�S0��(=�{���4W12�:d8�R(���2������aV�߻�1�}��HC����wv�޾�J��B�h��٦����@X*�H�'6�bH��'`o�T�WB, �b���g%�+@c�9u[�(��YE@u�ܩ�Sx���[@�:g� �?Pfs
t��L��F[~1�Ai;G_9S�p
�r�q�f^NM��ť��v�nc�F��	M�sdz`M�*ֺU�I�[tu���;d%v,Qc�8��!	��K�#zj�Թc[���n����>��<���J�
A/��)J��!�6�X:�ΐ0V4J�eA� ���'  !jR�]�����-�$�s�H>\�7ԕ٨�X�Л�\���V2�У�H%��+,�O��/NC��f(��!@.���ܣgC��m�r�B�L%w:X���0\��F�;�qh?�J�e�O<H���~R��c��$(�D)?H�4������`�k�X���,ֿd�1�,~�~�T�V"�c%M�u�s�y�2p�u��,�ުd ��M'B��tZ]_T�5�R!.�m�Г �D0&Pl*涔�J�c;���1f������Vw�Ą)���^4�15`a��ݘ{H�p~�0��@{���ܟ ����é���~�����?4e]�FwV���%݄w�Eb��� 9l�X%z�G�q�t�_���8H��]���}���6���E0���F����
�ȩw�����g��r�4�~�mh�����B��'0y�i�۝�(6t�B�*d~'�{vЈ�.A�J�0ₗR�R�.�L4�<�$�	���4g�z]��+�ps�ٍ�X2v#_0
O��O�ok�K)��`����xٚQ7��/�_�����ʑ�'�_@*��*q:=ݟ��7yUXe7k�UE�Α��Ly��gkk���%��D��D�-8r*��	���Fͦ~�0'_�<=y�|��)��˱�J���&Z�`����։뒟O�vQ��?Z��P��e�PO�);��&�Y��6�OX�-T�Q���8f���k~r��V��Rh�����	����d3z�A�j2�C~�^y=%�+9����܂��~s�Ձ��z����>�����N1i�H��((h�;��'��ǆP�E#��+�:�b�����T�Ⱥ%e$5���!Z`�9����xr��Z&�Q��h ��� w����p�hFr�{�.�CS�㢪ѓL�`Y�:�����f��ث��ܺ��VoY��^@����H��K�L6��/V����`
��M_��ґ���V���jQv���K}y��4|C�1����a(��QY8���3]�)5��jɻ%|(d%��<*���쀂q�X?ĸ�9H��z��33�:8�:V�`���yЌ�\\H��Ld�b.W����0��;C0M��zȻ~��Mŭ�2T[zb��ޠ.5��O�N����f�����
HB���<[uE͈,�;�$cy�[�׬� [R/��;��C�rk>퉓�pz½>#Pj�* {���1�(*�+��Tmp�V'�#c�@���cz�����(x)����,^g���ζ�4�ih �����ʣ��	�jy�4�g�6�̔|Z����/�pA���= ���&h��F^�24䶶@�ºPi�V����54��L���������[��J�xr��x��oe��4X	B�MC�2��¢Q��2̼��)~6��]�R঻���&�/ٞ�:,L�+v����Pk��K�H˳�ۂ��d��3���?/�#3.I�(����@�h����	(�k�l�����S݂oqJPH���v��ز�lu�#0%�|�[q����M?"Ov����F꠼RT���.�ȄkJ���<ᢧp$5,#���O�P�����ǉ9���������q�z)�����+x5؏�i�H����ɹt3�hJ.�5�ᆓ�3�I�I���LZd���� [������T/ܻ�l�b�
���C-+����'��{W�i�Y�Y5E��M�qI���_z�B��R�!�v���Y,���O�Bd 'A�/�$��4kX"����չO}�BXɳ8c�JRA�k�7�?��6�쑬�5��2o�a�,aY�~8"X?�0X{'���K2A��Фj�\j:rh
�C�ֲ�1�~*t�4��U E<��Σ��;|e�U�o�$��$���/���Ӏ�b���'�냎��7k6��yn/���.(�Jc��q�L64��RspBLڭN��4�54�ʀt������-S����?3�9[
ô�! ��IU�WvE�ۇ�[�hP1ٯ:] Gjt&5�k65W�RK*��W���,q�/"E��T�y\�em��DDX��:�V���xl^�zm��o�{�1�Zϱ�C�@8�( ���I�������_.8�o���JoU��/f�͒ݛ7-jv��r�=ߦ��׭xw=QCL
��2Im�&�S�21���'Ż����-�=(��b7K���RC��/*(�S�V�]EnPQ�dd�]F�4� f���k�ĄA1�Hx����ݖX���DvR�e�FQ��fT�C5����������z��!i��_��=˽�p>�F��x�
�D��vD�<?<v;�UpD�MQf;����7.I[��bM�����e���^L�j�>rU�v�i�Ly�k�������A����߄hdU��l�'hd�+Yus(V�a}o�	��D=o���erIғy���Z��%����c�?iȗO��J�@�ڮ8ف������T#sQ:��2����9���y�6�&�*T�Z�i%��E)����G|W'MR\y���b��x`O���^�yO�k�� ��O�6;1�W���o�;�[�TT>f��NCUTWu�LO2ʁT|೛I6��H~���}CgU���h(v��j5N#�j��O�>���q����Y������@[W<:Ϩ�ك=2۝����P�Ю� }���G�oW�>���\�Ww�խd��A��Kۿ�*=ɒj� �
?X�t-�W� ZZ
0�����pw�hv��Z��Z�y�0���@�6?��:�/e���`ĬJ�mm�=