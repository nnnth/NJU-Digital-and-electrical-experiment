��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��X[&-����v|��y����F���/88=�Ѣ�o�D*f@
kvZ�h>�s��dzUl�������n|�B���s�v�T�%5`��%�o2��*ܸ>%�/����SEk�����B��t
��,��;�) *��g�3)��f��ׅ����^��f�=���+�C��cg����	�~sp��ڵ���\�FX@��T���z� z׆'�mZzc��@͐�1�*Fmw5|��L�ĊU����Gr#������l��?��w�A���!�@鿕���$���Q����_F�s����kW�S�1 ڌu}} ��RN������h�N��b�}��t�Z� v.u���9���nK���͠n �������.!�s�ߔ`�[24p*VS��ڒ�W�k1�zY�g��>��u%�w�]�r�6l�d4R4$6�|.��^��M���`��~p~���at{x�,R�$;�G���8�� ����nf�ǌ
���Bɥ�7X��،w9�ï���<t��m�1`{��+�%��2�>�4�����O��l~	C�b-)�A�^���s�$�M�Ή{�[���O�G�g���r�
�0գk���'rB		8.p��]�ݯ����Vѥ{��f�#�5���v������n�SO�i�4�L���CL��v)���A�W7����fB�킨aM,�E4OU���1�'?���F�#ـ[��g���jJ$%�i���?���p��[����z��&)�?@�Z��ƙ53���\z�a�����R;�Z<F�9V�7���$fz�& �c�^�^䂡��z��K����������8HA�z�
,�����@�kp�����xKB�[F<�E;oI��[1�@tvR7H́�zދ�1�ԉo � �	A���TD�t2$�"Qat�+HO�%B>\\��Bqn@���S��,Z��ޠ%;���$�x޶�WL���J0��!�:�"�����` �}qgg�y�܃��#�;X��/1�������P� ��GD��E����ש�KNN�$�%�"�{%8�� ͠�{Pa�����lneˬ���r2u*��lN��5���T^�N�Y�C�е��g�X�A�RqBb�u��)�g�+�`�t8��F�S��(�Qq���j�E��g!ΰC�;��L~^~�<��4j�ق�]_���|�:,��FB�:RXȅL�<�U��ov�d����v4��ad�n��H��.�TǙ3��ғ��D�a�u;~KDEe?�����ٗ�
sj�����&�i���A��eNh,A9l��N������<O�y�@o(7��x�VIl!w���N�L,�[o�QB0y���q��e'E�╻帩��}`� ���e�Қ���xI��~%�a�d{#�>�/$�g�����奬j���F�M�5�&�k��;_V��z�	�8��4�/�wv��� (e��� %���v44ޯc�K�{}����V~Mh����?ӎ�^�7.73fTī�3~�1t��?u�W�gҩ{��(�&���wQNћ�G[<�<�AN�7Y���u��@�P�6Z��~Lt[��5��Q�Ȇ���#�-�GR���*����A)q�g�¸�F}��Ә{���́�8-5��⌉�Ǡ��y�+ؾ�B_}e�h*�T�ښ=+��ȗ`���	���i��xњ�.%�@�h�݌�F42G���C1VD'�c\~��h�z,�&�*c���oDY>ז�1��f	��߆y&o��b��<��߲ͦi�4(��<E�jb���F�S 9��cή((���)�����B�J��3(��*�L�6c�#M�n[�5������	����������� l{m����OE��vM�2QK�a��dԭ� ��0+��=�iZiU%p����x�-i����DI�Æ���}�dE@X��kS�o�ZO.äj9����]>rH!�@�҂��;]nWs�E/�5��gpg^�?YI!t���4Ӯ-����^S���ץ�����A_It�\�շVm&ܯ&#�qﱾ2�n�;�N]�@���O~�r�Fn����]*}�Rb0��Nq#sI�c �tl ���BS�Hy	H�TXK/ސK��`���;���`Y��b}�lxYV��T�^�X��9cPK�D�B] ���Q���̀g,m�Q����X�3Z�I�����py��b�\��6��f�[��׬琙T��a)/� �aso�>�MC�.K��҅B����"�?_7	����?Ҭ�A�˧�>:y��*���cmJ'� jƎAV�6-/Q��1X R����,& ~1�λ$r���-rg7��`�p+]������]�_4;Wޡ1���1[, 	/�RO��GIJ��5���Z������4�B  �6:��".�{�e�x�U�c�g㣁NMD��;3ڎ�5�k���ax�����Q�/l��dLqc�RV6T�'�)��A����I�?���:�����%i���k+���y��H���qk�o3O{;��M�Щ$H��2>�-���T�;����zK��j�	E��5�����g��a�`�9�ך?� [��*�#�$٥��yũ��f�sj0-���3�KA�|���+X�����兴x7��ZY�WOѻ/�#�L�UCDu`�CLY� oZqÛ���I!�������G�5�s��>��a�9Ў��������&�n	��*1u.V	�B���0�_��!�:��p8ڿ{y���Ѣ���;(�����*���ɯvI/�� �yZ�y���5�t �{K����b�ZF��=i�J>o��$#Z�n�5�}���?3���% 2s����Q �,��~�����l�h(�s���3,Wѐeī�����ꬷ�L ����k�i�7:Qq��㡌+��Gb %����jx>/�i�I0���c�+֟B	��N�`7�M�w夛|��ߔ�o���`��[�؜:���a���`rU��R��Œ���A?�k�C���q�:�d���!UԵR���!M���ŲEj^�W mze:����H�ι�W׮T�UI��yS@Og��S����̑92ZK+JxP��8�k'̃�e�:�i��z��v��$�j14}m��K�V�a�6#_�|�น�]�3z�-DO�ˆ���Dq��� }dd�R���Bϑ`���a�v'�:�YUk�X���g�=f��rM<ݒo%�<������
p��S��F��c�Yh	�DC��~�<�'%\FȮ;eR!�d�L@��s�~?m��#j� 88?����v\u�$ �T:��$m�<u�(�k�6��q;
�S��
kh�aXw�l����8�'�UΙؒ_��x��,��Oa�T�|�Ц������r(c9H�~��"����䪈�p�������� C���2�5:_T�,�)ܠ�S�sz���S�V�H�)xو����2��H�+o��v��Z"Fx�]^=� �`�N�FLe�/ً����R�L[�Ԩ�:�&ā�pj�?j;"�db���� ��Ňx���)C̐��� ��t���V�v��������
{I�4E򤶀����ޚ	�1%���&�@��-�c �d=ac{���K�w7�_}8e5�+�(
�J�w�Q��
����'"J������b�Ve.r�-H��VWҤ&���7T����W��/�
{"���fm�T�g�?�� %�Yϥ���+���tV7��(�E�@8y��~\�O��B���)Z�Rf)41�H�X"�yݷ8p�-�-�t݉S�0��]���(��t�(bn�O߸�W<2��Z��2�P���r����{m��z
aMǸO(��f�4��v!9\k)�q/��%�<$�Z֮�|Q@2O�ϐ_IN�$���{�#�_�[vOJ����~;P��Г����Dx/���q@W!1��9�J0����D���ή�v��M�d��X�����k�qO�O��9��h�K+Q3|�.���J�
��p���h�'�Z@�Ø�j�ة@��)\A�t������ٺ&�͔���"��i+koO啕q��q��>Q�mO�����E�hSц���hw��=v٬�pORA�$�zF�|���ʵS<� 5�i�,��x0����i����-�PoX��M|c���r�>�0��}����C7�n��Yd��(�(�%��
��Ҋ6���w ]�V_��{{d��bNk���!���u��o@'���(��6��5[�T�|�7�I����D�\GMc��Dx��8���R*�o�����s�`F|pEH�d���"�kz��T_���A��r?�E&s����&
�S!裸���ըL�m��#.iX��6�ڃ�����(C�Xjs����Ŵ{��nc$ڕ_�j�w�޶��[�︵Z�M�T��&�%7�_&�{&�G���Yo�/�Y7A�S*�s���9O5�c޾L"�5�T���Q����Yďp|������_�whS?� ʙ{ �O��aQmM^-X�P{��ps?�Q>�;��(��%��4l	�a����>I�e ��u�Ao�9�R�i��Y�9��S�nL��/bx���z���� ��h��tJ�8���n2�@�]u<!uѣ����(,"7��˼����Z��P�\�粠)G�龹]5 �&�J�P���1��!Y�ٌ�w<n��B����pl4�Q��[�&=~s;���;�x�h]�����&�FX�͓���No�t�nc{���G��xI�Kg@+oڿn��������7G�6�|F��9n�[z?ȗ��`�SW2�CO,�T�uUh�E\x��pJ��:�'#[D�(V����*��� �p�Z�|�SX��:�9�4
m�ZrVI�5Q4E�J��r����X��h�>�rf�ʾ��2Pԭ�y����q�o�UJ��>w/�55R nK�44������������E;@G��=�a��V8g��{��j����*�X���8o=]֒��k����g��^_k��S3��#���}zN���sXu��=5�*��Q��]���Ÿ�ԃ���0KG�E�]���گ�x9�L����-mk������6z�D#'&ݱ,�����Θ.�,d�'�v�u���F������EA�=�E�dC�c��F�-��0%��yd|�2����3v��:�=͑�k�V7���)>_p�f ��Y[2���̔f���oٵ~Z��wy����`�Vkq�b��*wg&4x �S�&�~�L�{�ӕ�ُ��*٥��ȿBw�&���.�O1�܍�j �'����D�в�n���]'���Ɨ.:qڞN�C:���̤��1���2Y��ϊ�(M�[e���+��k�H�4��7�º漱#YM풜�~L*	\�%����ph�ݿ��/)��2}�$�7z �*���~�b[=L� dت��^c�-gw�J���Q�q�P)G��`3���e�
r}�\���JK�fAJpF��vY�E ��&Mb淮xЙ��Vm�A��� lv���Qp�dX�MF��%�N'�O��)*=�>&&�U�B��e�s<Y<M$s���%9��L�{�0b,O9Lq�t�B�U����Vcj:�8�B���� ^�ܞ�͚>P�"cv:�D�o�?Fa�����@ʔW(����*�aޯ:�"<�D�����.����Z�yc(���&끎�4�1��_ܵ�!�A�� y����f�L+~�!�o4�d�O��控���f�XPiƽ,�U2n�q(�cD

�Cyw�@uN�*���J�&�vd�H�z����܈!&ˠy Ta�)�E���ȗ��P��&��Œ#a4�Q�:�_RW;�u��W�} l�X ��z�zͺ�W��R�����P�E�b;gA��vܖ]�!Io&-=���Y#���O�?/'�8���wH�R_Е�3x��cŴӇ�z� @OC��A���{�	t�(�����y;N�؝���v!�Xaí�K�,�Y�xI��?� ���Q�h5�mq��:Z�F?�P΂iܬ�ِ�#�$&?����`��nH��Z�?�<i|����_?�~x i��%'��XF�h��D��� ����QC+ҘÊP��]/҅5��0t��1���a����J��*ȓ!M91qd����*���b�<�:�s+�6�z!N� �B9kku�<���~sc?��?ר�t3QJ:�K}��C�"Npk�%T @�}����lu+��*�X����ѧ
�VDQVݳ�^��CR&�?"��Guu4Ar՝��L���o� !F¥%�ы�5�v���3��n��)�h����@���h����dXD�+Q#;v�Al��������<��:��U�9�:��4elstWLe���g�ڬ�����!� ���fG��5@�V��~|1*=3%��̀��_{�\��==�.���#�]�xP �ՏQ�t��1(�w� �Y�v���Í�-�3�#����"?���a�������6����cLz�iM5-AE����}j/1��)�دl[R%�`��:�d����qPG��ϟ��a�?��.m�ư*._23�^���B�L&Qy����|���O�&�;}*��Åk[B������������J���T�!���Ĩw.�.�{H�����,Qhv�3^��/�Cy�1�N�ں�����^ة*���x��K�9�u�������U_�c,�c�&�rm�*a�wo�_T1�O_���@�hɐP0U��̪�M��./엋K���~��۞���f���է�I������Je8)dx��_����=�ZI`��Ѕ�o���]��;>:� ��9,
��2���A��ZJ���5\rY%[�����.�D���jV_k�}w���16�BX8�Jo���
\z��p����ޚ�o���V5���S�󞯔H����p�"�U�ƕֈR���Jb���)?\�D�^,k�,�6�H|�b���Y���.S��K�^�:��}����@��-��[�^�S�p������%R�R#�^7dGN�a�s���Gb��{jѪC6�lO���%z�Od��KX���@0<�\O��߆x�Ԡ��B��5���$9Ǚ3���6�ڎ�?��JX��Ձ(/��n����"�����HG ���O9���
:sz�{�v�0�0�Xvi ��/���E	��Z$Ѽ�'`���^�T�׀4��IF,o��=D�����
�L�ф�5=g��禁�ê���V�0Q#Ͽ�gU;�
�碼����.�y�����P�Q:0|��*���:b?��9d�1�Z5h����@P�xP���=�7���1`�aw P���V���q�"V�>M�O�y�<h7&����P�B����P�ʰBɔo��(f,�{�`Yƭ��d�}60Ċ6��I4��y�ܘ2F8I�4Q�� �<�r���9W<hJdL�=S�a2%�7�MYׂ1�c�-%4� ��V�ؒ)����b���턢�zGvn�M�yn!�� ���##V�����Et׋�EW�{�U�&tk��	9�N��*���(�)�ǈ��B��5C�O��)�h�����oEZ�p�tWb��4�ʀTx��1�4�Ut�C��f������?,��}���u�%y�C��^>��T5thc/�Y�I�F�3UmG84��,�;Z�ZҶ�|�׹��yP?�G��I�m��2"n]�4�<o4a<�O��߃Q ���f�H�r:p�U���R����r\D�e�]�&�i�;\v�l��&O��g�N����e�՛��:����뼜o�g5�(��c��>�B*���o�9^iRQ��m����X�		�bsˊP�ª�dU
�3PRm��uh*�<�0Z�ֺY+���;���S�]p�N�JR6���Q^�yq�a=�g���߄`yj�~,,����=�����w?~{sj�	�9
=���f�4� /�7�J�ھ ���- ��ي�V��x���<�
�����2S� �5��y�a�3Ba�^4��VvH�U��?oY!v����q,u�ڹ�nJ?j#����y�o��M��H'�Kv`LF=�԰p�p5�]tUJ���o\U	O��gj�S�(�*�/��l}�h/P:�dP�5H!r�V��p-Ԑ7۱�<��N�}����&{���U����Z��N%0��n`իS���+��4Xd�$C��k� <gmWy<�ek>�z�t�G?&'~��p@ugS���v���=�9�^�;.l��VO���1$�[�&��W�[	'[�ؿ�*�КBE��N��!*��1$��`ƚ�1��GT�.��I�gD���q�k� ������CAG�G�Ѭbo�QAў���Σ$��0)�L��ɛ��{�$�١O9�E &3\&O��V#����l�U���%\sq�kT���S����햀rH�x�P���$lbK�2���Z��/M��D��~;F�A�/��w��=���r�ZK�S��g�-��j Re�Хa�!�e�b��\�8$�S�?�,a.������F: ��騩�2i������݆\|z��1�ჯgE���vK�8�Hy�1A[S_*��#�*���n9���}���ğ�ո�����2Ip0�e�M{ae����o��I��a�< Ą��/m�>�&V7�峍�U�e �=�ƴ��@C�#?y\)X�0�F54N�L�2�+ĥd�·��u�g��TyP��B%��]x�cI���?�d���<���}���"XD�y|kԦ@ی�NP��wM͛�m޹7��P
 �k�g���fX��3p ��+\S1)�!��P�1����<�جƶ��,��c��)��͆vE m�1&2�(�M so�u�Qf�]�S@O��VC�c�2��?�=��C��֦3�Ԕ�P=��w#��>�F�D�2d�[�ŷ4ƪ��Vې%�uy��i�����VB�ʞ�
�t&<9|���KAgX���8úMlj\�y�����.;t�u�^3�x�#���<����ᕹ��`�-Hp��JH���n�)
pE׎���"|}��Ᏽ̜*���A��h���=��s��G�~���⫷ac��J6x�HaL;mƼ�G0�֘
@��$0+d�x:�S���!2۾�1>�>=5h�n��Y8mc����/R�9�q��4"��(,,���R/�t(=�Z�F?}n8[�t��7A��IiR��~�{��+�&��p��od6��k�]�������&H��?&�T�mt��p�m�2�cl�l7E_u>��Ct.��Xb���a�	��"y��4��i�x1B��D�xb�m�r���o�ǒG5����K�6s���@���cӏhEڥ5w)~�%��_pX��-���`C�T-!�|V�a�P��H$�o���5_+�ْf�	��pv�4y�� h�����w�)�|)B�y�!P���](�9��>�W�Ĵ��2F;[��-j��$�����(�=��h��
�s9�Y�7��	��(*5w'�;^�w����D)�_��>ݼ�Up0�K��%{��H��Sz��Os�C˩�<��%�S�r���we�����-��}ݕ]8\J�U�t,�����b�#�u�g�<�9>^�q���_�|�����x~2 ��A���Ҁ�k�*�ri,ah����'�?శtš?�] ��^)�O�86��8�{=W��w��P2�A����uw����R�	�)���)��}ѵ�s�V7N^�|�5L���h
R�ȸ��댿��4�?LӁ�r-[����N_?#7Z�<	T�ti���ƕeKTE�!�fh�<i���S��6�Tj7�{N.	n2�q��p�{Ow���?*��!��6?�sW��HLr��7!�5[�G���zi/��t#x`U&�r��j�4�u��>R���+�`P�xpa2h�'���-��Z��|� h�I"�?N<��a��{.e�:���ce�4��֤o�
�;о��r���潑	f]�0�o
�9Z)����q�w��f�w���36��-���r�����I���7�{�>�@'��2��+�^�� *f\�rG2�#�L�B2.��6��7:B��D��3B�L㸎y��A�n��\ձ+����*���}��ܖ�5Mj��58T��\�+uS7U����Ľ�+N���K�c�VHeq2k�����.M����Z�a<)o��-�A��&Gy�C����Qk���W� '�K�<�EwT�^���y�Q�-�(�e��V�oIlS���O2���Q-:Qȓ1U*ˑ�հ�.��e�q[x{(��1r2��d�ޭ��L8�3�sYs��GĖ^򾃊�f���o���K����5]3\����=�6>��O>䮽�Ia�3`ȭ��!z�b/� �d6]��٦�`C{:[�=8�`h����"�t� �t:l�>� x����x8�7���[�����-/�@��m�&v�<��n�M�jjAH���*/%;U1f���}NK�s��sJ���>�R;�c{�p�������S�}��ߵ�-�f?�p����,p���H\j�.$��8f�L����,���é~�k�*w�1�F{�c��ydgPV?uNn~s��&j������,x���ܗ�Ya��Z�|4Z��ft����$�tX2�{N�Uy?@�T��mTM,����{���m���
��� �gQ�����]�no��Cfolt�V�X_#��\�Ȉ(}�bO[�e��Jދ� ���5��2��:=�nR��q7�HY]_i5af�Ҝ��yg��1]�C&���������N�8��$��A���"T��7S�{�##����Qm�FV�0�inU[��S��_*�i�)l�`��G��Ph^��2p�tz�g-s��G��x�f|l�o��a������n�W=��~>���0�䑿�J�:W��v�0��p�� ��x���L��Q�������K{���&X� g��m�=,zԚ�jn<Ā�Zb�_��v��Aen�[.��u��{���u�3�㌖�yՒo�Bn�O��p9r�ʼ���he�ʹ��~�"l��S�c'��. ��wUX���4#]�
�v)K�9p��*E����l�D�'���p�#u�N14�ce:7)�ص��q����3@��Ƚ�,�z��(Y����RZ�����6հ��}�"+jI8�4Q������>(V��>�;uY�.R�_S���BՕ�3���|ϙ�Jژa���&��S�m31�Hd�"��͵N��;ʕ�1?�<q>wW����2cc�iZWb�а��^�I@YF��n�'��w�ئKR�;#�vW� ,97x���LFyI��j'1�w��Vp�K�(��B�l���+m�I{�.��S���u�y��7X"ɂ‼��U����^��ͤ�՚;ҿ=���`��OZn��9ˈO��c��/��Γē�_�F����Q���(�J��q�z����P�b���z�n(�:[e�
�����Xz���:��-� C��a�����H5KCe2ƴ0�̃�9�i隽�q�����G��5���-�����>�,��Z��ZЏd�<h]���"�Si�n����[0�.�{�1�3S��Vq$j��³Ԋ�t�F��d[`~�hS�N�����_��;ԇ�^��W��I�}`�b���)�a}_��Щ��N�\�i���f8�������y��m�*�7�/����s\���	5�w2ߠ�4p�{Ʋ�ePt�����-��
�ЌRl�Dڱ�tʜ.�?O��`ٌ�~pt�7W�p#�K�� 9�[��E1|_��@c0 K�k���<!�{t�v��"Hf�5���U���~�D!B�@�  ����wJ��ʖ�H�?���o\N�4ٶ=�e3���İ�9!9b���KL�H^(/@�:21�yrj�U�j�c���2p���%R
z=N�i�|��ؓqҰ��]}���6�����˘�N�,0)�id�� v��Ҿq;��+tmti�;Y�!F�uv�l֬u�4Ÿ��WM�	��֌č�l��NkteN�}uf���a�~TH���56j[�@��Z�4�IUE�Ձ��W�	Sh���d��deC��p��f���o����-�t>�t@���\u�P:\�m�ES�ɈC�r੝X��|��6)�b������y�0<����T/� ����(4;�d���)Q�0��L���o"==%jѐK{-�i��x9B[�E�@�}7=��8�|f��+�Æ#/S���di��ŭ#oC4�\.�RWE�l�m=��[�_������[$�h������7o�i���5�	��E�I
�����[2�\�zmƁVnOhb
�m8�^;�g�N�k���k= ���� qݶ!�`Z��P}���a�:>ۋ�b/ag��Tݕ��\��(���Wߗy�;Rn�(_mHBr�dn$@�h}rnMg��.��"���0��F��TH��=������`@z��I�^Լ)�$��tn#����*$�;�7��/����_,�"�o
4K�|6uB���rO|��Y��>�M-�\�z�S��c�5�-��Z�_�k�I��� m藉�r�0u��*6Jn���k,f�����z*�$qcb":���������}�*ðfA:��p�_Һ��e�^ν"�����,-k����x�������Q!�~K­Sp�5^`�ݿ��a��U?�I��Á�v`���P9����'D� �[���ʷ�G#ۖ�H���h4��z�7R����nxC�G��=[�]��r�e�$���?��2+M&�r):���߫�c�����
����#��pP�$�`V&���o`.]�b�ZAk^U�<4�x�,lj��J��)���ܷ�pZv�^6��\���RP8Re t
,��_�l=0
f\��Sҝ��|�T�G�ʰ�x7�xYb�X�!����,d�e˞k�OK[��2�v���q��K,0mOHe������ڞ&AE����,��ψ���*��*]��d�l�1����9����$�8nV��W���(�JKk�����3��	&��(/��Ac�H�HiO�uS���}�$�E.�fS$3�>X~C���+�8 ]�I�D���'�~��K��i��x�
e�2���-��a~{Y�Ȓk�:jŴ�ɔ�=�t5�d��1
nd��]8��l
�1�_�y@�Y%k.3T��]�oQ�����M"����b�EX��@a6>��z����?Ø�G���G�����#�K�F;3�֕\1lA���?��`{���B+�H��Jm��+?{��
��4�!���F�[�f�\�Q*��۹hմ��=T�?Š���mw�58�K�.rW�?�G�8A���&:�.U���I�� ���3j�bM�J,��W��j����(�.`�4�+O%�t��C��4���V��3�Mz�Y!*�/R�������o�[z��{v���rTl,%��\�a]�~b#���h����ʪN�j;
�G��LnwJIՠs]{��s��� ��b�˿�x��Q��XM���rv�f��=��(�G\�3�a_]�@ M��IoU�>!�ꗢ�^�^�o�-����w�B\w��m1D�|P9��0eb���H�J�7���røm4�O�.�@ܲUp�`�6�)����y�@)�t�x���2�ZǮO�f���\����y��M�ŗ�	��U��D;҅�'�" dT*v�J��b��r���+C�+_�C���)�5Ի]���������+�o�߀p�Sk���.��b%�W�|����!�o�Ӹֲ���m���4� <=P	��M��qE��.!�.f�c�DpȲ����N��
I�<,���UOi��Ε3����f��w����l�E_��P�Q�ޚ7/e�%�[���V!�a~&c�������E�x�>iz#x���a)׷�`�
�	]�Ѳb ��F�B�-�'�t74�"�ÜfR	s�s�e��;u�`��{֓tX�b-������� H��X�8d@�2&SU��ޓ���?{3���]��4*������r� �
L��|�I.�3Wؙq5R"cp�B�Y�`*M��
�ǹ���,�2@,fٓy��lZ�lb�k�����J��d�Q8���H��ԛ[�SJ\~�9�H�ks5ը�u��6��wL1(o-��vw�2��.�R��i\vDҺ�,_�@�L|7�2��64t�.��A9��*���Hv�l�3�F_�a�a�6�/3'A�!�\0�*f��<���j�� o�9�5#�q�`2v��F@2����qO��U�������s*������k�y.�v�8���;$�����ƞT�3�,e�:B���U��Ъ����8�7�|�y�(\�^��e�lZ\�ٲ:xq�p�����	©��_����K�'0>��̢�c����Eжl��f���#3r8�c�6����� ���,�J�[ݐ�<]���5��	�o%۰<Z�B��#7.o��p<��tH�-GR�+1!9����Ahq�ju��"at%�<0��\�5�`��)�3�<f���b�gX�9�on�Zhє)�Bg���h����_v&HU���S�)Dl���"*�o���tx���C��Wy�K-���X�s~MX;��E@��E�t���MVa8�M���@p����wQ��Ha���K�T.��I������V���=�1���Y͛
$��}dL��(����e�T�F�x���+��Xʲ�h/4�|t̬9�r�s|�{����n Og���8�Q@���!S]�á;���#g-۔b�]�eiĩ6�M�M��m}N�Yu�� ��֢ ���[������2����I`����a����t���(&rY(�:6Vx�['3B�A}+[Z���w�K>���&�2���aw�ݫ�$�'����T�V������S_�n3�z�hL�vr�zI4J����6U���X*s;CP��6�m��,i�K����q����`�l���\UT8�O� 1�R��*uG�*ƙog��$�}��(��
���#�"
@ل��c�Ћjpc$ɥ�o���)��Z�N�A�6r	��YRM0�òE��u`�s��Ԍ�^Q��9\mxh9�A��6.��� W�@8��+u��A���vƛ��2e�+s��8u�g�.L�]n4��ޛB 41�_-G���("�$�^����;��C�����f�mǸ���5��8��,�ml�~̟`�����b��;��c4x��w�Y��������)ّ~0�x9L�mv�(�LF��2�cw`�߄����)~�V4�����Ս��B�$k	 ��4[�5G���RI��,�y�L�	�\fIΧ4����V�\J�;���Uжq���֥����Wv��D�L������X��;�h�,�:7ݹ'�^��YKwBm���gJ��E��eA� �ElG���@������QϜ��-S���XB�@3cK�]�"'~g����G��F�`���ק�3��E������-w�щ �[�����֗W�h���1/�փ����9br����P��k��[�q��E��M�Y~�����c�gH�����Ũ��偵��h���ޒ�೮��Sjs��q��l��	�2#�]O�R<z%")\���)�'�"6���+���������4�ӶKK�#��'��W�5v�+�����8�~{�2��涖}�m�)L� BFJ��ꋕf���`W�
ߋ���(dͻ��33t�s�v=BA(	)Xz�%
ْ�j��N�������t�m	�ѐ'�[v�!b�����tn#_:a�N�c]��[M����F���y~�F��)���k��~G�_IM�*[�a���l�PZ��ZߒS�|��!�")m���V]�`��gQW�V�Iü=��h��gao�&泿�߿��'��'(��^.B܉o<9��&�+��H�n��s���S7���Mc�J���@�|L����&�q�`D���()�r�����5LqqHLlȰ<�0wdk����s��qO��\@��FrM�wh?PVRlƋ�@��a��\AZY��{'%߼���^�e㪵C�L�c��s+Je�R9S���z������۴����z �n�A&﹚0�FX���l��o��z�9v�
�_4�L�Ӏ�7l�f����g�D�;%*�]̤	���g���A��n�Dv���"%���˲5�k�dTkg7I�VSY?`׊���R�����i��L�]���MO�~PچH��3-\v��Ut�� �(�p�k����kb� 8�XzO�5�m6#�S�3V
eu2�n���e���+���ܝ�`U����|�A�h�3�zx�D_�֨j �M�W T)=>���U��׭c^ؕm.`Q�:Y�B�fY����ۊ���3��*�N��)=�F�F��ا�_����*3�$� *�7��2�K�0�v����x2~��I�X݌���`QBh�=�U��W��TVbCy_�O��ES��!���sp0*S2?�x��:}@�!!T�J���bjDxx[����?!�	�:�ǟ:a�''1L�F�׹�V�Y��ْD�fT#��`>����3K��,>���$;8��H���kTl+w��4��	ö*{W�!ڗ�U^P\��yNh�h�rj�W3�`t��3���!�o'���.�{	-l�e��$l`�hL?<�(T���@�i_r�P���:Ó�b�ko���M�f]ܧ�J_����H�5/�D�s ������ty�6t�&�"SHI�	+"h1�WJ�P�ŪE[�.0a�3�)2�}L
V[�G���f"��e��"aGY����&Zg7Y��d�`f�8_Sa���+�Rg�*���d�;�$�xTn��U^)�C� !�-�i�r$<�r�p"�x�u��)�UT�'e:>�?�%�Y#��L�T�c��0l��p��9w�����Q�?����t,�a���G>[	�q��$�^�����d~�uȮT'��G�<H��D�� �ڐ��`5~���=��xg	�ͨ;�>#��F���M����4�]���2�n�<�o�������VC�Oc���AC��p��{8�#��U&_'��e���R��N�;�6�,-������E���h�PVi�!/C_h����/`o�}��P�:�)(o�������v���%�^ގ����ߏ�''�z=��8I��a���Q��1R�)?�&�e8��mN4���sPhEhM�2SOe��>�����;��i�<L�Ku�G�O&П�UuvEi_�a�P\��t)b�^�>[d��"lG�2�vF
��Y�
�MJ�0#g]��-S�	�~&���v������Z��~����O�i��@��U�z�kQ��Ď��@�ߑ�<���W��t����4FuX�[�b���Qu"hq��!V�q����W�OH`�ߎ���E�}��F|Q�|���y��*�MLK�;OrG7�N�S'��`G�UBG'=�����jS1��D'�s0�<�al�d@� �v�jA}m�n ˉß��S�`U���d�(7��ʧ�
;>t*��<AV�8��m9JH亣e.��F:�,��U�;�1a3j'7��m�w��S��s��:
u�H�D\?���:�a�TM�KĆ�d
(@㊯�>ô���X?�/ T�:��W[����ش��}�)��b�qKV�W�[@_��eهk@Q� �2����x��
�'�w�yt�}�^~xbJ��^��d��^��%q���2p�MޓўQ���| ��y��1�B
$�-��������������q�z9țK�1uS���������K��_�cN�~�א���7-e�F�2F\�$և��u�0�ic�΍�2�>w�x�ns(������-y�dؖ���b�����I�52W�]�/m:����T�%s��F#���9xy<؎S\<�@y7B`n1��uEj�A~T�4k��j&�d��=[+⽽D�g9�����!��o�j��]Ô��b ����_)���3촊�U�����g�I �_ەws/ܥ ٵ7�"w����62X��q�x�/��"�a�N��d4]���N�9�+Ǭ�|��)t��p���3��x-"y-C���ɁFͼ�V�*rB��Z/���;@�������G��x�<3ǫ�� �hiI�0�mb�L�x�A�;��ge��5@O!V����\:-&Jq�6��$�R_ҕ�^ƫ���H�"6Q�iB+������nQЌL��~l�v5Jb�b]c���#V�_�-$�O���%��� :�v0@yQ�^6E߈�D7�s]�%'aH&d~�E6�RO�m��7M|���hI̵%0U��̓��2V�d\�h�F�!����;V��b�4m�YX<}|X��� Gqz�	��0j�,�RM�@+�6E�[�P�T6�L���yż3�	8��JN�}i}���)~`��g�BR�|�J�i�x��T�W���o�\d�\�;�wL�&8:*�C0���#7��'�c���'n�x^jg�P>:R�q�l��Hד�^>���2�ƘY���
������ 1H�� �_��q&&qT��䘼�W#�����%R��
~/��"�y��ō��/��@� {��X��oJ�w)��y�E%�Y���/�Ps��&o�F�Ȏ��ڷ�(]��y�{����txxp���࠹��Ԯ@${!F��YP�̡`�-��2�-aaP��\���N�luzZZ�p5�
"�_�5��2�75��r���biT�F��8pr�9��FcB�Z苋��;�W^:�	0$�FC*<q��N���J��Ԙ�怜��]٘����@�8{)�I����wP2+݀�	Ѩg�1����R��eb8����n��ĉo�{�
m�I�'�)W�j�B�$c{����m���%��3P����H�P��V� I�.0�Qo�Y�.��9L6�J!_�D/<��Tl8qL�P��.)[V5!��j+@�\6p��P�-F����d�A�掳�z+i�|3N���˳��u�8��惁�O�Ȩ\T�!t�T���r��������F{Ak�%Lz.u���qR�1�����{@�q��Jz�eLJ��@�lz��@��!cE y
T}C#h�׮�o���bc���zE[�od�_A��ck����ǵ�@��Ƹ�ae��컛�%��!�ZI���׈�M��}�m�3$7�U��µ\a�h��ѥ����uy�t�����T$�b�p�a���]� ��[%��ѰA$�ѷ���x	jF�. .oD]�́mI4d�Ƶ��D��=��<Na�-C2�u"�,f�*˘6O)X`��hY"�Q0=Յ�������$2i��mkAq2E�U^������v���P�<3��t����n�8Fnf�̏���D-A*�0�"-�u����A��V�w�hpoz8�GZ�� ]$��,ܩ����q��@��\`AϟPa
Б!������A�"�[{%��
u�v�0��!��� ��7��0kHKqT�E�f����i59������2�rݮr�;E�^��:�D���X�N$���T�P7�w�ל���<��`��l瘐�����ƫ�G���?�X���R(�u��*"������n3�$�[�T4���r⫻�����O�{I`%n"%�/ڪ}�^$юW�^��[��=Ɖ�����$�����4��趔':������Y�f�$Ƒ��F�-xl@?����h�����8niЏ�2��\�=2J�2ȕ:*�(1N�`�E�Z,�9��E�L�p+�FE��et�t��^Of�c�E�ZD��_L���
d�3i��`M���G��k��#��-��xN�W�Mj��g��]o��؃��װ�u@\���IN.���dt`��:/���S+�����X�-D��Qp�.[{���,*'Z9*?6R0�*�~�_T)��w��zJK�[��(�z>��������� �[���lB)��
��QR·ŭ5-k��:2O��F���(�9;a�x���t�h��jY���B;`ګq�I,�$%_��i�$��;Ki�,h�a�>5�U���9tl�\ɇ��N��ٷ�A�v�����$�볢���D��	��k�V3P��㋎��^k��D.Z�[�T="� �%���8V��ȕ�e����3-�9V*��4zW^�؂|@#�tS�3����o�XW�yq?.�������h���f��I�wИ���[i�O�g�R��>�������s�Y\�����a���m�-�1��f)�h�b����`�p�2�v�zM��l�e����݅c$�������Ի����J�����\`n]k����؀m�O�vY*p���qX���$�>�yK��Hp��[	Lj?��X)gO�0��KC��R�oڦ<i���@ �E?�h��{S�'���v+y�D
���KR���M1f��s�Bbht�,�nC�8�����P�\�S�5��s_�*�.*���Mh�/�@��8�6`!�Wp`����W�E�}�3��.���DL�W����T;o�=�	�M0o�@�Ӭ7�_˪H�F����e���k�����'���h0��7Ch���-ݣֳ�o�\�}�J��{�������~-X�'k�"��ԩrn�m$:�d��"�[M�rH��[L[�4ǉ��"{L��-4R�ȍū �dk���$<oT#7� �.zYj얿ɓk��3hު���Z���=%����ⰷ
�Hi>J���0�36�<��mZ�ٌ˼�I/l��Bl?;>��zM�O 'D�&@b�v`�©1ڇ#}��̠�!e�lg�4��y���=���S��`{!Am�Gu�)L�9ޭ�/����%}qh�E������ǚ�6���X��7�q��>O�̕��!_Z-��?�"��ԮG/����(�/M#U�
K��p�:O�&o�l�[|tFI�ɡD�@N��2.$Ҋ7�V#Z����bz����E�U��aG�M`�%�|�{er��)�
ʬ|r
\>H�eC����
U���b������ ��l�g�|G���+����ܪ�������uo���sl#"��=آ�8�Ǟk���}�VSȔ
ƕ|����Ӊ��h�[*�eL��bL���0&�0r�,��32^�'܆v�C9�E�D�ʉ� uCCe�o)���Q����%^�|:#��6&~���u楲�zka���#;6�o�1i�i�S,1ߵ�ϵ�u^n�C���L��L|3ɭI��:����>F��)�af��]*���u���Ѵ�1��^C�{��K��@���X�*Ez|h�%�!����#��78(1F���5W���JJj|*�F�ɚE{�
}�|�����u���K��H-�}��v&6�q���|=�uzP���r߫7m1k5�x ؁��̓��	�t�c}�y�����7�g���m./�a�o�Ra#;�@&���~C�j��yt� ���@��n08�>����L�Q���>g�4��;Sǵ�q�B�	����Zq>����)D{L�R��P�;0�^����H�#���闀�םz&�<V�$�Ϛr%�������O:�\��+֑�Z�S��r��^�pb/������a�[Z��Gܵ�-:�
r����V
�Ȫs�IN�nzvAe�s�`��J��R��$���N�?�3����=�ǿ�t�N,�8���b�{�"��[Roz�	��u�V�ׄj��s:F�q>��s}�6eܜj$�uP��j��k�8=0���q�E<\d�s&�)����Ѳ���&g���'a���xIֆ�N�0gy'��D5p���|��(AYA�����U�+�jy
�	��.��u5m,ˎ��e��o��3��לx�Ӿ����������^M$���	n^ �����;�M1	�q�n\�VC���>?���m���N�eî"F���5*6-eD�s�H���ɒ�SV����5a��Z�m�j�oQ��b�����ڪ�>�,HL��M�H�$�X�D���tB��w�Ջ>^�l�4Ř;=�{��p�;���V��D���#?)5�O��	,��hn>K����2��TzƋs:��eJ�C�wl�gh�l"����S�(��"X�o;ͮ��[��^cnG��\N�B���W.c��=�n����i��.fzkA�,�Փ����W�/.�-a�)ҕ:������w�N��1��r��4c x�"y֓�E)[���,ͻ�6ۓȴ#�G�*/g��+��D	4@M��γ�*�lw���^�wϔ|u�O��Ϣ�c�w�UB8�$-qW<������t�B%bS�P�AA_�4~�,��"!-ϏpPi�W��N�_'�r(ێ3�E^��
����-i5�y4&�N6��<�U�=��'X��B�@��1u�g��ڿH��l��$ن�a�N�� 6�^|�YD.ʙݎ.k��t�R�]{���O ?�,o���l�a/��<�o��p�Pr|A���W���iJO2�^��n}2�P� /�82��[�d:�.�[�<㛭.|f�@kذ&�`:��>�/*����(r��Xf�Z!\r�h�P�8LN>����g��v���-H�Yq��k��������pQ��0�gM�4��B[�X��V�;u�������!lB�b�����g �'�:�:�OA\ʗNW��4�p̅<��kgS�5J�;�)�'�#(о�<����n�2Z�XM�^%w�L_a�yiaz[t5��)SM��Zfo'���!�Ik�~<��1Ā�ڈ�
�>i��a���`�܁�|�-�m�O*L',8�)��z�h����CL(���ȍ�^�x����p�r�������]��t����5�{_��%i��loP���X�J�a�(��T�&jg<�uZ
yL |x��sJ+����W^)u�v���-�"��ڲK�sX�H6��U��|q�:��F?�fy��V�!��%W=�5�HtU�[V`xCF��^Y��&6���6��P�zGꆞ��5��N\}�ኵ�]:��>R�i�L�ӂqﮯ�l���-
�D��a��|X*� ���"L��	�2��ٍ��	���w�W�ҎOde�pe[b��K�v�0�rO���b�*y����.�|M�@�!C{N�7փ�c&��t.����I.�z�%g�B+���'Z\�$+�K�/L���ͼ�+B�O�`bRj��/�Xh�U[�\�����U�\��b��e8��Q!g(�2�P}�6� ~��0 �?�rp2�`6���EI?IAnʙ���	�����t��	b.-��B���cV逺�1�ly<��������wՙ���q������]i!-��:��Su*|�>3e����)�'�s����[�+�7���`?�0��"R��G�0=��2�t��R��<o%��>�<�+t�`X�i��F��z;��l`�JAg)nO[�2��R��>[�X��j��lh���7�>�L���f��g��2*0��Gn`��Q�����9'F��y���� ��RSO;˶��� $�:a�/k<�����e%z���=[+pv�Ӈ�#�*_� ��4IW��m���Ls�ޞn�vq��Ѿ�y4���@��8���Բ��ʲM�U�C6=&��5�g����C)�ߦ�_G;-�Ld�<�O�z�M?	~[������Y{og�h2�����mZR���c"����¤k��#��.���=g�	�.n�܁߶j��M���c�@3�I�.��M�^�s7tj|R�m��E���Y|�A���F�H�(��<�$q�4�Uo�󩈀R0L[x��F� �+���
��!�%=#n'-�2��?п�?�_���(�o[勶����M�� �@���l �8�����&*��|��B5�,L�Y���BZ��|kB=�r�=��y�jХ�i��(cK���%��U��������>)��ǂG=��� �R��
?�7:7|<�bxm&|�0jj�UXXq�d�7���KU���߷V��
�P�"�6�p�h!��H��tg�+�N��[�6�k��<�	T���A3��*���(���R�V�e�&(%Y���S�Iҥ�k�&9eT��t6�t�D6ѣ�K��Ɍ&���N Q�$�(�`��m��f�k�mg��,#��]Snۙ����?����~W���Ǆ��w�>衫�$97�Z����6s��I�˯�,�H>}ś"m>���E����Ls����đ��ֿ�U�8�d���d`}�H�#+3K�G�y�M�Z !����I<�F7}dd6��������(�{�7]>�$����D#hcN�!�gH�e���׾�`d�x����n ��$JȮmt>S'��+����6��V]GۦK/	f�e�c� ����M�?��z ��o+�x�v�X�,<Y��U�1���Q�TF��I�L>�j�l���N�$�٬��mJ���Pm�11(�b�M��	ņ�=�O( �/����d�J/CYz>z0.U�@ Uc���*�;%KFM�+�` a����@�����,z�4k��N���HH	gO,4�Qі3_�@�c?ဲ3݉��P���
��Mۓ z�|}���@v�_�=�V�������k�X�@�Q4Lq?�!�*Ř���;��2�f�O;���ZO��7ld�C����sSL���L�!ݹ�Z�m.��7?�S��*�0�����o`pa�W�=��&��XIG�U�&�gfS�W
�R��7$����ݙ�l0ل�jɆז��$c�F�����CwJ�����p���(�K@D�f!$�m�p���+��X�Wq���z�6rܲ�&r�g,�^��Z=R�7p��cg��G~����{��
H�
� O��E�y�����{2X3�
�+�5�t*ϲ1�z�Dx�ԡ4��W�k?a���:,��r��;'�F��7�I�����7 �*��b �v���6c�p�4�{�ϝA��G`������1������v��������=�{;b����1��?W:e/���%ߓ[_6د-��`mr�P2�@���{;�E����_Ec�Y�l��l0#��z�A ��,��p�I`�QYQ-J�!�"�V�Pꪧ�-a[&�|�<_�3�E%qs���m\9(�/�I�a�5��N�o�F�4��Å#��#am3A��ed �7!�!��b�a$D��G'�0�lY3&�#��D������[jN$���	U�>mȦ<*�ps��v����aN_ �hi��	(���v�(��V���pUOc�_��	Ag?�|(禭�@��s��<��VPW�s�7B�*6 ����}�/?��,ڋ���tE�A1�s������	v����l�}�?�u�c�4cW�2�0�:-��z��6�e[sR��C27*��\ ����aY��i�5�7t�G���m��ձ�rl������*r趸V��/za�����F#3�9ǃ�j�٘�S�7�0�I� 
Y�d+�*�����,+�󿳥)yx�(^�+�������s���;m1��1�,��9ۛ���V�-$�9�,�G����=� 6�^u}r9	���9��p�@w}��.b�/K�[����"ʹ#�Ak�Ѱ����	z��%��I>*C,І#r�
Z�`�)EQZ�`���� ���aY�g	r�d�$�b����j��i��O)ݨQ�� ���P�y ��Ö�El�i���9��l��Վ�e'pf����S�h��i_�
��G4V��k��~�ݟ&��T�6��d���(��&~��I��p���D��+���VE&�Y"�-����lf�#�}?Ȋ��!IV�P|�N���W�a��N=5�$$�e#=C�L7G��6z@�xP����w��mni�ŰG��ښZ�Z��U����ŀ�)�.<�/����N`� f�aV���{s!�ǃeN����Em��nǣ��K��@�*����l�n��`{�j��۸��$oP�5˝�h��S�6�Ƒ +(S�+`V��x��cJ�
�>/8*���j���u�֑��"�3�ai���/'�