��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`����8
�2���:����m��Y���8E8�mc�`�#|�R\l����弐NҤoe�����ja��~���	�X�]c=��(�,W��~B��sTs�:���0�#�t R���A�s��17U��?��+���!�@���T,�ȱKG���RS��OpL6!ףPQԹ�s����Y($��Ж@��;NM�i�o!X1�B��� ��w����?�M7�U�
�a�=hQ)F.x�i��v��R�B������wa;��b�>!�w�뿏⍹s`�KCui����]����31��өB�;~�&�p�\�X������S�+o��84��X?*OZ��l�Tc7l��Ń���^�L����2)$t�z�4��F�4������קu�CEV��Z�,�U�}-UMx9�#�@u�k=DN��2>��R��ļVh�}ĥ4��?'��Wd��2���2~@��hU�#u9��:�3�q-㼎]^:�j/��Y�%��Z�/�u{���f���dns�,0�EfTO�%:��!g�E}���L֔fX��_��i,ε����/����mӌ�_�_a���L����W�y��~�.����ăA��5w�_�$^|�}��������lB�Q�o��}�A~�(�##n���8���q����ɘ���5τ�}O(f�-�1~$B;%�-N��D�凧}0�Fy�"��l��H?����
�yL�9�i�*�ԛ��XS ���m�1�g�&FX���_4~�b��aU[�.8nh�0�\F����C�	�ls�*�������q>G����$�J�5�,Ͱw�̴4�ld�	�=�| :�z�P+�xq����Wb(ڽ�L��+�T�QԈOs*��l�a�v���F0n+�^����y85'�G��ڡ��ݤ�>a��>�����bb�j�b�ά�E;�����	Z��y�21�vnE��ή?��PD���|xv۪)�c����̙��x�.��BC���о�T��ھ�M��rꞓ<�	���L��l�ꊂ�����LZ�J������i_d��X�1�l3� :���Y"�����ił����	M�x?@?��~c��,!����f!��e�_�u�N�qX0�߶�u^�(�<ܖ��3�O��Oo!�1�λ���B�U�{P�&zƎ����	� {�돈��3�2O�y����XK?ȽN�[��o$���eҒ\��dV�K��q��όsw�o�ٙ�
��q�E��,/�]h�3���4+�t:����������^�R�)�甡E�Bt�E�!�(��5�MP9s��Qo�T���� �R�aM+6^�2���u�f��׎D;ꑃˈ[�p2QϘ��z4�Gel���<Y���"��	���E��>7�!�,�u�!��w�"��2��)����k�U-�l�r��瓕j����S��9N���!8aͩ6U�}=���7�z���^� ��O�uc����6�GF��gs�OB����f�u���?AO�E���R��J�
����:x�[��Ӣ�(C`+�o�Wa`�=��|K�H�����Ƅ����N畗>2_�TG��3���+m7~�ގ�%��+�N��g`���IO�1|L�~��*h��,������ܝN��E?B+,`�@ˍ_�4ŠPRA[F\r�B^��T�������m�c�kC0N��Sm�[٦��3�"w<e��gdgLi��� `_���4�s���&8��\����	���"Q���)|ʶW��p��\����H�a�E}�i��[��'���tE��T=�ȼ�F
��g���m�TQ7_A���+�5`YNڬ�������zES%���T�zRX��7���*J���ѐ@�k�GZ��O��%IT:ӓ۞�H�I�a���R8@p�i�=��Ӱ��@E��/�^� "2�M$����]x�a�E�����ҁĲ�7kfDۭ�T���c�~�)�����"b�����^�����3ķw�e
w��f �s� ��-1kk0�U+���� ��	��G�V�/WW^ڄvW:�x�#!Ѩb��d���%S�:��6�/\��`�=$eM�+Ra|5��
5�ɠ�B�gQ�M-M*��fc�-	g��E���G.W�>�x�c щz�Н��W[�'IA7�w�D�)�䀍�Z7�d5 �]��v�)E�+���Q.��#����n2���"b���6W�d>G,l�-9�6���c^J��!s����v]�c�%��_���ŐEW�f�-v���:��}*�%|T����ՠO���G�zC��D��>}Kt:s�a� ���%&�} �Hh�r��mM��t�UEݦ|.���s\��>{�*V����4a��.\l���R��p;�A�-Tٮ']�պ���N`R�l��Uż$I�����I����Ӗd���(I�::!m$�L�*p�I�&*�w��d�7��MKX����&9���y
�3�F1䃷��ӡ��-�.��t�50l0t�H�bH�^?a6}����7�os�<vBa���V#���P�N�3]ч������Kw���aX��xg1�w
��	��+�H<G}�����YZ�����b͍�'ªx�2���D/O7�?X�"27�����J��6�xR�pZ�.������T��`��&Ҁ�N� ����������iG�����T��1� ^i��R��=����E�T�����%���u���aQ�v%�fW'A~ѹʳ��q� 1�~v���WÝ��itC<A�%*�@y�1�i��@t����]�:�U����Gc)�}}���\������4�s@�n�CG�~�@��^b �Y���H6�U�0��Q�����F�vir�k��]��0�/��p�aW��u�U�Ւ�2O	���ظ��T?�k#E

�} ��җ�7���+5Z�N^���,fDn>��6)|@M�m�o�Y��<Uz�S���u���S�����l������QĖ9 ���j
�ӄ���8���K�M�N��o4s�DP����V�p�4��,�Wϐ�\^�-��$C �jmŇ%�:��PY_���̍ROC�4�{|�!Q
-8.a(T/moU�3��V�����q3��_��3Њ@���QQ��:�nq�g�~?�M'H�)"-G_�|������i�a^|�6}�z�J�
$nXXH��g����~���ػ�ڛ27gRa��Q� �lY۫I����y���
��*|z�I�{^@���#�D��-i�i�Q����*����[�+�z�ƈ��{��w@�9�`)&�V�@�ݟN8�=J����n{�ڍ���Q^���^�,��д�x�p����ǩ;�E��]��ۉ�;��>b������0*��o�O�Zۘ1^�DN +�b�
����O������ I��)O���9D�ק��=@�T-js��kr^�fjʠ*�����_:{+.>�� ]��n��L����|�I��v�w������a9&�F��#U���t!wޢBO,2|o�!�)��43'�3rq����1�%�#HE��wڜ�(�L�w�=�S���@Jo2}�wJ�<�i�H�;J��j��|�y`xb:\�
�ŋ?�^�l�T�vP�f�(�iRq\?� N��Ɍ}�c��e���oT� ln��)�a>6K��Uh����ǫ�jD��% Q<Y;9��|���F,�_o��~��\���
�Ն�����k��E��<���;���U4�<�
��_���.Ҟ�&;��X�>����C�
��Z�nj+W㺆j���(�����)��ዣ��/ܮH'�'��м~-hIʗ̔
v��n��yD�ق�.�����E4
E����\��Z%\~c�,���'JzMsz�_YIL�$�-�d,�8ϋ ��b�x��SP�2�� �J���W�c�A$x�L0�|n��|](<`�٣�~���2e蚌.B-Q�?�����F�!őo:o~i�.����+��J7fH�r�$�伪�:]�i����͔4 LQAl��z+E:��O�Y��^��7��� l�F&��~�c~h��H�x�S��Q ����w�]���E�Ȭ3��O;���O`���"$����oA�ˁ�ڑ���&��Ķ�_4��g�9]������ ��#]�T3�p�}�_��6w�(��C|����m�t����Y_�u��76��E�N/�!B:�|�5P�/TF�$4����M�>p���쎁�mY�� 5��A�#��/�c�8
|�<N�Uq�h�+;3���b����V���cu"��B�j�B�]���=}�z(��X��"�5���V�F��~���[g�'Kv�N��'�K����c�
r�
�Pv5ٱ�q��SJ�ZcI]�Q�8��𯩦aB��ww�����e�I������9�rݥv��C��7$t�2���z9]*��bM��|������鑥t����V7
�-X=Eb�_:���i��d_��`�S��I���V@�<k`Q�-c�5�����5���Y�y��/����kh05ӡ�\kX���<ȤRYl4����D!��"�5{0e��O*ߝ��({-Bdg�ꙙ\�ȡݵa+R�>��0~��T� �8mM��r�b�1 �ƨ1P�K'�� �\�%�ۢQd1u��=�d�i/��o�r���GHM�Ҭ��Q}��MA-��0Fqӑ
 �����V��RP�GZ�}5�e,;=��GT�4LJ��N�4��ۡ�K��Hn�~=LE8�R<��;�b �kf0��E��5�޸n�"���� �r�BK���[9�z��(`�nH[�C�Z?�C�k
�\[�	gϠ+�QFb3L<ͨ���
�Ч��*!
�6���4����������"��\�#���/GG��5c枊��)f������a&�E �-��K-�c����8ke�ɝ� ���NH!���H|yF)���sjLf����w���l��JN�#�p�c�XW������h�	/B?�N��kh=iĎ����|F�){���iN���j�QM���'�Iڮ_��V����x�N��7wts��� �C"9]�u;g2H�C��r�iR�yT�l���%zg�l�����NI��l`����#�
�����L��^1|j��#$�����Q9p?��f|�2����C_�J���л� �����dn�������y,K�M��H��{��������m�W���b�y�(���3���}���c�ʎl!W5%IVe���{��4einu� "bY]����ŋ�(TΨ8�{76����o�ֆ���	���z;��ې�~���C7��@><o�#.b����D�bNn�s��T�I�-�d��.XL�FH(��r"=B�TM\�s����R���V1�l/�3}��N�jw��Ɨ��Iq�(4z�۞�S�nF8��6<������x:+�yx��OP��I~5�nңKNx�W��΄	�my�^�����^r��U$j��	��ؿ��ݤZ�+�������s6���fH��9>�<��_b�D�fN��9|�w�n@��q�+rG+Z��12���rF����M����PP�;�B��>?L�u�:�m�j;�|�J+v���|���z��2���}iל��:��{i�����Zn�nj��v�8ٌ-r�����#��-Q�ʤ�+�t���6�ҭ&T���5?�ߌk��vhd��5�� ���<��x^�W5i:�
T>~|�gC��+E.�V��	&�O��+F+�#�������˩
&���Z���},+�y瓷��Γ<b�KV��!��ݟ��$����}�XBQ�Y���]l�y���Q�p�&d��[u6>��<������a�Ya�ǡ�IK�3��	��UX���G��St
�{Mno��; xY+����� �}y�L�ڎ���Xt+�ڧ��-�m7��SC01Kq�?M�m�lsʀ�5��i�Y��$"]��O�vȌ�I�+��s���0��$X�M�
���:��m{�RXlv��9������_�:�I�@����D[7o1��Ԅ�4�*]�q��`���j�U�V��Mp�l)\�#���H��/g�<P�=���'
�*���坛��/��Z�C��tlS�诒Ps�?�O��U��'�j�r��GT�D��tٵ��oq�h.A�O%L�o�P�ٛ�.|r,j�B�B>S{]Y�ŚŸ�fE�ge\@�$k���TA�}�#Ƅ���ʬ��W`w Z��f���q3���A5\����_�%�h��i�]ȝ�;�v�9w�8��\���C�O\i�V���|8t:(�X��4����yy��ު륰E.�zs�Q�/���)M8}�!�_��՗>��/��@Ν5k[7��7�c�Qj�rlY��fC\�x�"_�Z�$5\�t�Mo	I�T���k�Y=�7���-S�T���؊�4�+�M�gG���Q�P�a��&�����w���KP�c��L;�ֆ��׬Y@�6\�ٰ���
��YO�_d�lPG�3R�Ԃ�*j�'����勅�",Z;;��)Rkd
�Y	�L�:�Q"'��o��v8�T�$� ~�w��9�����#��\g����.�R9_����	Ͻz�Y��8��j�}L�5k��2������Ee}���c��9	�2���y�N�_��3�?{7���F_��ix�C��{_�h� aT�AW�0��' a-Sk �!���=q ���>_E3M���>�K�4jM��S1J6� >'�?�|V}�ˊ痧�-������F�Ֆ<w�sx�k��I� �[ܶ�D��P�~�Uݦ��ٷ��P܎�V��!<D��>��!l�I���`�*n�3�����+yYT�g��%�Y��H-~L[*�a?z +:Z��W�@"��W=�Ͱeĵ��#���v�Ÿ�N5�AI8�������H'�F]������y��b.(���e�.�ӫ*�Tr�`L�3��Z�[� � kU���RM�������j��r+"X����b�����
@�>QjE�Ku�w����t}.'?��������\:��Ĕ���w�>*��n�NU��$��d�ݖ�GQ�B��83~L��y`9Px ��.��V��!���i��(��5���3�XR�;:xyX�K����h!d?�YG��L�$�Y(�'���}�u�viT�����)����dk��Fk)8|�Y��}�X}x���Ĳ8
v=��s��૱%��h/�P%Qh8�j�>`����h�wY�j�v^n�Y!�<��V�S"hT2��I6�%���8ZY�*�L��Dt�@�N$���G�����	>5�]��4�E�?�mN|_$�<��\�3G�L���p�p� xX��7B���/av�?��*T#_2YX�Pm���a�ݬo<�q��VV�V��T���a����o��F���a�5�(�A؁r��S?ؼ��2B�d]F�����e��v&3H	.�ӎ�GwB�l��UMS�r ��"��)m��8L%`�C��rC�Z)#*����ޣ�vz��D����.}�����T0����CB.)D��-�l��Fk��om���H,ώ��NV��w�L���#8u����η�DB5��q���pE�GoA�	��H�C�GTp�%,p��ਜ�r¯J�2��w�O���	Η@���y&=��A�[�Lc9
��X��&���U�M�ž"|?l�a<n��̯G�)�?�P��q���ߗD�e�10�<Ȟ�ۣ3tT�R���<t���+v/tFfk����
I�9�������/`#�n�!�}a��0.iX���s>@��`tT�&�i���t��Chqq��.6lL���4��쓚��K6$��hpR�� ��kJf �ԼH�>)N�mZ`{�ph3���`{���n�`�S2� ��L���%�_�e�Ǭ�^���Űe�}�2�� �����d
�y�����P�4���T&���q7�#�����	�� ���5A:0Լ��/����{,d�Ji����G�{}6e,@�㧳u�·�(k���@(GS�@��}�����pljtW������>Ԣ\����*�	~��ei�ڲu݀�x��U�޸��ߥ5b�����n�ݴ'��}{�\�� �ð�u%�2���q��cN>4���9���Zv�ʶ"��tm�~;���A�)�e�4���l��n�3=�T9�@㳃��[���OՌ�X���%j�&����أK�ᕯ�~�]}w5�Z�c��@�2��_cLh�nq�F�^l��-<L��U�#jJ�J�푮 �u�8j��M:.� ��X�&�j#���R������Pl�j��ǯ����z���W�o�2��z���X��[�qfӛXP ,�sO�Ԑ��d��,�H��p'�t���σ����T�{�8�����ڵ�K�3
���j�޺�ְq*j���|<C!w%p��''��+1�eI�Ry��KMi���o��,��<�9$q�K���:BR"W��(�H�<�Q�6ōV��3>p����{��w`FW/a�UĞ@�sv�r'7� �=z"Ttw�[��d+MI��{�� �9��'���pԺy�b�"��}gvWkOK�nu�/2v�W����M^�7n�,�>�Y���:�e��Qg��/�[.��X�N	|ߓN�,�kٞ�L��W�w&�v4󇈭}�
�0ڧ�7��a�e��1�e��|:H�T�|�A��4����	����K��@�1��o_��mo��"=j�-LT�0<#[>�}�����F2�>_���ޟ��1�';V�㔐���X��g���S�h��8P��^��$Ir�g^i�g��P	�V�܅��c����L7N��6�1��
F}�0�fD$���L�H��ޡ�s/'m�U"̂�d��=��)\0�U��!k��.�t��$5.R�K �N>1����k� ��,����t�fhh��L�R��gt�f>�1J���!Fk�)�BSd(�h&�~O�]��$�y��NIM6�ܼE<��1"V]Kmv���DA-��D��Ku#c�t%��R�,�i�ЯM�� k���$�yʈ�4Mm��e�a(oM�� 4sˆ�2GVJZ��[���v*�?���8&,NR������={7a☚���va����(��Hdh!��A��0��{4P!�Ծ��C85�וug���L��RJ���ZE�W(�|G���h���Њy�̴,��%��,����v$w��c�ǅ�k$�@�3>T����%�kS=��.c��I��k`yA̫�Z�d�:�/���)��!';/4�G��uN��9wz�������̘;� h
NNHk]q=9�Ӌu�R�5�Y+/j�2��?�^��+ԁ���E1 V �k.Y�r�7ҡ�`�I�e�ud>kTw����i��C"1��n �os����n� o���jj�-�Z2V�O���o�[�0J|	��t/���&Uu����i�j��'��� ���F�?4���E2�ݓ���S���Pv��XW� �vi�<og�"ݫ��'U�E����m�����1j"��*|E����CZ?����jgZA�nn.K��e=F\Bj��/Z�|�|�����Zn�CG/�uj��qH�V-�wgOd�}1�e�p��i__�;u���DU3�/
 �����s439@?�W��_)��(,=VHWB��{��qP19pd�??-y.����+���kν�g]K�E�k�M��,��m_�Hpf�ׂŜ����5��+o�<��\0�j)�� �>�@���ɮ�W��x>{�����,���"g|��-�EH2���H���o�c���R��� �|���G��N�~o�?�gU|o�gi�����Pj?�337��F������e�^�Pa�Q�
�^����|�qLp��i�(�掂-Wg{9⢔5S�G���eO��C.S!��п�f}1��&�ׄ���_��8�Z�BK�=��W�(��\}�8S��KT|JU,��H�,�4,���P�)����(���+��AX:��'�/�%�</#c��,���k ��>���Z���F�
�x=��L5�.	3칍^�tO�t�����	�0 y�يl��<��Y���5��v r�*�|�Oy�ʽ�T]!K�����o�>Sp��H�D~�<K��جs5��Z�Q[�{�	L���;�qFV�^}�6S�oDSYÐT��t��O��z��@3�y���=ʅ��k�à�2��J���fk��X�$����o˧{I��m�7r2�+��aɻ'	K��Q�(b�W��"�NBH�fM[@��<���А��wC�&D[p�]��j�r�丳pU�{�774mZ¨h��6k���<K��v��IK~,��lB��aV��/qc0��/:#�׍����6�5���±��@�o�`�ǕK�w�����)�o
�]d��Qܢ�~Ws�wS��lz�5=Z�d�c��pɤ��"E>zVʊ�VE�(�k�C��A>�G%��^�z�ɩ
,�Ѡ�N��O���A1��2�ۓ�nn,%� �q|�(�@n��%2񵛮��Rϙ�N!�S��66���s0�zCN������r�`?lXB=�a�p�ҩE�6d�����n�t�#��3<� ����Xi�Ui�JeQ����k���z�q#�Rh> �N1Ʃ��W��j�F�b�Y�6g%6�[.0n@��>v鰉{��Y����|�p�y.S2�oD�J���$�sz��j<3lL�5x�&�͌4��gI�+p8� գ�2�z�G��.ȡ�8�|L"p˳s7����rǰ�N�b�+��*0��;�C��y��F6��mFy�4g�s�)�;�+[<2���E(�=���g\�1k�A���m_Ö�BN���dðd�[�2P�v<�\z�*�鼤' ݤ�8�Ίީʟ���C|��:����������R^�}h�,�"���]�{�9�C�;�z�jD�� ���k��۬ւ��o@w[v�)v�P�lW����CC����z�?�5�J�5�jl��[�+�<�g��՚�g�?�K
���4sm����ų�ʯ�8VZ��(w��!|M�<1�	�|\x[���@��lT��u�V]�t>�m�[Ĉ �� �>g�m��Yy����D*v4෡�D>��s>&s=L*��+��/��~�W)U`~�z������-��]��[��5U�g�K׶'8D���?ͫg�
H,_��v���k{�vC��p$�C�es*���� �Cdݕ�Jb*�Z��x�Q�C\yU�Q�Co��/�19����<m���?�E_1I@u5����VL�,��"�����������S������|�"mv1���^����vlɚ�3�y;���<�Ќ7:~�a g��f����{�!��:��F	��smQ�w���`�� F@��%7�5DN�C��Ŗ��3��oZ ����>��g�̣M��(���B9Z�ڈ��WK���N��FYu��&��N�@m+=\Y�\TW�nSBd�n\�-�������蔷���O���'��kq��}��@���c@sU(�=M��\Z�s1Fn1��'6�l%O8�ܨw������0��v��Ƕ�ۦ���{$h��;�������9X�ʱ��$�u�d�k-F�<´ �4��V��$&������w���|�d�'��xB1��_HYNF	���\���\���i�F���r�T�����ѧ�J��$�<U��--���h����0��*����T�&ϣ����,m��c�R��%�Z��.�Y%�{��p�(��&7%'�<I�r	a����*�'�D�+���7�	G$�ՠG�@�wFc�t���0�}�6➃����y��_
������0^勸eh&쁔���;��hY� Kpw�/Fԝ�G��7�/�s��٭�nU�5����
N3�5T�[�[Ē��O���1�5`+�NjY���S8�1�^���̲Q��7��=p'
�� VPB�<]�أA,(����D�?�P���a������:�)"͌��1jn�*�]V/��Rz��wΌ�F��������e,�A
M�q�����n�0)����|�^�"*�L Q�z���xr#����]����+/��o��)*���z��53��7)�:���gIF!0��������o�����P�i�rD�
%K��JH��r��kM��_g���5P?�܍8�~�+_�&�@�0?��-0��ƭ�j(�R��]�nm��X���x�8���"�:!3��L�NB�����{I��~9Cn˻�3��O��Z�>А��Z�-��7��SR��
Y^m�ov��3T�w�����	�yJ�AO�[+&�>@*��C%E'�?Hq���E�-��#���O�0m�"�~�T�X}�wϜ|åT^�f@<�9��n��~.%�lF�"01�(��@͕-�D��8��-�Mo]Ĭ�r�}x;�EK��@��8.��a�A�i�0�a��T8�w�}�M���} ��wRV�N�ױUP�,\�A���6A�p�T�K" � M�w�)�ٝϹ��H�����eu?&J1�/PU�h�a~�Љ~��o1g�IqD�Q@7� "b!Lcy] m�aq��<,Aʋ�o.�ޓ�E�6��!]�K<�8^3*���ͫ��@��fjӴ�n�a6��� V%(�ܗ�NA�qJ��� KB�����7�Ɍ�Z�y8&&��%z������4��>c�fy�U=V�iW.:x�" ��z�%�_B-_N_K���E;�2�O~Cnxa�{u����mĝ����p[�H��Z�����n���&k�3����K!�GB�xs��q��[D2�aJ�����r{��O���@d!?(�������k`���h��^cp�l���@Ҥ�ǵ�vo>sS`y�;D���ZΉ��;��>6��ErU�[��8��W�܊�OXT��5ě�Z4�;a��Yv^[��~�(P�N�P�cKz�m�jH�n�Ο[o��P����([u�\}.b��E�����<L�{e�;R�v��
R@?��H#��Z��QA���/�+��N��)Z���x�/d�t��'����kv�59���8�H��jE�Āh]�"�C�Y!_��$�-6#�I��9?XRx�")��uit�F#��{D.���:r�.8-XP:�ù�0s��o!MD�X/��9�t:��-m��Y'�n�LT�|����1�<�����Nq�CuB+�<�j%6T�M�/�^r�'��m�!��R}�y�	,����H�x���<��\���pV#�����{oU�-��I}�I,-ڛ�pZ��}�L��VS��� �Ej毱x��KuA�#�8��͕�g����=4�|ֻ�jR&K-��H��sW[�8;�R�O��֏J���$p
:%�}��햗r��S}+�+R<�\E�n�LnH��iY~��[�(,S�TC	��ph@"��iUO��.x����A�B�����{�U~�5�4A<�1� �gǭj���R�f,"���d��3�gֻ}�����o�`8�?�3���R o��wO��p}{���'���5�,G~}o��unZp&�����h�����P�t����3�9K��Cj#���q]}>Z]d��D^F)����m�\p���~�f���y�WL��E%�w gw��!��"z�9���'�{8*?@�QO,p�������!�-���K����6��H�����i�X����p��"����9
��ݦ&5r��]�:�s�x���V� p_�Tr*�N���B���;'��E����<�ex��y�8����(n~�@ި7u��rl�ß1���]V�V��9�J�Y�m�T��aY���E֥�M�b)�|��$�jA%H�R�T�̃���pe7�O�Y;����l�� �����/�[�:e�*��M����Hf
��� `m�@^�v~o1�ɨ�l�$��Q7�H-�n�-Z���n?MR�DA���{���Ո�f���Q�=«]��5Y�3d��
��Dг��Z��E�����pi�+|%�1�i�-�~�X8󁷉l��Դ���y��}�F{2��H��1��U�"����Le�E�j#��6�{S�XK��*�0�N���"�4y�0�N���<��\���lX+��m���Bd�D�� :��|w�@yd���P�t����ǷQ�D�1r�>�"������^Jc����A���e��Ĥ�m���,���=ގ���x:�ڳ$k�4:��X*ըz�c1�U��L�pQǖ�#)�ظ��s<h�
���x�|��>
O?_���T�ϻe��D��c�y�6g^0n{Q.�n؅�<$1��������:UXPi}:91J�Z1<x"��X�ö�r�3�[Ꞡu�kKQ��q��JhƏ�W�w<�aifQ��-a�:P��el�!�m���js��_T0��s��p�o/ca��u�2�Y,L���S���UL8D���ڻ��I���G�A��:��$��V@�y�7{ݐ��:��Hn�'%��W�S17
�'�ƞG��|c������u��WYN����&����:S�K�
'b��Ac�bX�IаO#1��)N��{s�fV
�|�=gz�C,--���P����`)�&s��łԀ���.$�M@/�V���i׳[K�
}M��L��S���)��hX�uĂl�	lo�ױ���hE��~6���E;;|����|)!�؞�zi��]%�,�z�H{&?P�1"�!�W��ο�r����\pf��=CG�3���GC�ӑn�p�5Sh��-w�Yb/Q r@Fsy��4�{i,U?jA�G��/�[���3@X32�p10j�#-��8sC�b�۲G�Qw�6A������k��9��v��W�; ���l#��T�����>�;z�s>W�释���a}�3<��;�oR̿m���a��؍�co
��ׄ��yc����T�����1�_���Q/զH~u"=K?�Vm�)��z��#*�A�Lh�����0ώ:����wu��� �S�ð����X�>�SPzB8d�率��?�X}���~�y��0>s��M5ɨ|#� �3d��ťL�2���_m;9���Ӈ�k�OV�1�9�6W�:B��b�Z����6J1] �%kYꄑ�6u��;Wy_oK���}���?)�_O�J��*�O{��P��17C؅{6I]�.��V<Б�J�y�F��}u�|Ń._(m�{Ӿp>�B(�;�r�>�>�u��"8���L��rx�n��̡�,�s���������/? B[^
T*�ݦ�R�����[��걱�������%xeATb��FʀP�6�n�� ���7ZqO����)�=�0�����<1��Q�d��+�~�X�&]�����l�C��u=�MV�������!�$�ՀM��|���n�~��dUX��@�t�c,�I.S���/�emz��Bp�rE�Y;:&��B����H]ތ�<i:�IwSyZ���1k	��iz-D�aE����$}�� ���4[k�
����W�v����v��l=p1yHw*sO>�"l
�hu\$6�OzWh�8ղaԕ����Ȋf�ͽas�1 ?�^]&]��_nseB�yјMr[]1kb��nZ\��<ZG�ĒI��@��!`�*/>H��	��	��>�ktqm�_A�������p,�SӞ���CN�Ī,�4�O�#��0 FL���|�m4�����ߛ�N��	e�p�/	k�� �1�o��ǂT})t��f�����9}�
�E��+�蹨`�k�4��Ik�@zR}1�
�
�u����,��.B��5�_���2f�g���l�,H���G�3"���j� ����
��a7��7!N6?�N3��M�� ;�/�Ȼ����-��x�٫��|�?[����KB�>��:hц�%��5r���t6i�;}J�sQu�>Q`yD
��_���pd�X��[��gH#-���ku&3��#ce��7�yK��6�O���S�`��Ar�r�J�>�x�CK�4�?o �fsOF�Bcg�)!��Y���1�ƍ�_�iI�˙#	S�g���Aw�ZV��	�	�9F\Gauc�iC\�A�	���2H����}\w�H���6E�����7��z|2j$��xʔZUowa�2@+!^ݨ�}~Q΢*�Zg4QP_���'�R��� .ŝ5}!����֠U���ҟ,�S��(d^�[l_�~�H��٤r�LF��wy'�I�R���u}�6Q����t���Ύ�����?�ݣ�/�b��ʥ��
(K�D�6�Fb�)֑(7�����c�0����b�Y�Ǆ��DG�Zhb�N*���{�l;�����(�b~�v�J������;{����_-��aU��_~���7ì�j�x�@6;��C����:H�ё�=�wă��W{1m=�5گƵR����Z�y�瀢r�.��s����G�#ӽ�lu=�;�o����p��!�A����/.���I�z���Aq?�rIU�3��y�2MI