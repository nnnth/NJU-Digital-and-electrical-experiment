��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�x}��j��S�b_�)F�1�(d'Â,L.��ꙺ��e�˭'�{���)�Ilf\�@,�y��Z�n�X�D�P��c�����=���]Od�w��yD.΃��o�%���ƪ�1�ޠ>����&�t&�n�E��Y7<?.G4a;�_���y�_,�7G�n���j�H3�l��2�� ����^���^���C�AB��w��D�� A4���TU-��/(�����j��i7OQ�1$'���;6�q�4X��"�V�S@��ʹ����"�;K9�1��f�V<���=�\���'��I���1�g���4~gv���;�.YI՘�V.Oz6���7��>�Rr�<����#K��29���flfD�*����uf�0FE9�R%������9X\ȿW�}d�
$hX~���q��I%��iD}�Y:5��b���H�=��N,=�
l=r@A	�o� �a�m�!,79MF�:������K��?1�ȼ@m"�� M��F��"�J�P����i���5��c"a�Ҝ����)?w��uUW�EM�&?�©b~V��5�^t��� HSz�-���sƙ��źeXԁ^׬*�ڄ���TY&`RЂPj��y+vj,L_����Q�:�֕��8q4�����JZ1xaU�"�0>,�쯶�}N���H �X�Gy%(�
!A�~�N��.Y��:
�s��7��1m�hm��~W�K��Hw��*�vт���d�<r��W9
qi#XŌ�Pp4�8��A
�-�X���!N�oWNB�6X���npy�������J��S"Fs�����P>��WL��āϟ-����9;��y������Lx�0S�IH&�DƁ�y�6�hK2
��L�jV`��Kr�lR|y\�CR��/DT�߬�M�eN+����GjStc�����w��-f�W�#�����f��Ӿ�Ƙ8Y+1�P���%[����}�afx��� ���w"�ڈ�8��b+������^�^qK���oY}ҁ���Ĵw�[�p�6��S�*P�ܻh�J��y��	 W/p1d�"��PK�C�Z��e��H$��1ߴ��_ˡv�p��;��Jxܵ�bRզ3ay�PF ����N�=wo]Ȗ�z��I�~��� Z��	5)U�W>���W�4[�T9�p��n��>�������k�M�؛�3{3	�|aw�	�Rq9�k%�Qc�W�l)�8%
c�{ń��v��-��%)nnc�<����]�	�1��9Z������Rpa�eZ�a�9��gGS�t�5z��\�s����q?�^���q8��u�L���i�?���nB�NΪ�<N*�7�LK�.�{h��h{B���RH�A��Ci^Z)��eD8m�՜;.�1��_4X_�͵�Ϟ�L�3��!��z�sg׎��I>^�nK�Ѻ8q]�u�W�-Aw����y��l�L�sf5+��e�T/�z�����}E�g�o���Cp��L�BF%,�@Hf�����_V��C|�����GHԉ5}Y�:F��䦚t>��8�T��Ɏme�q����m��uS堫�U �,�3L�L	��=�Dg|���@6�%���uc�92�"X5�B��¼�4G�HIV#r,Wo�I�n�v�9gWQAkp\d�}\������m�߹�-��p��T3n����cs`@A�ڡk������ԑ���W�JO�4�(��"�D�*x�a� �H�r�V^D�Ւt���'�����|̩������q oo��	�>"�A�*���tK�������L��6H`��!N|��0tXT�}�����Ȑ�W�xE����c�mvſ��{���V�|�F���6������&;�Gv�(�sjM�.�dx�`x�91_�MfO%�M؂�U�2*��._�$���_W�J��S�Hg�d�񶦼�ޭ�ϛ$(�(wqC�n����	����W"�+&�;:\�}�a3A|"�c��t$��)?��`�4��*����T�^���g�G�S���A�P�lh��b+31�
���K�D�L?!�ˠ@��)����k���C�F1���k'm�;ON�)��R��k��MG�,�����*UM�?��7Hۑ���6ٌ+��z���`_r�]zĽF{{�8�]��� e~j\�����4nB�����S,��*�%�	���[}O�{y3;�p�LU�(��V���Svx?���H�?"�{z��F��K�A��))��bW�s7VF1���6L�����=��6bA:L:��cv�&:V��;�ʹ��ÀH���R��j%��F��wy��X)T�B���3'|mx2Z��M��6Қ���)L��
.�7,�,ɵ�6�6Õ�hlp�ZBS_$[�fSCټ��}Z�����f�_"�	?O�{{3CQ_�Ŝ~�#^�L���idmQe�n�����G�Y_��*�9��+MUz�.ׇ{�=���|D]��l��y���A���QVS�GD�[���J�J`�x�P�=�LK�=Bp�G���K�@� ��ٽ��I/��>�6N>����M�n�#s��`a=FU�ύ�iW��іusC���G�j�g����؋�FgQ1�D�r �f߸C���T֓-y�h"�*�b�;L����`������TҜ�R���tq���- Y2�1��qOkh�
��P��h��PVy|,�P�iV��4's��2C�]�Lr	cy�nmKd�
��;J���1�����K����
�T�ķtz������<��P��2O�ף��T7-#��7?@e�9�־�)	�W�k$9fb����6Z�تa����'�]2N���Q�����>_<����6��<��i��V��O�QO��*Z9�3 R�>�*�!EGZN���)�,���<Qd�qpC.���v�����\�4*�8o�zV!Ym�����S8.��]�^�f����8�&�w$�^;�G~�U��7@�zb}����q7�X����bI�!H/�����4����s����j$�R x�}W�>���=,��Ka�2I����1�W�}��"�S3��)�d�ϴ�`Ǩ�1w/�>p�,;2�5��wL�����g۷��f�J��'+�l��J��Z������.%� ^�̟탻�8h�#U�!�x�w�-GR|�3����D],�S9Ѧ2$�ݙ�uɲj|y�b]V�2�o_��.7��m���&~7�r�ΓJ><YY_��j&���q�d��XT����h%��ֳ��Q���=K��:��(mY���"��7Ģ�Q8E���~��V�zv3�����ĵ����#`�|�/�YK�'@hiR+�͍�}-k?�n��W��n����_6]m&B-s�wWN.,h?��ID ��Ѫ�,�fǵr׾�-�7�h2�,��S�P��dFˑ�H�e�'�n�'u�Eg�
djE���6_I�_�BxgW���p~�m8���֣�!��>US�%�����Ab����SV�`�joEE�v/��J��+kNU�ز�
�X�]_>z�;�r0f��Ղ[�/V?E߂����2�H{6� ��� xP9\���-�����#�U:��Iu��l���h��U�b]�C�8s7d��E?�����g�\�f6檭)ӀY��/9˝���9�5�F*P:-,
�s|Z��Z�.��xn�I��+����~�欃������4>��(~�nq1����o|�;k���5 �Rc�P�h�'hP���Z�����a�(�X��\� ��^���ɳ�QٖfM"_��ԑ�`'�9�-��i��O�@o����-!����x�b���&�������pĲ�f�W���Ly��> a)=Lrb��O�^�w�3�ԡ�e`lk���.�y���'��G�gg���D=�;^n/D1�.��B.V�WȽ]?.Y�x�|YT�E��w��NPIʨ�R˓���,={#�D����X7�0B|/��uAE,)-�jp����L��{�֌;��� �+	�l�7
���P"l�e�"��������p���?�'��G/���������66prnvw���A��rl܋��v��ٖ���;�@U�	���U���r� g���&�/P[��UV��/��C:��g��g��5
���
�zi���B�l��[���wO$�{�Q��@�v��Zaᅲ�&E�!kǂd�G
ӻ�E�L4V��$M�{R��3�a'�VRfw���/nq�J\?��l��#�>�N&�5�~@�܍��I�����p�#����O�s	rdvzs�+N�XK%Cn�"}��~��3�?�U",�ݲ���}{		B|'�@aSW��P�^U�o1�ҳ�ҊOKE�tm�����Q܇� U��(Ŕ�wx>���Lz�@�j��ۜOI�&��1�wh��fWj�B��},[�b~=Ԙ���;#���i�4:�\�c��,��a�>�qi,h�L�����f������y��8p����h6f:{S������R�2�&.����/��b��N��?ĀeK� 	ɩ6�m��{�l�|�|�9b�*1fM��C�N�a��5��!�ێ1;����9A${�`����)�P�{�8"�j���W�#�k6�[���s�*���no�]ö�c��/!�պ��z1E�{�г�b�{��k7��!���a�LVW�
��$�3��i:W��`��z��ȩ�W�7l�m�K���^}{-��/�M� ���r��3�
�H4Z*�* \�7Y]��3>��B���.�	#�u��{/�G'x]bP*��|'�;�;�S`�*�\���$A��n��H	`�C'|��O����u���m��C��<z������@k28-�
��U������+��p?5= 䟭��坋;�T[¿��7OM�x�W�om�['�������-���|����O��.�o>d�Xu�	�~�����������H�xfgeV8���p�-��G�W���7���
e�J2n����� ��g�a�R���	B�p�JKK"Tz����4<��HՀ��1�x@�r�8�������yt��kH�/N�_�|���f�%w��+��}���^A\���g�&���߮�1#X�jc��1���L#3܃*E���J�ݸ&���8-NS��B6d�K���=�d���!���f�j�`l�#�vA��tj2��84n�%��_CS	�+E؎8?.��':�lT��
9p�ꦎ�������.�g&�'Ie����A�T�ߗ�M؈Փ�������D��9tR�Z����J,>�ھF��$A��A���G�l��&�H�h� ����v���RL���yl�qYb ��i|��}��G��B��c��(��A�uy�
��:�����������L����c��\�Eӛg�O����<���v3��5X��t��ml�F���mAɲ�E	a:�D����|�c�6��/ � ��KJ&��`!���'�P7�,�(�BpV$E8=B�g��<�g�*m;�+��d�İ�?�(��_��]�r1=y�x�4��}��j�So=�^$�W&��R��Q/����*�9X��:��{��
����������}f�,܄`�x�:�)-Xg��ҕ�:�VT߻Y��2��4t��ot[���s}B���K��	���vܝ<���v�q����&*�0�t��a��z��<d����$&NҾx�[��כZ#@�đ~�7?�L���?�=���̹���I?n�s�*�"v�0�f��w%��L���X�X���kI����ÝRz��Ae/�=�s B)ޞ��qʒ_�x�7ڀ��tx��ѐ=��j8vШ���ћ�1m��<�P�O��g�+��gu��Lu���wD3Ad�P|����(5�ľ��$��˺T-�X�бk0fSzZ_�qD�ʄ�5��~�<߮�؇z$�Q/�J,\@������u�͋���@���'���te(cB3Q޲��$�An��b��v��EʉP�Bۓ�EÉ4��T�	ڨY���T�-� ��+�mB���7ɠ��+ċ3tj�ֈ��M�%�{�\SJX�_��5մ&�4���e�n���
u��|���zWR���LU^�_�*Qf�����f̲�,�������f�T�ݷ��˪x\RL���3G��܊H�l�,��CG�4���qh�G� ��x��s�q�V�vl�`7�p�׷u�\-������q�����s�����sp���Fn��r����N8Z�+��l4�b�/�|�=��Wy|\=��M�g`�E)�і�M|zz��ʾ�Up"|�gz�Ld;���?1X�)G~��t�E>e��R��p�?�=��Xi�H�I�Y����O-1G]��N
N��NeF��7<��K�TT:K��:�>��Pj?NHȮ[��!� |b&`�u���;��	\�tT��Ц�[����L�k�|3��P�N�,]>�����?��S����/I`*�*��ѥ�[i�5�2Wp��Z�qެ	1����I_�:�'.��.4�2�ϊ�Oڔ|�:WR-ʠs�=�/)�D�TI���B� ���>�T�y�U�G9vR��`\�UD�埖��j�,;�n#�ILˣ���i�dnB?���DA��'`P�W�\(㤷Pk�i���h�SJ=�N�>�d��VU�PV��kc��3j���a�>��H%l��'e3OK�"r��=Jg�'�zt��1���H�	��R�����bՇ�s���C�*H�Y���M%�ůln[�ܚIk[u�2Q���+=޷Vs��UYۊ����K��{� �u���R����ŵ��b�o�Ԁy����Y������:S�$<�	t���U<&�Usn���l��u��Jl̾�χ$`�(��Ԉ~)�:�Lp̭�t�=Y�e��U��ĕ�ah,�����,V��w����l���9c;8���^�DV5+6�%�\�H9��K�L��@�P݈t����v����qN�4��t�YF�S�ڱ٬M��n��4�j�k�����P%��W^�o�_H��o��%꽱�P'�JȜ/%/7�j���t��O)��l������׫�G���Q&� 6�,��V�$���
+vLY^}���HH:�f��h�����5�x�cqf ���gyz!�87�S�u��@p};�����+y;.�Hv���/��g�%����'�bٛ�%���Ya�S��b�t�MY�=�,wk@#�������c�!r�p���k����C��j]q�*�pm��g?uG´�s������A��bMP~�3'K�{7)��Nh�_e����&!����9e��?w���U��tdf�ȉ��ĕ)�t~�)�I_�|�<�?��2y��ad9�t� �cB�����8Uc1�oA%(�Ƹ�ZN�$F�;�*�B�9��S��|�>@�y{(������ uq�� �6�椀 s�<gP��*��ʲ��V"k�T��?��q���iN�?��H�$�z�gt�]��`+cLv^�b�yߣC6�fyʤ�1E���"i=��x�X��EXf|mC3 ��߫��BUҨ(8�:u�:ju�N��3����?(�p�U#u�*�W�O�/d��i1�����n�b�b���c�BPl�Ss��īEp��wع���b	ej²�)Q�mW"\G�YXx#�FKF,�(+Ce,��KN!'��
ua3��.l������:`>�T.*�brW�7���u�6�����&ؖ2UK������Z��UQ+�6�Son�e���A �ZN/x�s~���[c��m�;�(�D&!yY�@,ۧt����w$vK��|Z�c����� �Y�q�''�b����h4�<g�j�$��;B� WS=k�5�5ic6�+aeJ�yh,Nh�FmǄ��E����(-S��,E�Y,� ih���M�����P��1ɞ�5�p��t�E�1L�q�E(b��/�2�a��h��P���
�D�n�A6X6���̖��6�_�Tn����E{MȌ�-9pb�۱��0Ůf��]BT$��j���q��L�nʮ�ï{6�Q�^�gFn�	`����g���Q�C#g[���J�_��#fax���]S>4�O ���Ч6�:M��J��;t�%�ζ�UW�l\�(ZUL9�1b�b�v�S��h`�kH'��%��T�UXop�s���еZw"��ـ�7o�T}f}��xܔg3�W�<�͈n���b��o٫�'�����6�X�+�sLݱ�9�`l��>y�a0�?9���k�3��q��I-W���9&��� |��\�y��K�"S��K����7����J쁩��S�b�Ƙ[I\�� Z�+/f�����:ia]�GM��:�<�u~4:چ���/{������@��X-�H3X9g`�R�1M��N�db>��ø�d;�X�&��1f0�MZ�x#d2��@���n��t�x>b��7�f!��j3�����`|�����7�p�4m��+����a�wȏ�m�)� ɳ���/����&˳���x4f��Z���U�Cu+����<g��@��L!6B�Ie"yTG���Q��U�˅�������!�p��\\I�*=�Oa�����L�����n]�iV=$�@j�h���{�yE251�Y"��j�U9�{����p�)���bR	�=�נ�T���7�Y.��
Z���e�,��/ܥ�CG�'i,[y��rz����H8��u�,��?��XYS��LWᵾk�Q�j%��[ #����E��-�'Z]
����d���d�k��o�;An}$�	{�I�aW�t��}&`B7�j{aq�Le�Z ��o7y	U/HFo������ñ�+�(�)��lN�����2�/�(\a(YY*2�/G��?p<c�JJ%\�ɣ`�d'�:���~%4�s�9!k$�U:�:kO�G��a�N�s0�Ӷ	*fұ)�񿖮te����ӏ_�$f�H�;0���#=������TK	>���˔����"�ӳh�� ��N��a��-5��=gN��ٗ�*��m�{���S�v��O�,��>;;8����/y/^15�,�������1�mZ�)��up0�M����Yz���uI�<MPk���W��۲xfA}l�	V:����gb6�9KD!־֤�Nk�{(;���{��\�I]9Z��S�6eI^��/�w��]Zp�7� ��vUcLS������+r����h�.o�`i�Rv���1^�$ض'��A*6o����G�@�ԣ�/�q	nh�YiL+/1�����
,cz��U�!���覘��(���֡��_��8��6#�j�����K!������.��; �)VZ�&��y��gRa�M�´���#����i� ��� SG��7� �r�;5�6�������'M|��R��B�� N�Ae�bN�i�tu!�	�E�`�ֹ����D�B��$�l	�/��D�l�rȗ�j�>�>�Hx��3�6X�J�V�m2���f����r��!c������;k�����{yh� ���: dj�7
���,����u�j��Ɍ���
i�oӃkFe���Md�<IX��2���8g�0�Ny�a#k7�M*�#���/�)���1c���-��>���D���<�}pZN���naY�-�?�>����1����!;E^�$'��鐟��X4`�>�|^l���"w����j��.�X�wGb/�B�tgD0����\x�Y[Z�,8��V��p/���Hx����#��|�03]�? �/�_�p}������BgǪ�z��[�n�����h����K����Vc��/�8��lG�z��ty��v�]Sq���#�� ��_��v�(�e�m�d'�%�j�a�ׯ���>I<0h�V��q��6J�rOـ��|����p���h�rv�����UW����|C���ߵ�a�����c\e�_:8\&p=rni�Y�|	��)�Ȕ��e���Y��^4����⍅��uL}k,��EW�3S�G����Ma�����)���F�(�_�K㔢݆6�d\�ʯ��r����0���|�q���V��t����4�7��o^�{�D<���m�������{�{���So�D�����?��	z��se��~�������ƀݻ�T4>���� ʝ��
��0��BP���8z��ط��?ұz�ِ�(U��{}ߋ�I'ЙJNf������~,yΨ����[<T0��LJ���,{���-f���.U���I�?��*��L��3���l�@�6�9�	�y�O��|��n�r.C�G/�*�Kȝ�
�>�,qy�>Y)���N ;zF�V`��
��k�+�tQ�vvWu]6��0!��.��7�y��|��+4��l�l3�jU�¦��	*����T��?+�������p<�H��5�98A?z�-"U�v{ku��L2�0=���:JV`u�4�A���;v�	|��E��\����@Z���v�a��
�::5Ӏ|�g'y3���/��t���)��KB���Th4!�fG�	mz�ʥ������?_�rU�0'<���B�P"$��eV�-88�`1&����G��8p���@�(��-X�䯾 �V���t KGJJ�v��:N��I,�0��c��gؓ����(�W�n����<Q�V�e�»�=�)��
-}nr���k�r�C�%�� 0U+WZ����V�����T���B�y#a��b7�G�{kG�iB��6�%N�o��ML����m�)K�CU.�E�*]��/3�ڊ|>�Վ���v���8j�,�N5��nu^H��aX��G�B�	-��~������=�����w����nQ׼Ŧ�97�漚����(l 1����$8�����O2蓦&���LY���AKj��}4�!𲹳���N�g��6]m
���}�\>���o�2B泘�U�$U`�=~�u����{bg;�P-��=����,�OD��݊��tl&�O,r�t5�G�ǔf�s��e.x0��{���w�4�`���7)Nj彗���2S�B찗3��TD�5�^²u����S��ms*2[�@y�cdB݌���Q����dS̠��S�TS6K�_M0-Ҳ@�oe[7�.�Ld5�+�*LF;�#��x�������Ӌ:kvoB�ߵ�%j�<[\�d���	Z#.��e� �y����J��K�������6��w�� �A�{�?8��+��У���z�h��n/�i������~�8Z#�6�m83���bu�nXJȘw�C�H҅�Q�>x�I|��)�b���1r$G腵%1B��w<�8�s�dnk�l�Ff<�w����T�,z� �\�c�Gw��忖*DzF�>�F�_!�`��^��T��M{�o�:;����SNpƛN�p����3~%3�4���h�J��P�z�\O�l�hMUm#��q�j��=�:�C��k{{b���HG1])�k��"���\?���3����:�F����y��2��;?���0�1���� 4}7��a�L�O�l�T����׆4�.�N*�o����`0]�l���߃u;i_�9Q���O]���A��v���L�"�R���DW�0q�T�ۤ�(u)]��$�e��C���aJɖ�ў⾆�fO	C�e�p��;�E����焪��W� ���{�e�ڳ����p_�_ǽ�nC2�R N�d.&���X��ޏ��B�r������v�'wc��ޖ���N�(q��?y壎Ԕ���f�2�ln����)�o�Q������`D�Qn���a D�mj���jm�,�⼭��p���O-�\rߥ�����qYG,�G��m���۔Ê�c��^%��+*��ȫU��[�h��I���h/L2:��	���?�
K�(��>z�EZ�[i�1ERhڂ�<�{�ގ��#�]�c�
���k��lqj�\��Q*03;l�/`�֞��*��f�?'�=��Q�`xc�)�d���]�=cD�l��B+��w�"K]��E��˛K0�p�F� ��ĸL��W1��ۃ䙁�DT�c���g�M=%��D�9�^'����݌�؋��X��r�_�zj�\IXG�8rm'����صYٮ{��xPM�4����[<y�	����^@��ϳM�9�<ߜ#̌a�:��*���0��u�W�K��l�M{����r*��ѕF+��=� 
�a��R)��x�4|ȅ�r����:��q�P�KM9�����8��� ���/k����[	�җ��"��f<�	ǵ�����u��3�>�Q�&���Y�'�1����B~�����"����Y
D)��7m��$�������.�߀2�%Le�����ώ�bs̮B��}���K��~ا�9��������_>�@�Mִ���x���%)�<v����o����%���֒�{�����gA��|L�K�A��m�Rz=>�)�S����l��-��^g��C� ��D�w>�� �x�q���{�J�0���@�f���t�ꑢ��6o��0�X�	{h��u�zF���ͯ$��p���q؂��xʄ�yE�L��c��4؎�9��l͛������F�����]c�
�|kS;`��x$|�$F���ʱ==?�(-{Zi\|PkiUmRب�ҨH���3e�pjG��yFݫ��[Hf��z?�H�ֹ�]��z9W<�rF�ן�軌���~Hw?Y��#x Pyl\a�(���ps6,���UV�8�����o���x�σ�j,�O���Iϝ�C��X2�z2�u���w�,:���nH>X��|07��3��+A&=wŽ�B9���q���H�G�oȚ���!�A��P�D{�?����*~>�7����s���./�W-�*i�s���s>O��2���6u�*_#�9h���Ӭ��,Լm���w�,�f�t�7��1����z���:|!UW5A����,���{/:�Zn�`�uة=k�p��[�M����z�����{�/�8#A#���Z�y���HF����[�z�Ҧ�|�n4԰��T���X���El�g��4sz�����N�I���'�RԴr q�kɖĜ>.]M��Ŏ	����&iJ�\Nef��Щ���9�C��� ��erU2nT�Xo]�4(�Vz]Qe�!���NY��#�k�C�!!��G�݋�gwf8e��џ�Q5���R��a��8�-��8c��yy�+�Q�Na���Cw���#+q�#�?VB!"��N><g�T�_99����9������b�mW�Oh������:˱��}:z`'zv	�t��^}��i\��ׇ��Њ����g�V$���hS�$�fZ��N����[&�a����;�r6��[ݕT8:TǷ�/\��)��N��\Pv.��:�W�W��4|��]�@���6�^�����\;ٜp�D���͟��N�8䙌���uNw� A3�l��Q3��B�	4C�QO��o/��Nqe�h�&������K$�3�t���5� ��;o���x�|C ff0^y��H�jR%����Sw=j��",�e�����b�9�$��32��P*�!�)x�����	�l�gd��!	c��i��	%8'��σ�{����4&���W�@.�Ys�sA�B�<	_,���˫��P�rXgQVc+����pQ�P5z��}Pda0�$\����[�i��%��W4}�	�=�ۺ�ƃQ纍���Յ��wu�R���-C!�}Q��W2�����EG&9�lg1��u�o�_'�����Yi'*0f�s��G�����r]��pH����b1�{շ-Խ�3�=;7�:0�H4q��O;Uc�pzc���#Q��V������yC�MI}.��|���@�4"L���뷮?�d�+VA���R����"�|�" �_r9���|�y�����f�~W��d���G�����|�x�O�b�YPy�R�Κ���xK 63�~=��B�$���|�a���WH���D� �1sx~�eￓ��Ħ)]h�Y��9��	>v*�M�ph덡3�&��Kr=q��|�}]e�4��U8�\Y���_��]�3$5oy��x�X9��l�St��y$G�eTQ�����E:�	
��-���:�����
��`�	=�%� AÌ�/�٦� ��A�}t��FGrP��P��;�n��S�8;y��}"�Qet�?�M�=c�?��W�C:��������KU��&�g@�{��o>_�8�VZ�&�H���]����M�oѪ��?��$C��Mv[B��+9���c�ʹ�1A��l
s�)c9Q�o�ʺu^��G�
��[C*&1��l׀�����L�l/��A��4�m�hI�N�!Z��6w�TQT�������ۘ>S�j���*;M�ҽ �L_~��X����22��w�:�V`��Yy$߳=p}�R�d�+G���U�oJY�[��p�R�^7uxw��	�E�11�a,��a��E�Rɑq����o2��k�y�IX���Ŕ
/+evY��c�nQ��"���O�t�@�����C�m�Ajr�[?eR���"��;i���F_'��9�%�E��GiL	���}2ZpEa/.c�$!k�^츫X�qN��0��7�6�Y�aH97��0���Z�����������1^&�q"Zz����DQ�ǀ����Nca��[5wJ���4�k�����*Pr���+�BE��R}�Gq�Օ��Q���K�F��߼������t��HtI�����=ҧ	��g	B&���^S2��0��OT{ƙ�f3�8��NW06Z���g�{I�\u�陫n~�wJ�m���[���H�+��j��nѓ�|�����e�Ȳ6�Y� ���X�b!.�y{���UU�À��Y�6��)�b��N�	1�+\T|�kɀ;�+@##WH����b��.p����]�MK_�3Z�g�Lى҇F�Ȼ�|�fEƾ7<I�~L��2&G>�L@�2�C��#]��/��M�	bv� ]���j��JR�hu��5`�1v>W��j'Vy��x֑��)�9o��}����f��|k�s�WH�
CR/��~W�692�Bf&�v�n�c<�K��,K?�ւ�^7"��j��UqI�i+�A%����^�>&[�XOG�ڡi���)�^O+P#����o��i �L"��*�.���5���7�U2�	z�P��En�Ӿ�ă\ौ�Z��:(X�`�������6[e��,��T"����P	��;4�-E|	í��������4|�6�$��wt�M~?�[9]S���R�ϛI{�[d���,�n���t*.�~D�Ї�.@�E�тp�����o��G�q�w��N::c3���m��ATh�:�x��+P�;�Σ#��mY�ƽ�����)`�6�^\���A]�=w�.�L�u���I)t���5פ���i�;���_;�Es�1��A,?`\]��������ѯ#R׆� c��".z�����J��{L#PA��}C�f�_���#)��eaK[q��������Qj|:w�����Z��Dާ
�9�hR�0�\�y��#R����������i�dh~��o�?����K�6�qz����Ӕ�@�����q7���l�N�h�O�i=���P�a��)|πN�.[�\dqğ�8ϣ�u��ߣ��fK��Q;ޚ�[���h8L�;���һ��"7n��������Z��3X�+�����2gz����	[� 4I�"t�*0���-���FA�@Z2��1�ubwv�lO����T��ފ�ႄ�&�@E'��A���ل+�Ґ�.���Sx�N!(R?� ���v/������h�,�~�AX�>�C���E�$!N���4��4E��Ҧ����A��&���<�L"��n� ^�,��p3y�\
A�A�Q�j8{,3@u�7�X�T���R�ߒz2��s1��V_Ӑ2�õ�k��g柵���<`�Fb�u%��F��@��W0��g��p�#��[L=�\=V��vi5�{�L��h�BIO�*ff+�xdo�^L=�$
ԉ��gd��{�M��ǂ2��1���IN%y�a�;��f�r��ޤ�����e�ԫcI:+���S+��G8(��#=�v���+zՁ��,�s΀kb�L|}-�*h���K� q��&0��y����1�H���b�����	G�oE�mX�^�
�5����� �|m�2�7\��#�n�]�3���Ο�K�9��ԉ:3�g+8���g��H��}�$j�S�����Qp�� >�9D���$�r,߬ �����D�<mF��;�SJqރ	zX�U:��m�p�˳��Rݸ�k��,�\�d���P`y�qb���bc0OՃE����(}�P��C%����0��(!Y�t�x��s�Fyˁ�y����i�؀o'Q.���@5��lӸa�YX(� T�V(E©�T���^-Mt�	��x~�}�6N��qT��w�bJd�sSK�]T1
h
1D+_�*Y��e���]�,���fz1�k���K-���'���!/akSk� ��L�������C-8�����=4`T;�;B>5�t'�l�)��Vx.VwrE���l`���]K��q���G��sB��ʡL�ժM_p#JNz2��'��Κ�K�i��l8J/y�\ڶ%Z��h^����7�U����dO��b� ۀX�S%��a�n���2_�|iX����!r��%��r�U�&�� �t�f��ڒ�(�+VI}EpD���^@��]���Nt���9^�,M��'?�V�fH�$j>���se�ċ�p}~�Ob#O_��Bzǀ��C���l�y�2��t��	4KpDi8��Q}������@�Òƭ��"bފ��tT>ֈR�Hj(�eU���9��V��X��)�u������H������K��ۧ�=�@�L�+�d�����_�E[JyU&�^�<�	���yȽj*�)X� ş}��5aO�����7=.�;%����=��Z�q���Sy�=?���H(d��!4�
jv��iH���b�'�Ś�%U���B�!����C_x�L�A����n���m}�����<�J����E6�����+���d�N?�*X�D��F�r*��������@Yt���C���������.7�
N{�F�J�?@/��!�m�;H���֌gF\��@Q�]��N>E���YV��<��Rw�*�*N�^�OKTT��B���ƨ�;����m��RA���E"0�P>�uY�L3����|�l�b���i�$�5�_��T�YT
��$w�\�#j�ͱK'@r>}���-S ]b��'�hʮx�:|]�c@��xC�Sqè��)nw�6
�%��\�u�ewc2YK΂祾Dիm���o=fԆ����� ��F�6e�~�S [����a�a�?sɌ
� ����vb*��������6Q5�Jp��*�|)Nv�Q��P&���QB
��S��<��T
��ko��|�޳3l�@z���x�*���#���ϯI8�Y�|�����x����B�C钖jM������U[�5�Ϩ.�Uj}u�En��#̨q{E���8��7��BZC5=��6Z���6�9I�Z'J}���e��(Cg�9�QG:ӽ	������� 6��2D&S�ߑK���X#��#�=�v+�=��L�n���+��<�h�>�r�e]]/�k�dc��z�j�(L�y*"���@��u��
i5�ɕ�E�ٗ��س��4��� ��������%"3��y�V�����з,@'���ސGO��k�ׇ:#��To5���Ѽ�>\¤���8�[`%���:�*���ˎG�'Ƒ��gkHf�(Q�$��+���}�
n��>rz$�ӣ[c�'��y���l�� %)B7.\uI�~���ܩm��b����o"�d`9����_.P��a���{�M��'�r��G�r��R�����n�ǲ��s
�C�-�`�6�p�������,������:�<����o��d9z����fC��w����{�WI��4(��<n�GC�*<��Z��i@��)�=>� �Be�GI���4��]����8���l��CK��V�,��n�m����2,��[I�c�A��/]H��,��Z���K*H�Vyt:�y0I|?�L,�5�qIpJ5�u�@O�����
�QL�^ˌ���щݣM2��{_a�D�ڷ��aK��r�g�d�Ji����z�m�wd��`{*@�n��7�P[�X���c����G�u��po�w_/&k"�A�S�Kr���Y�5�<-�s��-l�n�������e锑ᜩG��jC�.�[�=��ȶ���9���V�E��\��Gyx@�0����9C�fJ��=��iz����,�L��|p�Y�B��6R��q,n�4�$�h ��K*���5d|���I\x�[&����r�S:����|難­~L\�q}���X���1�$5�f�L�\�Y�C�z�^�X�(��a��Қ�-3����x0i���f�0깱0��7m�O��mj�k)ls��y��Fq}��˳�gw�CLG�lΚ�U�?5K`Z�e�}�[J@���\R��'�9$��#�� 4ͯ�F�M�K���eL�����[E_�	��	��>hH�t�,\��.����4�+tW��W���@���/�3\�kC�>)$0�z�a�0O5���y�����f��Y*F���iW�I_ �3�z��5�:���V�~����(h����5�aiFA@r�}���А5'R���K�c�YA7�_lL�)�񺀋4���Ea'#�)"��X2�Ć;@� GiS�q�T�=��/tp}������i�WZ�um�0���Iaª�Z���P8t( �W�)�@Яxj��o�`���#���V=�Gn��`�!���ʴmR��#s��XIy�
�1��FEU��[J�-�1��}�15m!)H̢�S<A�H��e{�M�p�Y�� x@*g\g�'�0�Y0Ec/��Y�����o�9���ei��qA�|�>x��A��LM��,���$�����n��g������j�[w�����JT�/��ߏ>��FӃh�b���QL�U�Rh'�l���ɸ��G-sz�g�(���۩U8�������7+��\�S=༰.���=����An,�ڗ��[ޫ�� ^Ut$�>b'at��8�P�A1V���C��� 9r�eH<0ФV�ʪ�O����z�H%
t�KU)���7�+��mĳGgh+�e_؂*$���=�����>�B�C963g"'�!YJ<��W�o���_�t =SA�di΁���Ɨ������ᓺ6r�!��*ɑg�[�۠p&,��'�/����=�L�j�0=��sK���ϙԴ�[��&J��6<'�2F{��D��|5/�SpO��Ǿ�xy�ՑpR��0��>�5r`}�e�v�2�Z��)?^�l�B���yc�
�-�z�c1��6�H����5E����s�q��$�����oZ���N	��uo�4��U��b�ս���3�?:1b`��sB�=�)�`m�w'ڶ��edr�m�s�~p��ބ�݄a��{��<IvȍMT�wP�b]����k���e�n/�Wͤ*N�|�������� ���Ț�-�|�b�i�Q�M��*���Bhx�@-��Z��F������׏g�'�"5<���Ņ�:���E�E/|rS�U��3V���h���RZ3Ϧ�����=+m�=���_^9$�b�{5�t�˚KN����j����t����͉%�C)�@����3��Y|r�-���s#�E�;��K�'�q�ѐ��r
���q~��e;� 2:ۯ3ɍ7���m��A0Վ�x���F]BfL�H�2�Uo��{Y���o߮C����:�>Q��<C�q"`�l7s�v�����J&m�{�+�W{����{ð3ɳ:,��=��Ӽ����d�;�Yxb��uZ�6�|�ұ����@��^�Ωj����i>��<��VF�jW֐��x�Y�l_%��q�q�X_1bE�ӿc���m?	&������#[��)Cǚ?0iQ��O ��1s.t|����*K/�L8s�;4_h͒���B2[@ �����q�36kI����հ^�b�8��o�%^P��1
>t�n_���޶Oq�d���7����SG^�ŷ�&\�:Z@�A�8�1cGH��(e�F��j�;ׂ�+��N�K��9	��ݢ%V�ʨ𺬴�I��.�i����~ˡB��vj�K'KO���Pz��}��;V��r����=b�[{:���4A���b���\������E�&|Ms�`��v�7VR���	�[V������S���Z�t��qﰆ��1���W��B�/��o�(�ꛭ��Zp�؂���B�����t��/l	�B�gڵ�CJ�/�_�����ާ����Uk�Ǿ7#�5�L�v�$s�z�"F���R�c]��mj4BR�#>\��4�ߣ줘��M-�u6�� �͝q/����"��G�ڞ!��>Z�o5q�zs��
����+��@3a�r�*I������z�Ԏ��=X�Zjw���֦}�c7��k\w-'�����C�E���Ї�g�}�l���Չ�tn��:C��T�5�E�ZZд�:�7� �K"�}�#�g��,v�1�j!1��N5������BᩤK	���i�&��NMt���~y��>��tra�2�-�իв�g����CZ�b��m������7[7 �!U�)5�zŗ̂1�%�m�5�q��m���6'�1��n��҈���;��|�U��&N�������
j.�S�*QH$A��5�o��i����ƀN��S�:���k%���.�wO����%��D�ؕ}+�7f�.���njf/�?�l��-�� wC!%N�v�9L���h�R)O-q�r��&`�gI�f�����_��
��dN8�5�$~8��|��v��F��n[���jw�Zt�%C��O��g��H+�:� �h0R�	�#�M����_���C%K%��[�����o�[ap��@9��C�J��nf����!hXO��މ"j,��0R�WM'ǎ��ӷ	'���:޹@��ѿ���=EJ�G����n��pHy*��HVD)���͇쀂x(�O�h�*���Ę�Q� �	|zo���a��(���H'P�o�D�c�~���e�����3��O2����Y���~�E"dgP��&y]ոr���-���?�Z�s�=MZ�O �0����ݎZ3�C���)��%�Z�N��<��§�58�<95Z�:�A���EP�}��X���㍧S�))X�u�§��	�0ch�<MN�Tjx��w;�����w3��g�ȁ<2�����.�$�TƮ�p������7��M;[�]V�L�wE�8�c�G�6��d���5�����f�h�Y�1/��Ò����*���Ɵg�a��㪧�h����k=7֩�0�� �_��K�x9I3Cd]��U���)���p�b�m#�G#�� �����=�/��qț2���Мݚ�����.p�Ӎ/Ȟ���"���u��`N�˅�\�w��)���x1ҁ@Z� �a��j-�ȶ<������^c��B�,+�p➴�r����@�����K �g gt0��%~�� �cY����^+00����%j���G��H��^�o�z⇎k�X�,�*�g�`�^�x�;Y+��mhL��h�C-�_�FX�]ӄw��WO���b�V菎v�w fV�Ue�����q=�k�-�Բs��z�<?Pu"���@� Ԡ����K����_[���T�9O1�C�$��mW��E��p��[i���oʝ��r�
P�p�_�Ѧ��0��y3���@,�2B<�Ű��8ۜ���I[F{�<��A�Բ�\}ݐ]=���<�v�ĠQZԲ��~c�y��!ܾԞkr�����|q#��=|�X�c��NZ�RD�)f�*��&�����A����ej_��"���Ҷi��j;��C&3dzLG��ԱS\AUŗ��kS��K'ֈ��|v�����P��SY�ʈ��ITG��3�L/D���͙(��[s�8?��$�c�v��ނqblY����I������q�z�w��Νc�A'	�.C�����J����0|f?r~+�/�#rո�������	\^z� P(�թm;�J���Ά�N���
������� �]�NO�[����>�,yM�~�qm+N�XE��\�_,9}�w�ʐyu쪹裂���q��~���W��#DV�r�iW�0
	w�&p+Ǘ���J�& ��Z��|���^�F�o{�Q�on\>�υt����m촥A�Y�3/\D#n�!&��M�V	%�Q��#;Ħ-�Q���5�5n!����q~{N%����l3�*kI���+S ���Z��Q�!���'�[��l���Y�#�1�M�+��P|�(é7�	�'�/4�r&&��,)�Y�W���D���ݷ.�-�83���.�����n�E�>�kU9Z آ �3�!�D_��ò��W�OL�q��i�qD�X��M����]J�܈��)yP��P��� �x�h7d�p	���%i���](�(ό���q�beP?�h7v�q��	c�o�>���Vk� ]7����$p9�G�)�5��.��j�3�ƪ�}����m�I�t��p��)n'��e�&��6�tX<10��]��4a1��hb�Ob<zG��+��	Ǡ���
:��i�$�/z�ntTݡ��i	���J��QE;V���8ar�"3Y��7��K_y	�ی��F>K�1�}��|给�A2D����M^ӯ�TUz\Լ����k�l�V&��,3��n��x�"`�n�'u���;�ч~��/*����sf+�,��S%��8����X�h���+|�|�,-$�(`N�/��/y�wi���]# ��&�,�vX�a�<�q�ma��ށx�Z���t�VpY�)A�MaO��������}��٤A@�Ȍ�ѽb��e0+!�����T6��@�e��:�&��̘ {�z��b��c)8z�
����=����G%Lk����%���#|kj����Lf�J�ϨM����"�,�� ����ܶ��:�YZE>��Q�[�hr��' j�O~����׻����.�D�<K����V�/t�/�P�9�A�7'�t��D����V80��?��1�0�"����\&�喠eF(q�E�$�}!�2�֯�� S��?t4��"��7ƹ4D�U�*��+��ւ��!��|v���[&ぁ;95v�"� �	�]�a���D]�hv�Z^6ufp�9���^m��?�T-�^�Z���J�+�����魍�X����ת� ��әE�$�A�*�sz���S�#��3u4�놲ӊ��X$�8�ڥ-J�A�&�S1�o��v.K�S{�:D��Q8�Ұ;��][����o� �u��F7�K���
�D��5s`.a�
���p�I��J�=����LchĹb�dnF؀�2��˹8Eb�8���DQ(鲶����X?��C��(6O��}&�D0��[���0�;��Z�_脳<��}b�)9�دa���tE�n���{O��A"��3l�lh����:%c2C�f��U����B{!�| Y@}�p���~�~uM�[�E'�{#�%?�R��ej���b���X)?[w�v��{�-��vOm��#�m9�xު�+:�+��k����i0���[;Fx6O����,���LP��%�*�e`7
�@^�:�
��V�n�a�_�2�,y���ۄ�70,>���� �L8�Bi��[.���`/<om}���*;�� �xV\��.~�38�v��oDd9����v�c{����n
&�w4Q �
��~���ϩ,	�-�A����h0�`��.��R5E��J�T(j�>bCȭN8�{v����9�!�#��
�҇۱`դ#c{j�6((iH�H��q%q�Ix��{Ό�雓eu}&����[ʫ�26����7�?�dˈ�n[���>CK�4j�O_���NcO\����`����&$h�k��N��o�{!ܚ�#1�J
3���a���B�ހx:wԶ�V�� 4^�'�=]��E�ࣼٔ8�y���z��L~�
bz�po�āz�͙��X;j�[t*O�@��h���d���ϟ����B�8�>T��B�1s�`�]����PFG50��4�=*��|�j�p$����[#��-�4���TG7D#�:����,JQ�d7N8H=��~�=�$�7�q�����Q�j�#~݀֜ �g#���Ȗ$�H�
�s\x���b�k�8��PT]:���?o�,��u�>��Ԛ��C���:�D��`E��P��2�0��k^
�̵�L�Š�ͺ�}>�Z�YbjqKv%����?�f_7��t}�a�,�@��n��`�G1a$TF�)M�i<� ͣ�M+D�4^!�M���IDee86 ,��3�ZS��y-m47�hm�;h��I��S�.��- O۲>7��k �輱�.C��~��q}w��`�hL+��.�y��W��	�����i���l�5r�>�wa��Jq۵jf��twz=�ŲSqȤnxy�>�`��0Ę#�x�slV`wQ�΂��8~~��"��
)��v�7I���+p_�v.�pUO�`�����=��NMl��~2~IN ���wx���b�u���:{��|^%O�\>Y+j��O�ǁ���?�5Q���khW���b�wÚGya��]!q����G!C;�@`O�-�b��ဂ�}Ϲ�}��M{1;3:"z>ݚkH�(���}�9�$��������F����t��*[�!������cS�����u�&�s�|]k�U���;��`;���
�״��Y\v�w�>����k|o������|;J��J�9Vu%v��S�+R��2�&�^Ñ��lW��OĐ=�+�������?�l�(-Tڋ|�XL�jmj-�v#W��cY�H+���]����q|v�J��a�=���gH���<���Rx����;U���{n+�Z�`Z�GQ�/qپX�	���7g�%�iΕ��<L�����V��l��e�����o%߳��\p�6z����� �{�?�5�B1����"�7�$s���hw-#��u����^��_i/�64kl��w��/K#�;Ј�bۥ9����-���a��Eٸ�\}t�4~D����;��H@�����K��.�z'�R5ie_�G	'i�������U2�N��} If�?@o�6�a
sN�U�)l����ʇK���Ĳ��"����IZ�����z��}Q#�i�aˡ���P֮�
�mI�6��	��:ƾ��NV����y��k���&����f�����.Q�#�yQ�nm�Պ_�K �h��?Rg/�#10��L�z�2��.P*�KJ�	E�v�>��LKOru�U(C�^5�Ө�D�6=@�5u��^I���o0�F�6ʬݜ��Γ�� ��L⛺T�X��_ۘ�u�i���S	�5C�v�8�d�U�N�0EQ�g��.y���V4e�dA���Vl!Wפ����T�ɚ� �j����J���u���'�j���-��X_�t�uP�4��0.��FbHߐo-��j�TdK��5G�.�I]��.�M�@w
G�) 1��(�ş�n�u��'ش��0g{����eD�P)��N;nL�H��=��4���sM"B�m�mn�_�����w�)mKKJ��~��|V��x�v���m��%{��K߲t��wkSۢ�?�6�o4oP�J�P~�~K�v5��1(g�� ��,�%Us&ݏ�<��l8��sF���n���G��z] ��ʲ����J]�g�M?(�F�ho�|��4N����Wy�������ܽP�_���?�Dw�1+���TM8�>�!�&<6���%ٕ�L:�F0�����LP�]K+J������A�+%�ŸՈ�Р�G�����i�`���!M0��p#�k��3W��^�FqF��V=Km#7��:�n�ΰ0�@%sU�n�G^.�~�b-3Hh�B|a�c���R��~z�*:����7���2��k���X�`����:��@K�iÅ���ރ�4j����܊�Sr!�wL"�mK����M�Ű��Q�����ð ډ�&9A�5u��/Y�$JKN!���)�?��%�w��_����!ߧjsC�q?���-��6���T=�O� ��������-_A���P��O���d��g�� �ά�F�^:eS��@HP8R/���Ze*:Z�K���J�w�ǭ2ִ����A�b;2����=R��
I��߉⻤@���՛;���U�m/�����	H��~-ƾ" Y�Ȓ��D2c�p1wN��rX�D�r8���B)�Jwζ���iֳ ��/� ��"��1�a��Q��y�^�@���&�;U�W�z���F�4fv1��GWA���1jȵ�b���tH�u��bq[�`���+�<�Ȕ� ��\lB��f=>���L%1�^�㫦Ȗ����$ʻ�Uz���z|H���V��0�ȼτ�mp�"2j��K�"�)��Ri�JH�2G�e����w�����.�أ�P��-�*=�����)㯹�*��<p|:�T|~呭���#E�$�s�1�=���Ɲ�J����|!�l_�ܖ�Z��� a�8����C��YI)?Ɩ����Gx�y��Sϑz	X���r�@�,��W8y�2��p�!����j�� �����m����I@md�i�q��G�e���'�Y�P��3��������כ�F'�����6�塉�ݝ�6��O�u�_	�f�0�ǆ`���[j�B{�C�<���w�U��.�!oVT�'C�\;bl�=�A��"u����x`G�~DK��C'��%O5T�Ƚ�k%*<�j��=_��!jq��RW�/	YMf4wn�FF3�����0���K�T��:����t�+�1!;�Ѯo�]���po�|F��x���G@��I�����.�~�١�yt6ɿ?�^����?Ib�uf�uԹ��SK��F8�[b��a����D�$7���_l���1�j[�0��i�^w��SU�8e�c�%�}��׬;H��/@�툆{W�9���#�8��M38�ȏ��fe� ���d�^;N ��驠�hk�eյ?������e�Z����[�r�;[/�1�)��U�-:Ҍ*��j;$�A����� ;�NД�/l���W3�dn�H�v�Y�C�x�'N��`q�<��s=���ɥ9�6�AZ�
ǚV����^[�V+p�Q�`u_���-���g5��GZ��t��&Č�<ݏ��4��9Ėf���ل�;�ݫ��~��
�Y5*@9�(5�"KL��ꏫ�3s�c��^\\�#��0q0�Н�R��s{q�|
@ǁ_�
OD�6�FK����@-4�4+z�k$���$�{f�F�t�������0����X)�S���,� ;O��a����TI>`5������8����� CK�[�G�&��F��WZ��]��T]�� �Nd�Ց�Έ�O�}"��T'ؤ8x���߀pt�Ϳ�* �3Ӆ�8��s�!�J��:g���j���FB�SP����F[i?+��S>�_�  �������Je>��/��G���a��G�qq�[d�����<�L�3�M��l�z���E��}OC���s���{�˗$�b٫�K�E����Ȫj��#gV���ᗅ��-GW7��;= �l����'��H��cI4\+�Y
�1
l!5d�,�e�#�׏����:P�
5 *(9=�A,�c%��.aZ �b�-�(�ߞ��:B=��S�{�W�]�\B��b�O��H�SЈ�k�a5��51�'�;2���l��Z�2���ў�]���`�(�ٺ��f��L'�	��c�e��	��B�޴%k7mu	�0��[Y03�M���:��jL��S+�)��R����e��̬?��D
����C����HR�IO��'���ɻ0��`nZ��M���~U�n�ա�i����T�d��|W�A|{�~��1����7[~�i��V�5���:@0�oѥ���&�͜ο�l:�`�ņ��O v��qffZ�S�}�Ώx����o��;yY�G.u����1��x��IAR�R��3�͟�m���9ϙ{�DS��TOH�o@<`�/�uG�>9ڥBN3�qY�;�W*8������&��_8�j;B� ��L��|��H�$A�j����Q�u+��D����p�U"b�,r�Q)��\��d�PZ}S,q�^>:�A��h�Lٙ�H�N�B`�o��J�1�|��i^8�o?���z���(�'3"�ݍ���O:,bÁ�mW��҆�Y��#}�}�������!���#ָX�_ƅxV�N��v|�]����D=��V3s��u$ 6�`��}Ձ)���<�����*-���%�:�C�Jz��޽cbh�ޝ_�z�KeJ�K��%<NMԯ���6	�uE�+%}�ƣ>3/G��CiL�N���#K��Z����5Az��KX�CE��.;M{IU���*>P}�14>���x���T��UV���+[�~�S�f����7�Հ만j/�Z-��y��M��!��;�L�D�L2;B���`*o*&ځ�=�P��񌵴y�]��R��]-���u�[�"��ONCY��i��u$���9���iػ�^��"K�/F���G*��	҈qH91�uI�}/�+Vh>7
�̕���P
nꯋB6p�=汑G�r셩�?_&�&@|7��I���� ���|<��t�����[��Ki"�)ӱ����^/rCƬu2&_�>��h����,������`]d�����u�|��2�w�ր� ���} _�t����ʈ�(@�Fy|êEx�%>���W�������8@-=���eb�W�䮲ls��k����CӉ,�ѣ��:ٷt�4����2L���DU���
Dޘ:�K�_���끄�@��7�
���g��49z�0�m���I��g��Du�]�Tx����t���EX���?�ތ���[�F���f�@���5�h�+A@H�|��Ⱦ�,&��G;�]3���:�U�풜���9(9 GK�ľ�@�M@�>�bd�+c��U���D�V\���gh��`���d58�L9|-b���n���Z��� ��3?Ɍ5�MI�+��9��,ɽkN�����e�9~/���ȶ�)e�w\~n/6�s{!�u$.l�W�@	I�%��Z��q�k�H�XD&�E
�_�0�.�(�:�V�rM�Q�,�Y�Ga+n��z��sZ� 7\��u�g��dT�)G|�)T���y��)yv]�'���yTt{���QWb�.K� 
I'�� y4xXh��$=6�5Bhx
�*��a{a��Pif�IS,��ZH�q�/���[X��:\�����T;� ����|����u�g<^/�fZ�{�Z
wa�`
�~ۋM8{p朦�v���t�@;ѓ�ۍ�����BB�tqd�\Q-h������%`��v��ϋ�r&S�I˚FZ��	2��2}v9���m����+-� :�~�B=h��4�:O����;b�?5��i��e?��UTZ٭���ͮ~��N7��q�~Ĺ?N���r4�S��Ce�j`T���Y�h�
7�p"}��O��y����2��*�N��Co������穋��A[�$��,�#�s�����\�$=]:���ǎ�(�^��´�p�<@�b{��<l*p��,�]mqON�hH������[�1=��"�F�W �v��nm$��}!����h(���I�0���A��W�H���,��V&B۷��	3��{7#���&���;��nߒ/� �"+�çӶcm���;�گ(����B�U�ci�a���~I?|"2H,��������0(�'�y�qF���p��� �H����EE���p�S�4G�\W)�2)II�j5��d'�r3Hs����5_�@u�����
� ���.8ߐ�����f�����/�W��d�w���Q�O�ܖRS!��E�ʾ�ٿ�}f5I^@ܵq�8֊� ��Q<=)��M��~���tF�~��8�㪋����F��y�'=�iEL��'>��q��?��a�d�ٚ�ƱpM��j�nː0��Gs�����X���O}P%� i�3~{PF���̿\����#��Nq�H���ȕfQmj�x-*j�q_ڤ��~����W"_���ߐ��6�Gr���_w#%#H��	ό�}@7��rYo�ߩ-Y���,2����+�ϸ�z���i��h��=����G�@OkW��C7A��nb�����U��Y�BV4�a�=Vފ�8�G�U'����]���Ӯ�h1㇘��[FѲl�W�?@�_�n�z�M`���N�W��0Gp�����N$����/+�%��l��taE��������
�&g�Ku��%�=q̤�31��i7�'�4�ؓ]��%������Lj�p>�����xC�1I��l�Vt%���k2���I�|�_��e�)��.�_c���1u9�W/�2S��zJ)�e�{6���0�����{ȕ!����!��)���GV��gI�J��gl0v�1���b��~R��dw$CF����BC~�#촑��$�1��"���F�=c�40�b4�s��]Hu_�,XT���'N» �|��?��Op���ܛ����v%W_��W���܅FGZJ�u3�FB�"�iv�4��6�
�� ����R�����hns$�VG���$�4�%r�M�@��|�ҟ��ɚxH���0�|X�8�W3��^�0�Y%���c�7\r�m.��٥��J��,���a)I|�����j�Mۃy���|�T�`L8�U�u9�5�~�����.|x�)�c��+���c5�ȉũ��k(�D�G���OH���4���"a-�od�SvU�ۦ�o�7ͤ��:Py�%�Ps�i�Mb�|b!+��{��	�u����9���y6�cJ��C��s,�R{��?)|Ed�4�^mn���ُ�e��Ih,`�a�Z.�q�G�:��W7�i�vxPg\?*X922J����0���P��0�ٜ��_a�P8J�ˢ&:Ea%�D�;����`�Eo�2������S������� �8l-�	L���'��203�U��,-��l�-l�*�.x!��g6뤰n��`�*+uA\9��-j|'6���*+�	�UG��
bdw�t�_���j���y���m��p'8�z�Ç���8Ve6!؈��,_� Y.�c���̩��\0���>m����4X��������'�R&ᏭTX�/mT{�>��|]�F�:�(�a?���h,��r��2� \��z���V�[k������R���� -����{}���P�:������|-m��F�|pcÔ*��Y�V��2e����U�ܐ$Yw��+,�#~��x{n��zp��+"��"50e�֢J�L�;�dqׇ���}�^%L/�3�c�rˬ$�>)x������P᭩��	[R�� �8!�e�D����xWi����5DN�:�>0�F�f��h��i��M�p�B����d�J���۬:n�UR#Ǔ��V�@ _�9[�d�$��<�738��b�KQ5�%�s<"�4�(ih@��Lm[ �Z��F�*_*9(�Ύ��R�*���J����$ٙ��L�U��E�ѣ��z��cODs�ʦC�V��S�4�Q�T��<YC>�3���JV;�Z �Sc�>�~B�b3,\��B��gBqy�)5l�=�z=}M�P m;�6��"�8Z���k�wS֖`&I��0�����If|�黶V�˞��+C ��T{�f��������~c���/<�5��ԏ)������`��8���N,M ��
#B|�D����X[=�#Ԁ>��{!��
4�ƄX834���+��	���5r�����iM�:�0�<�u8~�C��:EO����xpLn�.�:D��jb�f���&ӟ�����k̨�0��R��B<:X��׍�L0����uF��ʌ.�M�e�^TvUK���ԍ*x!*�G��cS��ڐ�R����eL�v^b�{É$�+�����|�Qi"N�n���
<sٙS<b�:���� ��':�3pH�0�79ܭ���Ǒ:n�� ��u\i�B���������B�ff<Px��wv��Q�D�q7l��	�X��Y|m|�"��'}Ijt^a��̫��z�_��'�o"��j5e�'N�(H�����?d)bNF�X�$҄x�nDjChv�����tqC�7�����-p��G�_N�9	99t��r���v<�ja	y!o�ŝ��Wm�.�\a�T.�^�Ga��ΓS�$�cCj[�,$3}�K18�3��E��ō,%���B*X�}�X`6���8��>=H��?eK��U�%�}��x'�&4B�!������dx�·Ӹe X��o�J�dA���js�2g *M�l~}p����C>򛢂2 y�}a�ɲ3~U�_���i)��ub�$8���ꖭY����
���h3�^�SݖrA�s1�
���|24ϣ�&��=�v�|FM#1l�����x=��!�@��CɄS�0���s��^����, 1������|���۷�yY���*`�"Z���B*H�����ia�{ju�Δ��:�.��{��i ��þd�A,��F8��s�����O��8��u�<�}�;���ҷ�|�G~�7'�"X���~*���N.��D�f�($X=�B2% p!������y��{�[Zw�;���n	�j��z`�����H�*Ȧ��y�Ĭ�5eɉ=�L7���ZT��Zy�英)>���`���,��!(n�����B�w�{��hA&/�:�bF�K�S8�g�g�<�L����{���v�����+��3��Wf���}�-�r+S������o��T�Һ�Z!���P����?��V�Lvz�۳Df]X^}��Y}Ҝ �S�CϏo�~�Im����V��
��}N�����4��\B� -bM :L���t� [����3�B���\�R��
�����<���&��-ZTb:)Z?���\�e��t�xY)i
�\����*�8R��X�zϛKўY�����5�\VGN�5�ۼ�ݵ�r	�]���HXC��#�cB۫XK���:�u�^��hꮧ��e���ʗ}�e��D��.{���Jq[��:plﻨ]t�Q��0�m�h]}<?� �#�^L��`�i�a�*��%�������H�Cf~�u.*�[�#&q 3���q�-/v�b��������{iZ���*zm3�U"��s�mRqƛF��mBM��vU�~xQ��h��-/��~R�ƒ0���۵����,�;�<��]'�ϒJ%z�t��;e4+�&�vD�$�4ІA(��`Mi�4��Ԛ
���z
zᯪ&]��^��!u�eN3�y_��NQh��S��J��ܭ,D�����Pg�ƌʡ�pjzG��to��V�G,��c��0w��������`��l��	�������{��N�G�p����[><�,�&~|��N41�YacM��3p���{S4���q��̝��#������y�M�����=�J��B/�9�{2�?G���*�A�a��h�ߴ�6��D��\�)��F�Ξ ���;�6$R�>	��7E���_��}a]K��ͅ{`%Z���a㟇M��!��f<�RU�P�v�>4�Sd%?�u`��y���Z^9�Nc�N�p�ؼ��M��(#�w{��K�r�b��L��vڪ\2^Ki�G[��^�j� V�#�Ņ&�����q��4@r�E��22�/���வײYkk�S��o9�|����`�;T���g�e�O����`5������'�e⶘���{E�E��R��[͒;� 	]~6�fWk[Pݢ"Cg2��҃)���ܶ5q`%��ڤo0f�=���;����"6�ŮM�ʸ��+l�n,���
EĚ���U+�a|�����8:�n��[ҽ��ػ�vo$�x�VC(���Ƒ��92M^��]Ѱ����C���Q9�&�n�p��uqj�����
?��N�`��u܍�H�%'$*e'���2�p�4Mۯm��9�����EE��tvb�׊d�����shZ��{�w�,��;׮j���&��`��مtZp��.t�2�[B��:XڷC�y�@R��j����z�J����ԺWht�- �%�*�b� �1+#Х]*���GT@�ՙbCȪ��B��,��|�%�YK�v>Ϊ���)����׆�H64ە�X@.���8G�pYqe!'��/>�W�g����9F�f�m,�������
�$�b�l�x(��l?G��e�L5��M�}�Uh� ��-�9�*�����M�I�d�!��~ gI���C�������paj�j�n���<��J,�	?������
+]Z��Nm#M�u�>����4�W�x7���� �g����H�Bq�A��t"�6�*~!<��Гk�ɸ
!��U�	F��s��7UB���/������k*Uc��>Y�Z=C2^�y�p�UH�xJ���ďwҸ}��\r)��zx�CYp����S��� ���p�<ơ9��ں��=o��?�%s)��6��?�b�+�GU!�����ư	P�������%P�3�)�x�����Ŀ����<� ��W���I!�:��=WC������$��v��u�Wń$� ��zB����g�R�����kɝ`��дb<��%Y�G�{�Xzy�W�tYB%�����S@�w&�+��P�w@�6C@�:����mHWbX�+!p�0�?����G)sҌo��)v��z�`�(���	D#�TK+�*T�=����\�F'����"�@jgG�Q�g�r�������D��l�l�d��̐�V���.ޛ;%	�K�e�1�����w�\��
+I�����I�x{z�"���wŻ���Cj��c�3C�s/$�?	� =�H��ڊ<�<�˓��ƮF"/�����}�G8�w��⛍���i�(��P�����(4��g6����]ʭ��B�C٩ݚ�豱.��A*�/�_�-Fr&h=x��7*f
���Î,���w}��?Ig_�'K��&�#��1�ր����mQ��p¸��y=/cIģ��I���j�}��77�^%�<���*�fۂb�T6�F	/)
>�k8�.�Pih�f���_֘��u����i�0	3���A!Ny�[f�3�إg�mi��UH�L�fʐ7��. �W ��I~��T�_�L	iZ��[����!�<�r�.��^��`��7�������{�������_X�B���y!����
X�@�/� �ժ^�7��[$�8����F�Rٷ ���* ��H,q��~L�lf�[�(
�QF�.J�X��мXK=��㪿T�����V�2~�[w�uZd�V�J��
EY��:&�h������R.�f=��t���G�ű����[u��?Yc�K�<�w��g��8}�S:㞭�|�Ҵ*���%F�h?%5s֝{ %���ާ�,����T��W���� ���{�_��7m��0]�rO�F�� �JK9���'�m���K��@���%y���'�44>^FЙ���-Щ��L?ݙ� �	���+׼0��6�:�>���aS�ܻ��bͣ.8�!R��G}��+�H�N�1(3�p�V,���e���=�Y��`��뉝U|r?�~(�α]VGsc�@}�
ξ�0�!���u��!��<7#��`��T_��Fwr�����C<���\�c6�MP7��D7��3-|(�  ՛d�7�it̉�������=L��6�}���o�/kMKO:��1�wi�i��\#�=�q],��i�Q,M�=��L�ѣJ(C���A�*=���0�y��˭%7�]��᜷�5� �e�x���!޻�������~�7�c�	�e�C�w륮>n��;�2U)�
I)�Z2�ݍ��G1D�%4�|�.sg������Mz��<��<�ᖭW�����=u|�oĻ�i�1�^��6��O t��}�5�6��^���i0�
�i�tP@�!+����:M3�[��F�F\��0�8�3/���0��F~��K�kx`�����.:�tka�/��Xu!�Uԕ5'�\�����{6,c����x��V'���,�4:�)�t_?=���"(���J���Ǌ��]V��\��,�E봣5|EW��;o-�D�F����#�;˹�rh�k�ϻ�x�n4m��'�z����7��RlFE�P]$��q�ό/䘜�$�7Z�bޖ�|�Tp��1��2�O����3�f��dR��.!���M�#ɢLG[��r�ިZ^�/yep@`�J}���1�c��/3��;[�vVإ��s����Zp�x�0S�)�����(c��;�#��cٳ9.`��[V�p@�k]���ģ�u��l��&����+��N���t�A�5g&�����k)��H)��ev.fjΞtz����U|:��1�r�s@*����3�YT�%W�P��@T����r��U�6x/�[*��^��k�(�oZ��0���5����x9�k�&2�>����L��V<DfgӖ��l�BuM�g�עH����s�	%*����3@a�"?��V{G��Vg�����GC�w�+/&ih��	��YS�M�f���ۤV�6�����0�m�D�u]��E؏~��(�	�0:p>}���&��I!����z�~�o��@� �W�gr�'2�j�6IVB/޽~t�%�[���l݄ ,J|�E��N[(�ݮ"����#-��(�.�C�2����� m���Kd��(���g��.F,�3���cDr:*m����Q1��k��#3�.E��R��pIJ�a֌X0z_�O��(�IOu�h�
����!�`�s�|���$��]�#���Hny���F�QVL~�Y�ݐ���Y�`�;[�܊�ٴ~�I'T��Ц3~�m�_̻(=&�]$��ݥ��f	�+���D��^%�0�Z�_z����\DR3n�,�-�7�r7P�W�8����$Q��(�͉�9�VQ#nȚh%�������G>�$���.��~��N�ƫ�<]�n�����n�s�pB���ak	��
9F�U8�=�Ѣ�������W�Q�Rb��˔o����o�n��J�f���lfwS�h��	N�$�<y�����p_�eZD�B�ŅV]��a�������%�϶`ON W��,6/u8M�x��<��m�i�}�*d�A��݄`�i����'�Fz��z"壘/�ÆY9ڲ�om�[/��	o|8�n�U, ���F ۭL�����/�9͝T��=0�VC�;
6�jׄ�r�G|�@g�W4,�(%�� ѓ�lϹ.VҰ��E���z�'��ς3jm��=<��4Vi���g���R�]H�j���~�"k��te����D C���iΈ$�#�nA���Ϭ�%���Ҥҹ!�r�H���)�W�W$�7���m���[V�FQZ�1�!f}��c��Vgz2|��a�yJHl����J�ѱb�bG���̣S�n����U��Oc�W�G����'/����ݽ�j���8(�dh�,��3$_n���HMIDڑ݈�NsӇ�uMy5Ar���x��3D�� �H�4�fPG@����p�L'�}�1���X��#g��:+��Sȇ]|��v���~Y�Kvl'��	/�Y�A�!�=]O1˃�.�&�Z��a��h����<��:<�l�p�ZF͔�5������k�Y� z��$�'�.WK�g�����J:/\�W�]���['%
�^�Z֣�u<� ����"��:���A"O�!@����03?���NC�����Γ%mA�v�s+�����_�(� �p���t?���H�K��y���s?�m�K��RNN�j`	!��P�SN '`�-߹��r�`�_ƫ�������4�,,�c�5�����/;�1K��Sč
F���,����^X4�jy#���%:�D_c'�ea����\��]�;�&@�@M��ʥ�i�[]���.����"Oװ/������=�'��!�˳��6�3�.u���r�Ek�"����i��nl���ښu'��8Ȍ��T!Mz�0��0�~��s�Ex�A����n����V�o���hSۑ�����{����V��줗J�Q����7�����Z��,Nm��b�[^o�ڦnJWj��͠|>g�-�H>���w,佟�z�~Jʯ'��]C���57B��`�ч�RVJ�m�r���:T ��5y�Hj��7%	��X�+�0��ph@~�cX���"����~�AU��k�P�֔ ��H���	ay��lċHR��l�#�L�A��cu�fYtVs[�`Jκnoi^����p�/U,"�����i��+	�-<fV44EȜȞ��@a	�9|��*"�'�t�p�2��q3������A��qˑ4#LL
{؎#$5�2�2ؗهp�0���q�t.^(�Mo��a�	`��G�v��/1��V�k���`�9k�Ϫr���5�.�K	���v>/ytR�����,�q�cKY��0� �og`�N�F�{�3�T:�պ��Щ
�����}����#���E�	�\!�&i9@t�͍��oYpp3�>��g���*���E�a<�<�zR�&蟬aXHZ�'x���oh#�L(�L}���:�-��!�����Ce��S� 4��������P�]1�Gw����qi�ᴓ�Kk��c;��vw_�ΌB:�'P����z�ΰV��Ihs�knF���S��pN���	���	|�cT�v��4(֗�n.;c��6�#R]G�v�nv����Z2�&f��=�)���	�U�"����·u�}d�L����b��b��~�⺐��n������c���c~+�����BL�%A�S�ѣn�rU�$ ґ�7U�?���!�{Ig!.���;~'�6��t+� ?z�����>�?yi /9�wo���T��u�p��,f�:��|ܾ���C�l��].�߯_2!I���U�$���y9�O"=�#�)f>	Q�,��izy���4��n����ׂ�7�������/7�eQ��Cs��m/�"�e�C�笥O�[H:�ϗ��M8�E"3# ��\��I�����R%x4OM)�i�iO�??�n�^�(]�(GI�q9�+B*-fG�Տ�)ЭC�N�U����I�\�Т}D�\Bpn�V�:��1�¸4i�������&�7���t����yU�$�%�/?dD��bx3h�L��/G{��^��j��;	��R�c�{<�>>G�	��*B7�M�d��K���e6��ݣ}3����9�9AMJ�K���T�Br�6���û�k瞁K��qg�L+L��w���̏W�)8^��NS/���Ri�ӪӮ�W�{Mյ~Q��N����'������?�H�aIN�Msmr�s[�Ԍ���܅d ���K��E�c;���MR�I�GlGe�h|����u˗��Rdzw�=
��c��E2�0�ZÁQ>����d˄;�����+2˼��6��톖	��pA� ʥtޜc��t��zq~k�x�l[��R_C�@ۡ��a��Bi���k|휼pn�G�m��`L%_��ݼ����]�yJ�h����\�bD�h��5�%��r��]�nDq�b�=�P��B;O��oI较�6��u
S)��[/� ���:O@��I�U�Y��B
�c%IA-{�#���|�KN�%�\�U7:�7���
�e)�6�]1!��voaJj�G��㘯��&���o܁@�6�������F7�>,�&�&�����j�e��"��Q.��D=�+�0%!J5�j�7�j�r29B��z�Sq�� h���?ɇ�������L�И�h}��)�;����t(=\�]��(I���v��AW���X�Q8���T���P,!d�0�d��-�^wҁ=�]�'=�l��o�R �D���q,\�u,�qB	P��Qs�.7�:I���6���Ψ[�ڍԧ��>'PKxS}4r�m]9	ʼG���2}������2��l��-�)�l���w:@@�XC��/0���Қ�6X���� ����:Q���rȭ��0��HU��z��Ŗ4�͕k8�EL�4��&��0R+�z��Ѹ�2$�\#�O^K�2J���Q�x헖�TH�<�T]��Nn�b���{����W�"��W�Ǹ#(�>aE q3�\\ǒVB|Y�f���i��U�&"���)0�ȷ$p/d�^���]�x�=�p���!g?s���k��*��1n�Q c�D�� �l�2�֨�ݛm:1Yc�&&Q�|`��@�p�#����(��}��o�N5����B,������\��f
�Q!kȕ1�p!;m��>��b�<���J�)��]�F�XR��\���Dt3��q7�-�2Oc��P�w?��5g�� 'h2����wE���� �O�rwc�Y�s�����nb������'��RZM�$��\�H��� ����ԡ�p��a	,a���6�[���\��~�M͍��b�;�B�X*�;cn^	� d�^�$c���&S�_Jcf)P4<
 ���]Dc�I{Q4�*���o�
Y�~����!6�8(me į�Ɣ��e���� �IE�����dƜ#��_���4�f��:�s�h�׀�N��_��`� �)�`�y{/�˽`�����8\�!z֛�՞��KL6�n~T��m+���qkI�lb�2-��� A�8�W�7�`pb���9Kd���� ��<o0�?�&�$	q��j9[lHT�^Y(ܭ
$���u������eG�X�xCV<��n���l����uc��",��Z�f�:w˝my�K�H����s��9��m�XkzB�~;���`���6u��:|";�>�W(j�/ŧWl>}�*`�߾о�e�DT�c&+;�u��R�X��ۈ7W�)ܔ�zDc��]�� !`W��#��}S��[G"���j� ).%
��*5Y��P�چ<��΄�i�[!�Oˍ!�~I�P���a���cH����hW����綍6��*���s�0�4����|���e9g��/�ب��A䊗u�[gWu���У���a&�;?v�d�H��FXbL~VCՊ��ͫ0���2���;fI������_��C��#)}9�\+��w�O���:0�Z'_H�5}V��%��3,@*�@�
�"�߮wy��_����%���vWK6�������+}I�� 7� ܡJK�M�<��K�\��?�ВV��5a>B��O���z�J��!���7�*�7�Y�_��O�H���8�䓰`c��	̥T=�pV;^l�%T��w���x�f�B|�D@�~�f^��T�������#X�l~���.ا�'a�6sh�O����-����6ߪTQ�e.��Ag���5?�&�����'B�25�����"��*�RuWP�Q����u�pQ���>r���TP����ny��r\���v!��Z8�ד^�u7�`*�_+y�ӣy�J�����y�w�!�*�7��6�ڲ���< �D
pXhֻg9�R���6���5�y�rc��Ab�!z�x����
�S�>Q*�A炵�s����phS��=wI�a�n-1ӓa�
k��@Nhd��雌�a�
A�#�4�j+_,[�9:���Ff��9����f��_�Z�M�t"�V`e� UK��s|8v�wVjC������b��hQ���	�ue/�y�{��D�S�Pw�f��dx����ʨj��r=��x�hY�S��dj8j\�
�0g*0z���Qfld���B�u���n�o���!�4Ȫ�������G��?���J)��$�c*�+L�k���k���qtS0E$b��Ω��b�)[�>�-�y\�_�1�h5���*T��(�i6qg��8�]��$b
�pLu�10���u�8�'�Yp�q��J"Kn��\lI��ч��.A�%�NҒ)���)ʍ3Xp�Uc�W��$��K�ԭ�u&�5l����_��D�fKk<�����eP�<�HQ�H$t��}���Ta����rDƪ^�D���{��.=Kd;JY*4T'>m�#��*]Y��o3��#P ��KT#e7���
`Ɔ7J����d��[����j����gYʲ�`�#��T��0=������jm@]U5��M�a�Y�����a2��Q�KxP�!X�ߓ=��	4o:�|�9�[�Xc���z���-!�9�+�d�߸_��t7v���0f|3����_W1w��QJƉ`��D����O�S-�ى�?}��,8y���F��1 h; 0����g�7��PK�iU��	�H�{(h�1�&�rs|��)�����C�*����R7
�gQ�e��w�J��� �A{�u!!d ���q�\<|mF|ɍ��*v�vW����kX@��_4g�/}�aX"���Ouy�%'�u���C����o��o�s5T��|Ҷ�.��M�|AD`�!Nр�wn�];���)tlK�e��;��I��M�y� y�<w������6��)��Ҟ��M%g����d�c͕�17�l���?��ܶ�`�n(��c���E=T��P+���E�t^-�(;��aH��U� t�[�1�Wzb']�ʖT��3�C�������+)ي0H���E���mi��)�\���.l�{0���`sF��n���ב:b�� :dw����l�Yc�4�!s�s���{�Vl}�.�)EgJ��m�l6���$�p�Cl�'/ԥ�t�MEjΫj�-���?�I�o�_W�+����Nj��
�`ޣ�{}�> �G}�����+��o)ԍ��+�W�j8ղZ7�.��҅���x	���1�p�%PДt��V� �r��{f�B=�?�A���i� �ێ���0�?�q�Y`ð}�(1~>kIi�����L�w�+zq��1�2[5�k�߱�,OD t�1Hs����L�,�8��j��x��2�`�Ӫ�Zsͯ��t�hlH��hLđ��R�e_Xlk����忴l0�n���q=���&���0��|�h�0
 r�|�\���u�+1T�*�9��Q�mE�ꎠY.J"��:<VoQ0�e�Z�{��L��}R���
�J���gn��z:�7x:�=���� }�I��'�K��EEr?m����v�|\����������x�ɒ�8��j����%��	Gk���i�$�$�����)xu��y>W�I�� i��l�G��KM�O�5�Po�b1�O���N
�V�A���t
��'�}G;\�zd��RX�)�lV.�� ���|+���1]���>�����<�ٴ#.Kiߚw�8N��2R����riM��������m�� ��.|�������^O�V��FV�2&�;g��|WTG��Y�[��|�$��-�L�(�����x$8H	�-a6��~�x��Mc�0��ҊfAG�������8��4��Ѹ3��.oqێ�)�{��(���-D�t���@P�"�`���韒�קz������V1<y�eMSmkM2�4��o8�l�J�͇��/E�
aP�x�Z�ݥ��	��	��uU	=x\?�jw�b�� f�3WLi���.���1�^�C�_%sVP�H�YH����y��*s�?�*yw82=q��<��r�6��[r���$�z\ n�s���J�	O~@M���dn��k��o��,5�)e��gl���O}=�����9��rxl}n�=W>R�B.K��v��S����~И�� �E�z��X]C����obC�"(�~��&{�O/�����,����k���P�m9�bہ�������%F+��j���u��우�K�ji������4,�we?���O���tY}��䲯��x����

���. �"L��G��%���׈x�'"ք0W)Cra����ֈ휜B'}���!�kzẑ�/X�
�u9�j��e,�q_���V[�"2��@��6%��ZE�p'�ˬ�E�&Z��{e7�Ӌa#�����u�6v���ݢi�lU��ֲJV݄J�Ci�����s�T�4>����Hel�h`��(+�P�^[��cvIy{�e�X��-�Tb��"�S��-���lXn�ܺOx� 	8��]vV
C[���*°ld�6XŚ~�RT1;?c��e��iI��{����5�5)=����#HS0}���t�؛����4Ol�.�Ӷ�D��ub�yI��X1��O3xp�1x45�f�U��.6�dL����������b�޷[*Eđ�Lo7���ctr��h�a��aY�J��?��F��@ǳ�T��n �x�1�Q����o�;����jq���'��YFN,>U+��i4��N�*dT�5�<7]��f��$�H���m�&c��G<��1�<i�jw���#4�3�.�gWuj�+�N��'�
2s����I���	�������x�f1ƚ��^�,��'Df���4��|�uؐ�S���ρY�m4<���X�f��B׷�����f��_��6�[q�����o*�4��WB��!iC A��a�>zR��@����LCH���/�<��E�n{5��yo �D��hµ7R�h#�t��G���s�atԬY� �h�q͚����I���IeB�Q�LI�/h)����n��u�K��Ih����)���Dϻ�����f��O�8�q���ɳ�)W��� �r:�o�`N �4�}��)Gͮ�o��eY?;��9z�k:�ރRDv�b�M�7%E���=)lw�j�&�Ћ�����V"bem�̠<���i�|��;:}���֩Be �zu��E��%�q�נm�����z����(a\��Cb�ç�֔�S�͎]CQ�ZQ��+�O H#i=��&��P�ĕGOelZ]x����XY J��[9�L�"
��;mi�w;��#��i�	y�aµ?���^�ͯcv��4Dl�MX���ኑ�Ϋ@=�9�+�������|���տ�� �f-�]�֪{��C܉OE<��K���P�p�|�| (]�����yw���;U�>�FUe0䗵�o+}3��ܪAO�7W�$���*�^�*{`��X�H���\��0��@C�c�δ5�^ɗs����8��'�l�D�ʌ��|�^u���[a_0�{��c���ngp��"��B�h���b���a��$�4�HN���<~��W��aIL�9ʞ~�z��UL���N��bp�_jO����b�V"Sߪ=q��c~���8"���JﴫDKUg�q��E����%gҰD≢�$/<7)�\�b��(9ż��d�~�tZ�I��t(�*�e�J���1��_z"-T;�v_*��q�ٜ�W�� �ҪYI���m'�n� v���P~��	�3`�`��yA�Q��`�E��XN������#��2㘹#�
V%���)K;y<����c��2�/gǮ����v��m�C^�Z�.��|���|��}�U� X;oo?$G���r�i��u�A%�@�Q�����~v$�#WCN!�31��������\5V��:=ҸSDV�-�x�XX��`�מu�ty`��r�ۄ�$���P.�N�WT�@�ک!kɡVL�P82�bl�� 2	_2h!/Z��� �
u�)6@,)d��o]�nӉ�VH����:�hu��-�A��9����r,`L�r �e�6YU�ΡT]	���z�+ �V������[n	u�"�j��N��YzN]W�p��W^�>��y�V��,$�� �ƞ2�/�!����=�q1��87��w��5��)���p+�Ķ�A9i�H9�U�z%5.��2;Z�$:�a3��z�"TL�VLG9�u�o����a4��XJW�~S*��N,:�JW�2U�YHbX�-ʼ'���<��l�x���d�-�C�F\q�wD�]c#�"Q��a=�R`����'���<��'��e������R�����7����tm��Pi�J[���s;��|�9o�9!�.�
m�a���8��`a�a/��m��k�3�	����H%���@y�L�k~+�Fu�\��笃Jr�֜���8���L�2�V)Y���n�h��I���=����j=^��1�>�xv����-rB'`KA�Y�F�Z=}����%�/�d��e��$jqW��l����`�V�T��̔��X��V�?7b��1_4��ɧ�����*�`P���5�ӯT�侰1���e�*W���'�.M�b~gv��Ԯ�5��O�x{T�
�f�[�W��TEHI�c;�`���DM���q2�� # a�X��8/2�,���3������x�4�x+��m,�(�(�&oRFg
z�> t��IB\��h�ɾ�q{�2}�jttv��4{��
��!��&/��<�I���ts�9N֘���0�1Y��-�����2��v���nX��aM�����=h5h�P���@�V�=�̹��je��dz��;��c��˝�$hHL��MY�'��'�ԟ&v�ʦ��؅C`{.S�#Cu�H�}�۔ۚ>��7"�P��AQ�p=��=�(Ҋ�+��˥��cK;���j��|�xVe�zV\Ƣ�`p�T��+��*����V��@�����E�_�|>L��9��1.o�\ 8�r]��L��8צ���/���}�Z�>��ib�3R��NH+��"���܃xC������r���"!�x{em��>���=|n��������a���Hx�7װ&_��c�ʽ����'���{b�
�F���H���V��&��� 0а-c�^9H��­�*�"���Q�,�>ہ� |�"G)̉)b�+L�y�G�C�&�(�8h�KZ���^5��R{�{��њ�K����6�I���^N��o�p������6��U�G;��w�0��Od*��qg�)�]�0��8��H��I,;�W$;Q \�fQJ�,��B<&�@�Gc��Ԯ]�KE^I������Tר����@r��@�����������r&'���!�ثA�_u����Ӂ-\Vd(�*����
���T�>��G�_X��|Dܒun�Ae�5��|�9�B�o������\)��)z��̫���K����T(�PF�O��7��y<�`�K%h8�+�B,����&]��� L���
�},z�7a9�na'��=�g3C�b4"�u,�:��A�O$`�����欣s�|�������U�0m��0�g�Ϫb}"l����c~X��%��/C�)�
�$��З:~Q�=:�a�1/P3����j�Yȅ'"?�������)�Ł�.ɵ���Z�g+�r�_'@�B8]ѵ�*}R�wgq�{����`��eY��}��z�_�@7d�~J������6Ín,��]�e��HF����q�Ęߨ�s��"Eh�?�����\]��5�&�/D1�N�L�����6G�J?�փ��yb\�$�.��X��b�	ӑ��zlɇU塚<B�*^#x��vgk�Ԭ!�p�ed/1�DZ=�2��_�K&zt7^����A�B�v2A?�nگ�:G�e,���l+}F�]��៩Bk��o�K~��S���*ꅅ���3go�[a������ES���ͼ���'�"�Ǎ�P0訢�%"����\�UȚ:�Ir�a���~>3P���.mh���a)���À5�T(�	Z7��q|8n�O#�P�+�e���	�v�/(�#Ej��6|T��y_��>��=7�X�K�E�u�Uo_��@~��wArR�y|㊉k����
��o0�`�ͻ���텈I����|�)1������$���3�5�3��:.�5����u�ֻ(��9�>�Q�w�s H��dt��.E���ž� U�������( R|���C�_8	��	(B(*���4�X�|��@���ɦ(KL�IrQ:�W����J��5"�1�)ϰ]��
O��
��H�3SFE_S�w�;�|�;�f,���=N��y���J��RNB&�����gKR��s��d�86��җxA��4��UB�*�X�ҳvʶd�hF9��l'���0��K#0���E�[&8�m�����_�[�u�D�.��Dr��i��m�jl�O��?�16��	�]�� �}�A��S���_":Cp�K�C�#��-�.:��G*PI �F��BE\��㮨I�$��!�T�tQ��~����n�Ȼ�	1����G\�©��H�|ZY˟�:�ʲ��R�Z�����#$���iUF:��utk�0bw�$�?i?�ͽ:W�՗Β�v�,T�K��NA����iHQ�7��֟ԯ:h������5`���З��+��e�=F?�C��2�D�hc�����ԥ�a ��(V���Nt��g�y���D�4c��>~' �k�;*�""2Kf����nw�۷5�jpFS[�r"K#�>��qJ88�®��w<�6��R�0tv�������ӽ���:��Bu����β��-�΀�L�'_�5�̽��7�X1�+H�I�I�Kb�����$g�r�-�j�d����-S�lG���|{h�n��I[^���}������'��9'��Òc.�S�����āԔZW�����b�!�r���e��nM���+2�&��p�;���A�Q���P72qy~�{9���_�G���yܴ���'��mL����|[�N�T8�Z��h�Kߙc]!>���i��u���	��v��k�㚋��z�Ys;�I���!����*�\R �7���F,�_���c]�'�4;C��f!P�:ԕP�am`ľ1r�!bJ�3��Ͼ7v�|��@@�c��Г���QPײ���էQ�j	9	<�AQ�SD"�
X�����g5:4K���/K-3�U�범�̰��7os�Z0-(���1G<?:�:ol-�C�WL�5�j��H�Y��¹�gbs�#Ղù�����,&�K�nr��D��/�cU�p����K��!�н8�P�xȫ��[ٸ7�D��$����f!��y%P=of��Ħ�cv�� ��A��w64�g}'A�Bc�������`�f�)R�����O�j�<@�sqz�OJ޾+gւ'T��;�"��ٻ<]`	agȥ�}3����hH�&3�L��+��l;��d�.���O����?��܍�hZ�G�I)��).? �CT�ϱZW��>�����3k���u�~���Ȇ_У��LN�(�V$����&7P2� ��e�H��v/���7W q��<۪B,��}}�7&�u�4��������S
�0R$uz�˳��:F�"Nr�L2HR+l��uq@��X�"
\�خ%ez�Ʋ@J���X=3u�F,W�A1���Fs"�0C'��P��Æ�]j��'^��m$d�:�V]�닷�?46n�$�ƕ��)���#R�տڂ�ʊ���=��/����P����QO [�˞���*�2<�+F)��8{�����=�z%j��H�B�����6��4��0��|�m��3:Ӱ�.����-ѻ����)��/L3ܠ���N�W.�,����'��o$frX 6����ϯ;���޽��:k����qy���<��>+�W0�"�����KR����}K�g�Q6� ��!���)Y���"�HԌq�Lp�����P^
�%���<��4�JP�%��6�D�4J������`JP�T��j��r�͐^��)){+�Ɨ?tE�?���F�� ��_�Mf 4�-��|��w��h��*u�`��ݲ���׎N�����x�J�4\�oZ��j�D7Z�5��c�$֙���{�s���H�q�ؒW��c&��@"|*�����F~�a�ҍ�̺�����@\%Cp<g�6$�<�F�ֶ�1�g�aX�c�� �����o����V^*����b	7�/�-a�鿿<V½K .�g�����?������Are�����N7���K�D��e�Uq%;W���_ufʗ n��k�4w�Jd�GA,�r�x�1	{�q'1���`�F1I�kR� ��W�y� �{�
�\]м����5b���,2�O̾��j1@��Lj�B�,Ȩ���� �V�����7�B�<B/N!�YM��a��4����ŏ�$,�����+:�=����X;0'۝o~Q���`M7k*>�okK'�u�5�Mc����̟f����S�Zz��Icf����\�<W�0���p vd���m��e&Ap����Fo<6��Z�Ƚv�>�jnTBa 0;S�S<��ʁHCHpw�䇑�vҒ5��#c���/�/��v�Ȓ�Rߓ�!τ���}��޴�
�*,�|*�iÀ9F@Y�m���Q��j��@9��e�N~��d���G��{+>�o[1U��_J(0T����R�v�/�1�H�B
�5�Q��P�7PL�:���D�CQB���ʩ��&O�Y���#51�=�i�-A���aW|�z��5���-��@�����n���J���������.��}�ghͭE3���7]V����+�uԻ���&5��FP��l�b�8���3���z��\Y�E2��wA#�Յ�kӄo���PDl?��|[+-�����>��n!O�ͬ�4���iV[kBX�Ŧ�_�a��gh��e{����������v�ٓk��#��jcI%�5vEA]ž�Tu�X��(��&��J�p�{D�E-���<�t��ng��)��d�N'�H�n��_4*�MF����>w���l;��X�ѱ�U�A�ɢu8��!���̪�ƫ�F�@��5����+%C&%��M!��O��W��_Hj&^�O
_IMe�g?~��B}�cQ!	z��]�A�[ޢ�}�D�9K��7��N(�M ��n�1P�;d>ͪ����� ���U�bT@L���(%�ϒ����s8�(��b����p�>sP�n��s"~a�m@���8u�E� �����W���?XO���qI�병'��Q��s�%��Lj���qX6�g�%U���a%/��ߧ�0�Z�t[����@I�H��$��Koۦ 'yb�_���:m��A�Tb�@.�
���h��3�籚���sj�b1�Ӹ���i�b��޷/
1h@�6ᐏ�Z�0�l-	b6�xupI=N�j���� ���w2��e�V� 6M-�V`���7�Ԥ�aoZ��om)5��ul�!���*IX�H䞼�l�����~Q)c�^�l���d��g����8mQ%'�E�Sq�������z�
G�T�7�E
��0j�}v��xol��*��p��]��m��XǃS�P�o�5
��{q��#�Ԩ��;��@&��I��$l��߇ERj���v�O�P�}=)��FM�
1�FO?�b�3�p�
���~Y����+�� ���R/�]%�.z��"P���[ ����5��M��"���4/�o�k+q�|��sS�����$��O�<�v)� 1��x�
����WΕ�)ZFtM1�zq�l��V���-�^�@f_�J!�{M,|�!V�]6 *��*�w�����2�H)�e�m,%�`$�<��6cIڝ���?C�#��45��ҸI������B{0jv��(!�g=