��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȸI*��X��{�w��h�C��@��D�Iy�Jz�������>T\�)%�$�Ēު�x��$X���d��<7"#U�n�ą�(���3�t�g�WԻ��.�����-�0�NB0���R-n���g�"�pO"Moc}�}X�Vq4�y9�\��q��B��7�V��ӳ�zkot���>2?t1��Z$�������MV֤�D�;ye�t�ӀQ��bN�c���G���=���l��i��Fj�q�}������fI�'.�i�ag�!��̂<G#��Z�%#�Qry��?����ſ���X���Տ�a�40I�G�YDQ0wB%^s�U�rk �&��H�/O�8	�S�����Gq}Z�F�u��C�VM���q�t/�i=i�&+�̦T
��)��bc$���c O��.r��:��\��aO#�ƭ�h�P��P ��41X+�R�PC!��.�\'P�Zr��c>|(��2\�.��tXq9�=���Q۱��p��k@/v�,� t�K����W�<��͑Y:&O���:�K�� ��.��~�㶭;��ܚ���| ��A�g/y>5���`���Lj�/j������%c� >E.k������IU�c�LN9"oI�o ��:�SU�j��M5���h�^���˃9�c|�p�)]���sװ$��fj�2�0|�6���+����/��y���^�*�y����ؤ��7��
�㇒�+gbX���@�%�0N�(%�B� 0���(	1�"�4�1�3��0ja�%n��}�� �Š��_$r��l��3���� 3�g�y2[��j�ߟ�)<�d`���R��`J�:c��Rmn.sd�ۣ�_�NQ�T�Q�!j�i2t�cDK!e�WT���������}$f�?�z�u$Ei�;�$x��)�{���:��j���[�&���5�:2��LΆXDN���bWHN�=}�Bg���xQ�
Q��4>�m!�6
����?-��AX����*��1}']he�<�y��]�T{�̥�WM�F=���:�`�������=�7��!x�X�'&�����Q8)��WxA���ߟ�#���dj^�� M�b�,�ٞ���D��#?s��ˠ��Cgp>�D�6���xiH�3ŵK�J��S���$u����LWn)�7 �'O{������[T|6a���-���X�h�_=�å�-۴uȫ�d6��8�/�I��x�_������s�����i/
�%��#>p�Z���z����t�?
��ʬndE���6�� (o����+.u}c��(���z��Y�!�Ð���W �lZ y��?T=L���<��h�f+FM�??��q�q�,7.���"�ZcOp_ؐ��Ν<)�H����2D���k���nc�J!�{>���|����L;��A���h��KY�����)�jkU���If�A��(2u��p�)f�~�f��-�L�%>p���r�f��H�*IB^�c#�v���3����3@#y�@E*[��ϕ��@;^u����w��]gh���ǧ�t>����}|޻�I���D�IX.4�.��a���K��P-��6[���������c�{#z�^Ѱ��0�woӠ���;��Mmz6��_��8{�o/��D��*��!%��v�"\��)��w�(�Gp���e�c�~��6��׫�
�'�[y�c�H���=��E5>g�z����뙻��&�B�u��HH ���v���!#��ꕰ��%����?�� ��[��VԤ�	����'PO��gJц���/妹�	��8�e0ɑ[%�؀��&�ز�C뻕�⺲s��-�:F�O4zF�8��a���ɘo�ps�� �#>�u�D���4���>�w��0i��*v`�n%@d�y�_.�xNJ� ��IY��Y�v����=�3Z�I���*�?<�
��߻�t����T(�C�7�]F��}t �*�w�n+=�&>���.����xW�
6L�@_�֎��w���	N������c�Nͬ�p��5]Z��q} {>�
�c-I���'�U^�ʳ����z��Kh������ADp�k�tp�b^+Q����~\��M~��iKX\�}E����A+�Q����T�(�;���2�:����|ξ4Uy�R�_�/'O�!%�W�ˈ�&@�少B�'x��z�eJ�QBW8��l��J|�gHH �N_�f�0 ��5=""兰�y7;6�'^}Z{m#2�L�p"�dɋ���t�.�g4�w 3�����{�D��2�U���R�朁"
S�	@�ͽ �g�F,����{�b��LZ����8��\Q32B4�B|݃�SY���kRcO��լ�������;���P0M^6���,�<o6Lu�o�/J�
��:9&ɜ��~M�Bt�ms	��"�j��Qb�j�T�5��2M\uU>�X6>��&�<Oaĵx�$�:_���OذM�%��I,�~�t���+T	?�'�Uݒ�ɉ+��X'&B��(���A�4,�h�6����"������H���ß(��f}�p徤{����ϕ���)��7U��ۍ��\`'���z���� �C�OC&�ͩ"2�?�-��y+�6�p�X�w��N�J�m!5�� �,Q�H]��@G�D(5H:�c&�I��s������)��{�ihw������F��qD�CN9�~�o�u�����M
�)k�V�]%- ��~��yĈIǎMj���;�O�ӗ���g>"�g_�<L{�)�,C��a-� ���!����ǶB��c�+ZJ�t��!O����7�i)��²��>B,�-Z� ��y��HJ $���d(��@g�.�b���Y�!���ij�\%�aŏ���}Q�rH6_n�'�z�zۖI3���8��!f�N��v�i���t 
�y�Fd�'dv���B�����-Ϭ�^��#�g	9i�+����X ��ۡ�Xn�Q&ml�, t�G�������j'q?pS�(��u8��L<����y�xh�z��c�����`��*,,�5%�U����K�S�|��u����oGl.�M��t5/)���|׹&����&���)!ak!<�v�r�:=���MR��>b�Ь
P�/&!�e��:l�ߺ�ƿ�W1!�8c�?d*-AX�ҋ#�p�^�d�F�'�ZA���]]�[K��gr�?�-.�nz*��\�yDƌL�h�����E}ucQ1љ	�c�TY6��NK)��^���(2�0�)
t\tĺ*6U�鿍#Z!o�Rң��w�J����|Ѳ�v��3��O�g��0V�K�b�Y��Gk�q������l�2B���3��bt���;��iJ9�47ԍz��ݿj�Dk�(��Z�̘�A��mܒ�N�饡  �N�.6ݏ{�m���BlȂ���c(��i�j�'���_��_�YF��
�J��-�,�F�xr9�9���(�`$�.��)U�/ewY�H'&�|�> 4�#�	9I+�ֶL�l� �Yx�^׀*�.i�"E�[r�J�K�E'*ǳ��x�JVc���Ƴ����I�Q�O��iͰ�鵻�77��OQ9��('��VG�.�W�� mΔ�����r�ut�)
��� �O�����I�a���ʱ�L]��ߪ;�N+�U��)�?\e=����vC��l�y��E�y��v�MX%����pely��T��o52�
~�|n45�^q6+t?�xL̖��Q-��ys���3]f*%�4��B��D>��X$�`�
��1.���]�~���e(����H6S�S}�0�ˆ�5�/l�uadw0��ڬ翘;����V��2�7����C����O ڻ�S�>���*�����@ߑT�>p�R�[���`{d+&	W�\��$d%�T���D��꘤��P /������Q�ܬ�q�сzI �9��(|8�>ҮVy�O#{/�A.ɩ=y�rC����MQ ��]R���-S��*?����vs�>e� @�z�}BT��.(�X����u?�h�K0���h_Z)mL'�qP��Ս��EM���Kȉh�}�sУ��j	d�Z@U�[p�v���~�BE�GH_]z�J��zo�:5��ժ�-�<�<����#@\T^>N�/��mQ�wZ�Htg��6o,�����!����|�!:�4n�������|gN��94�Ԓ�Ak���0���:ƿ�<[�9I�ZC�^�ZH�`9���g�� _[�� h�uh��ִZy�Rs9oQ����$Lq�pޏt�A`.�XJ1�O>��!	pAv�<����s�ןKz�l�q�q1���'�FBH�<g���r{<���T�jG���Yx���<>�Y�8�gA��`xƊ3�}`[�K(O�v�c�'SP�|�dG�V�Q~����s��tB�Ϛ��5
��OQ���|M�����o�@z ���U��X����n�|�)8�R�t3�Fw��z�������~���������1T������������3	�I��O��fSf١E�e�����@\�W�d�I��Aǖ,��	o 0M(��C<��q�>���XF�F��q�X7�8g�
`n��]/�x�w��_�a^\	�ٲL��M&Ť�ڬ�4sf�M?�ߥ�N��<^�Ë�c�+�;ۇ�_�3��@�G�4����k R����LL�0w��1����ٕ��A���'�4��2`n��?c���e�de�y�b�Zc�e�9g�צK@�=�KC���CEZ�^�G��^���.E�Qe̓�@
�$�@+<AW"�kU��9��Hv��~^"B��5�	$���@c�{4��}K�%d<x���~&/�R�og�|�����n}J0z觉��:D��Ğ/���ʕ��Z��@k��yY��"����	�� �k�V��N�Zc5�|KXM#��2G����	��i�T kc@v�k���'w>�?F����fI��^jI�����_�1,�K"��K�&l��b�q3�D$�zK�Ң��3�ʩ����;U5[��C��,b�VAN�_;�+�#%�u�s	��� ub�1�Q��ٖٙF���T� V�C�K(]n'����j>�Xn�!	O�Ή�
�8p,�O�Is���XI��2�c[D~��U������~3(�`��Y9\
r��Cm�'���2Ge2%c�d�F.�Kk�iT�=�S{����L�7���*�O��!Zfh��wBMK�\��U�~�'�hߌ�T.\�Tp�G=��o�{���_�Z��N8s��e<q%�(��.*�������P�_���$Uƶt�y�ݥ�UDO���� �\Bt�Sy2�{�@�#�v�����T�]q::��@�mL�t�c��B���N��9쥱�2�Z]j����-Ni�c'��?�xO1��G�P���� )y8���(�0PN�Y�t*��\����-��5��\#��Re�k�*,�Q��4!���0q=B3w��)��}���,$��-�XP]R>J�rϻ,W	O��c/7��Vm�RP����A�$��j7�A�&�e�����
R$���P�����+E�4B���*1��>pa���M����Y��/{5o�:�6|�"i����?J^/��A$��8�02�X�++�����t��ɻ����(��
c���o�JqI�t_��`�z��#C�ڪ:�Isj��%�X+؄Zmd��Th��Nj)j��5���0��R�%�S�kfӾ�Iq��!J|m�u��ZY�z'0f���9��fG~N�q<X3&�l����Ke/qi�)�?�>����l=xn8�h����~G�v��ղg�ў��;��vy�l+~�j���OZ1.J:r��X\����\_(��JH?r�*�&�==ԍAP� 3�Yq�^5��pE��MW.�R��#Epo��c9����B���3��W?�^��7�m�J"t�5Ցm��%���R��"�N���^��$Lg�NT��gc�h)�N�W��>�}T�(��~����H���c8����O�~0�V��֟�X��@�g��CG*s��զ]=��r#��B����5vr���E�vH����^��J�Ly$o������s'�ڽ���&�r������G
X����x41K�܀�o��#�R�8H���k�OZ��f��,����·��Jkq�l�aM��|?�I��?>��u�����BK������"9��o�Y�i �����1�8Z�u���b������đ�)7wN�hq穬ٳH���O�'�&p��^�zq5ŔN��v�qĬ1ˋD4���H=^5���~�:���c��C�ؿ
��A��
tsƎL��k��+Ίh�NM"r�� b�f��ײ�b���=[�V�R�r�Ć��f|���xcr)c��,W�I�.h ����c��2�b{�ev0��w�S����W:a�Ie�L�
��G����H1C�5.s�|?�~�+�Ԭ���|Fu-ѰW
K-%���~G.72R�f�r�jҧh�-���$�Q�\�-���#�^6a���vLhsAd�5�������QZ����4Q�oQݹsҁ�g^���1<M
�f5��ὶ*�D8��g���l�cuA~��'b�&D	϶����Dm]Q��A\������2�'-J=�J���M� ��ʼ�+B�jC�Jfk9�!�{;�+��tl�*����T�e�:�8�:raC�3Jby�Oz�^�md]� �����5���lRC�:C��o�IC��قm1��UW�.����{�iFb⩰o@��v0�Y��Л�go���2��h�6��X/8;�
��ZU�P`
��)�ւ�&���C����� "v�8���D��v'�d����],�*'oE2�����;U�+DH���\F3-2:�X/
];�
M�AO��_��	۹ČL�IT��Y�I-m�\���S�5�.h��md��(&[c[OO?/����$�b����mp$�f��Ff+Yvm k$��|����� cz�G9��b�-���T\m��e�������O<J�iX�q:�ƞ8�*:��Cys6{M�	-���}�ꝭa������ū07},1"���k��elչk:v�0�ߺ/ϛ7������U/�SQ9�u/%����*f�;!��3?��3R����E���'���z�㲯�i����fu���Ű�Hi�R�ͅ�\uH;e�����N?�2���, �K*#�*�����+����P��~�^����k O^io�GH��+� �B]��u�����,�o�!����Ϩl��CC�搰9LR"&��4��=<HTA�����=��vr��ɳ�tD������P�Q.��9,畒x���^�=�+�#�x3f/D����9Z+��hdnp;�Ϫ%Uђ-�1s��fХ�3�c�	윔�V�����A~
Tu��B��!����RL۬'z���s���nyl�Jd2��#�0�E34��C��0-L��?��Rj�VtǢ@�c��J��aݮ[EP�q\�\~��P}���FOz�����2�.�����=r0Ԭ�b�zD�2Zaw�����n	��tU`�*f�|�\�ӿ�N�,����}�H����3�-�f{����z%��J��_���ډh�_GL��Гl�Q-�����[܌E� 6�s�C���iX�����L����	�]���v���3̦��-���	��S{Iaʫo�ix���Bi#�Z՜x�t�BńaP5�0�#h܀+y����W��E�z'
|�~d�;hha���4��wbF��vG���x
�V����TrVf�Ei+S�߀�G��O���g�\?vN��� o�m�`��da�ЦV�>�cb�����y+��6�%�pmroq��6���QVu��1U�
"��j5�3����<�Y��UJ1F9�k��4��!R���yƒ����:��Z[:�2����\f��1��u�V�R*��zt�4+�XEë�LQ�H[I� <�Ub90�DJ�Z\�,�>{r,"�RO�j.�Ø�#g8}�JӪ�� �>� �m�����x��#s֣��'ߖA�Pɋ�R�R0b-�5��6?uAߩ]8���2<����|*�T�GW<�(��UwM �&�����4��3"�T*���U	��ɻ�Ѥ6g��G 4G���@qʼr�m�ʥ�l�<�>����:1S��.2���Kn��s׬�Y�XF�v��<���1��d��h����a<�Q�.fT��wV��p�!X�	:�$��@ ���Q���_G��9��7޽E^ٳ��Јi!�#�j]l��rk�������`�W,�z���>�%�z�}���!�,�;YI���\�.��~�1h�t����^}������f���`��Gĵ�Wuh��E�ĩ�MC�L���凪Y2/�f�d]C�?�Ӱ!f�>)#��_��W��]���Y'��4V�����i� Jol��@X�B	գrJ�>�R�)��Yg��!ЩYѐ_D�~1�<c�O���(���ڝi�r׉�~R���iyi(� ��b�Ks��*?�m�*ျ��>�'�г�.��d�Д)�v���	�A�SȾ|���?���P�m%� �Jt)�Nb��s�����	ӭdl�iڬN]����@L�5�&q�0�/h�Mn�V�t�N���B��UǵM/9���w��B�mw�"oE�����Ҟv��dQ�`;�M9��������9�1��|/i����H�|�}�] �@�4+����c-\��zI��]���-~̢W&��Y��Y�rW�^m{Z�a��`P�WU}.n|���[B�_é�x9��e.|K?���ʕ4�[6�),�|m�Ӫ�P"�~BxGƹs�8@F��22HS22t�E$t(:we���`��f��d���M�Q���/|Ki��݃�_j���O��L5�w��:w}�D�ݕ}�h��l��YJ���yشRasp��=7�hXK��1�'qǼ��-|��^��2��.��v9�ͳ�U�-�kFz�y(��-�!�
p�N��'�`p�T��Ѱ��'_)�Մ>Aڗ0)��_*�%h�N]�_C��")��V�����<�D�
x�:s�ϿK�]��ITӖ1/����`��~��yZ\I=�˙�Ic��=<�L�4�.�u�t�A)��a����H��3[VPeO�2��E`l�2���#���&&|Nuh�f�fA3k��5
�T.�����}o���]sݖ��\,@�`��H�Q�;�Ro�i����Rx=���Ϝ°���� ��8�����k�ܚ�)�s\�,�A�>$�N�1r����G=�+z�$��EN/D�%{�W����NT���5�Q�ɷb�_F�)���_�6����h�$�ݒ��a"ԹY)R��Ђǋ���E����	�cw���ca�7��Y�g rA���� ��t��M0�ؖ��`Ҙ)�� ^�lٛǭ����B�Q�"9����+�oNw� �R��P���s���C��=��f�X6}t��b�%�:���a��	6K���y7����L��G��U�1���&����5d�t��ƃ�!0�W���p#w᭏��V+~%�hI�Ly8W{��!�x�QO�\�&ƙs���`��$���Y��fb�e��n�2�Ǧ�)xvʠ�Gd�q��#s��H�WcuԵ\'H��զ+<��B{��#(���>O���1��!�S%.z�y�R6�e4�ʡ�[�S�ӧ8O�۱�Xnjg�$�c`f���7��0��/�W<jN����0��+%J
b"p�,i�JP�4,W������&��f�s����$ԅ'P ���	- �2a�?����r
-�7����GtܨY� @�m=,�Bhs�$hrL�`�l�y�����LS[:�K���f?w�w���ʎa\a5�g�k ����$�]��w��|�g�*;�h�g��843�ߡ�mOP#�z&�9j�GK�����j��[�*���P
m��e���Պ�>���r*����q�X# XT�?�PzE��-��4�J�`fa��˴rNn�@����&V4�8���̯�Ȏk�d	��NJ���O�?�/���L��p_L�?P@�1}򨞗�f�`��=ã��bX��	������@��ڔ���:��Y�aPk�˗U�'z1�b�8B�� n�V,��!����ҏ�>w��J�R�U�?����<��R�>�7^��M��&�F��d��į�����d�\��n4�qLph��� ��][N<6�=]룱`�[s��}�n��.�>ıT��)�[��w�Ɣݝ|��
C9�����,ϊ4ꆱa��Հ���EiWQ�� 7�U���*h��q�Ι�A�eٱ������Q_w8���J/�_����U�Xf��j.M���i[~269=!6ԝ�Y)���9�nao��O� �G (!����4c����&-�	�h���̆I�ؕ���lb��I�0F�y�t_��ZG.��a����>����U$?�'~L�_h�r�E;��-E{MK�5�*/��<^`�q+<�s���|A��7���Yj ������7�\� �e���! ��]�Q��5���6?t�/aW��$��;F&4(V�B�{�+R��{U������: 
�Q�_���H ��KFʘa�]c���	�0ُ���x�P��4&�k�-~�K7o,RU�L&���M��#�G+��9Z)�	�^+���J'�Z��Z�>��i�5�-�+/y�Z�uG�ꉭ[���45VWE���E�;*�� �ߖ�\
�~��y�f�/U�D��X�R��M�<��NNA96	5[�"�����B~(S{"�?]W���
sVL"��_��n���M0�M3B�+��+hOCR�>d3R�R�Y)����_�����B���Z��`�}�:�VM�#��1�G��\�?$��~4�]��v��1�ڥg|� � kj��|��m{��PK����PY�Ȕ�C#����`�=}��^�G�v@�������C{yq�zt�$Y�|�quϨ�7����+�]�ף
v�])���ԉYts?��eӬ�X�H(�_Գ�͖����-�ܳ�O�ᾙ[o�8�%��Vɦ�����k�QTg�FI�P�23òGC��U�\k��������)���y�{/C����ۘ�vY��/�!��Y�������3���b`ԲfР��[�2�C��ge8��+�6�U����LK8��H��P�i݈�j���'�CqZa1ۂcS9���y�as;��N�;�
�}�O�q�IxI��.!���\���b�֗���o����`^A#�5<�/�Q>�*"c����z,��f�u�O�ϵ�դ�gY�G*�^@����,&�R��]�bqf'��C����󢰧ϔ�%�fڭf�
̀+���P�[��k'%vG-�}����㏧�ȣ��ؘ�_�H�y�cW�5ZT��B��Y�4w��8֪�a���&h� k��z�j;��������8����2�Q�:;�AGk�j )�-�Ղ�W�@>�=�C�$��zU5�a\���&k�Jݿ��{�"Bo��d�<З�%�#5Cl0|FD��˵=NQ}�/�g.+��W�H��_���<K�uO�X�8$�/  @��L��_�!�>)�~�Ⱥ��}wm�J��,Z��0�;��}zɧ�^�_³>�5D�@����;%�!�y+>�#PD�RL����U��"��q��:3�b�u�?�Q�Q(������p@��z�402�ƹ�D�����C��
��t6���C\�w��z�Ґ�z-��K�_����f�}A�>���3 f� �#^�K���e�d�<I������w��W��Đ"A��8f4�*�/r�N_�/V��;$��S7�|���i2=m�Z\c��%�QpAt9O��jr0�o"2���z�9I�����d�%%��H����� *�<���%��yuW���ԏ�}���q��]�N�48S�� q@�Y��TD�}m9Q睸b�.f�aT�0�2�ܝWpH9������
6Kj�گ,v8���4F��p��)��H����Sos�2>]���S�>s��fz^�v��~�}����Сd� �F4��B�(�>�Y	O�����/��ا�[U����S���I�n�b2ߜ��ږ�`����hn��}3��/萹�vK��s ���IL��I��h�v��K��=��e6E,s~*h�c�#�3����Ў���:!�&������h?�[����/�|�DwQ�6�@�݅�,����HG�[36;�����_��`����x�}����q��0I8�e;����kG[�}O4V ]����JFxŰ�IK��T��&Z?�א�}.�sY����Ưa� [`�	�"��>�&���Zh�� .Ϊ��*�X�t�*IRC�"C��l�0K�jSI�W��'q�yHM���f��-�n�N��t,��HU� ���ʭ2�~\�a#��QDp�[�hRi�zI� ����q�Yǲ���ܴ>ɣȑ�*8"~�y�ʒ�;7�u�TXەb�ʪ�f$��Gg���v�����8�Tw�0n�A@w;��*�P.xWʕ�c�\`��Xa�$p-���h<[$6d�3�!�2B}�O�*��8��I��"�;�t���o;p�R,���<��WaZ~��^��Ym1�,T*�x8��/T���W3��[GA�lW&K2n�5�ɮJn�=�9���-\��7�-t�tsp̹����F���+�#\9����].�h����ؕi�e -B>���O���G_�Z�bw�в.H� �dD(1Tғ��V˲��
~�d�����O�o��T|5��X~S}"Q�l�EBX��f_iG,:�حJ��Q1��YB�0�=�<3`Vl9���Z��B����T�@�����[�hL]��\�|�Gi*t��n��?�G�������
2�[DZ�(��6��ٱ��m<\��U�U��GSMd6��S��T�I��D���ގ�X�����=��4H�1."������uX�Z�CK�ƕ_ g�r�eM9)��8�,�N�B9CQ絟A�Â1$Q��0;��YJ�#	@�~}�G��f��GS�|�&�c�N�U:�c�S������LpW�]w" S���w��d��B�I��NH�޻S)��v�mU�$�l)���>$��H��.�O�g���#'�PIW����d��]߂���@���dG�7�E4��f� �?z��Q��w[z�Z�#��~@��fx���-����B�X��j{#����z�g��i�y��*��I�
6��ݒ����XX�0�hj%,Ȁ�iW�̲(�3Ѽ�Q����ɮH~�)Tl��~�R���j�z�M]8������D�_���x5�
i��"���s�:��c乩w�
!sI��P�}s��1�-f�d�\A��4\�1=P9O���W]��&hs�:P�B�2/\ř��&:�i!�Oi��#q��j�)K:���y:��#���H�0z��"�� �CW���Ŝ�6&։���鴄�.�s�S��^
�tk;�O���N��.S�q���q��¶q�d^�a����;y�������l~�g:�8�g� 3�գ�jͭ����®Wm�m��.ca*|TY���x��)ɷ��'��oN3�M|;�p���҆�)Ĳ@�M�el�g_~c��6L���JS�������T�g�g1��;2�l_�;�;���Tq3����.1�Gu��'Axl}*��=X���$N-ݹ*.k�]�T�G���j�}Z�[��!ig��d�����Hp�%���i�,��)��0Jc�],ű��L��F��佳 w�v�8|Pn�c��a�ok=/x��d�s��]�Y?U�i���d!g����Rt8�"?�:��lW�&�#`��+��������I���F�Ӷ^'`�Zmlh�}J���L��{�Rw�%��P�4ճI����:�fW�8p\+�G�� �#U�� �@�3�^2������sa�C�c1uj'g�h>��f���@Z�̧�A�;�<�WC�h�I;��Xi�R=�^�[�Yq���#l ��p��k�y�S˶$l�h�Wº�J[�����Hu���X8]i4��04�;Ҭ�A�%��J�@�cnR��Ծ�nü��/),3ȞޜlrFY��aro����,�
��x�f���Y���D%�
��!�#�<����>Li�K�����&���`�\2��6n
5�#�)��7�].�K����[��4ĩ�G��m���������e�p.A>ih�K&����R��ȁ�uĽٴG�˩7��U�c[yL��89MJS���� ��7f���ov�M�"��74�t�oφ�K~������&0�7�Z��|�x?�c�X(>h��}���9��j0��0� ���zad��-Me7!C�>b���Te"#�r�
-�T�?ɨI��iQ#���M��>o�6�F�dw��V�O&AC�G�&����A����_�3��������W4#��3���^�:$n�̧+u�߾;��k��P���4&rR�r��?t;2{D=E�Q�d�;���$ƾc��_>(��� >�h����2�N�>�	.W#٧W���L4a�R�`�W5�$Mg���pmC� �U�Iʓ�܀��-臰���L��p��`�c�ۛy�>y�H���o�K���Z��m���͗���w�&���n��
�ksω@o�p�|d���yѻ�R��!����҇�z�)��
ili��8���V���ׂ�¾6vJ�Q���%��]M�0�f(P3�C��L�|��a
�:�!K5��qy��?��#`�7� �#e�̲zfK%�r��Cw���m��"��e�-��ܟ���������^p����d`�ȭ�w�|V�I�������:4��ꡳ��ǐ�ܘ61�I���u�<���4˃`��v���/@A`�H��c.)�)��w	� `|/�0��b|Jp�x��z���4K�8�b��zRz�C��b����}V:�Ԁ>��=� �\���P��GR�w��rӍ�VE�����؇NS/�cȐ��G~w��c�}�,ƍ�"�@46�^���>՗��y��W�j����s�����^W@�����,ط#�J�+\m�L�#���N ���$��-WM���V0Rm5�D�/��W��U�/��R�%i�<���D�N9�<��
l��Է�C{�A=HzZ
���Q��_�1^�<^� �(����1��>R��P�VT�1Aq��W"�4���2�f��3�6e��mi�DFʑ�uo�ꩯ��-�,�oNa+�k_�5 ���A"��d��5F��<�37��r[pb[����T� V�5��@V����c�!B�.}��0��S�1��Ѝ
)������}���b6�f��P�Ӹ~���Ǵ��-��o�ZMP ���݉B+��U%0�3�<y�����o�ځp�!˘d�S�}��+BL썩?�_C��y��m?�±���R�3yZ���Ќ�6A�����ߡ�霙l��OcB�������N/7�u�~�;.�3'fO��c���$kB�(�*6\�.}S6��x���:!�����eb�D��)�=�Y�Z����h�"dSzVa{	������ڏ�x�l����mZj.��%b�����L�1(X��вد�%l�x�2�נ�"������^ʈ�Sƺ�+6�OoZ�����f���֏��0�C��ɴe�Yν?��E%9��d�x>>�R�"�lw�Ϟ{͘���� c�ۦ��!=e�τ�P�~���Kp�H��E�JX���W����_Ji91�$C(S������Ѥ�vu�f��e��LWy���&B�!��R/J�fۨ�s������Ͳ#>k���D��1O�9L�8pCm���ƑX�k�1�Lc{�h$.���1Q��_yhC��nS�d��@G|��fΖI7������ѿ0_[���嬶�_p������̹��)����Y<�}gkݹ���'Y����k����%�T���nH_���q�y��%ZaZ m!/��.#r6k!����	H뤫��g6H����ve(c��3��ҩ���x���8NĊ5�fl��@$}�.o�h�2���s�1VX B�S�V���S�B�眂+��[x[����r���<�� ^��[����tQW����c�[)�Ӷlc[�~�dv�����h���ݩ�y2n�I�*���z~��O�7�/�r�d������
�|�>��X�@t�ِ�Z�l�z-ž��:�>]�u���IW�	W4��0Ѵ��>���W�.�L��|�2��ݩۚ)iV�,��]-������ư���~`�8&�Z�F$*�Z�`3F�S�u��PZ6�V�{h#�G� �&k �8��;�s.MTg}�?�� N��n0R�* �s������i~c�J�b���Y�y��*�6�Mq.�`M��EA�VE�.��oa�f�~%5	#!�^� �ኧ�����	d��L3����%"�|���N]�Cz.YC}�O~P���"��'2�y��t\7~����3��:h5Ah�*J�U�3��-|��)B)z�Ϛ�s��2���ΐ
�U�9�R�.e-��<xv�T%�f�%-��U�B�>2���gS-�d�����?�	��P|M= 1�k�Y.2	3�`�UR^��|��A�������C��QRǡ�@���q��x��P����&w��VP�����F&���Ϻm�A�|��GW���!�`�A��	ڇr߿��o��X����c�5 �!|^t��A�i�D��h[c�ϐ�R0ݗ���7GK�s�/��t�	�8g1�Qr�b����	�ѯTL}�j�R���,IƖ��"�ߨ��s�p}:��s���k�4�N��O�8���\�M+�����k��ӊ�@@���`�;g/���X,fXA�p\�qz�$��#)F�@����v�	�`ޠ��
�h�M�B�&�߁Ye$����z�V
�-��[^4���%���_�Z��@��l6��nRG�:�ɈW����R9��7	�*c�r�y�� 1-u���@42�X'��Dy8 ��5A�U�9Bvطi�2���t��ԕ��l6 g�����g��.�S	�]JR�f��Uw�B��w��p�B2,����R�v��5N�=� �`Tۜ+�х��(Y%�[�Qvaulhz��W!�*��M#Eˤv�L�C����&�Vm��%��ջ�&����>��O�����Ř�%`'�������4�4�k��u/�MyO�$6�tр�a����������ڣ�b�.}>����
�l�L\b� � � ��t�����&ᢧ��`xn\�� F���{�&��ي�o�[D�� �mY��t��D"J���'��됑T��{Qs-��ӌ�^��Y�	��������)�Xp�Ȼ�z<+e!�.��^��cW�D��|ּd�=]�0�G�~LL,�0r���NE `�h:n����u�*R����sv�-U�RAc�(?��v�!��+�Gl2!�h&b�|n��B�����!�-�LEx��>��_!2�|��X��V���s�/��"��ݖN���D�W��?=:���x�0�
�օ@I:���Ǣ�k6�6��櫄z&,6ԔY5��@^��7�Q!%L*V�d��e��q�k#�N�������Q�C�:l���dҀ(U��<FF���@�v\�E�s�����b��`k���9CQ��h�X�ȓ��q:�hp8nD��a��|v������J��ї��Q�|���&6`�C�V8�	9_z�%Д;�eK��A�z�ڻ�N�莩يj�3.E���m) �O�G�����H�2��W�.��5s�.�-����hd��j#g�2��kVʮ�~M�(׉��瑷'�e�=Q���e4��gjP�EK9�S�X�|	 �-P�s�$&�}�Q%@�>����0)de��i"���	����3x�p
z}�_B
��Vs���6<�v�L�����s�R���{�ݧ#0�����$ꀼG�|�&"��+�1���cD
�����1u`N���K�d��/�Gj��a|ћdH�pd:��V�6����?�[sQ�r�rzg�g������0��W+n���IoT�=��b	 �(:�],�9���`�+dRS�/,j�~�{�24R�FaU���T���ݲL���؜�\ouV��bx���=Lj�>��l��&���\�K�o���R��$���w��6��T���*��<H��g�?�w,�j��`��/f����9ߍ�v��qM�)���8��h�|�(���h0H�dR���H3��BefB	�����r�ԡ��.��,7�����O&��v��rt��rӳ�E�٫&,�s�[�h�m:,
�#�}:蔹�y�&iׂ~c��}nc��[�8��~���H�o�~�lyn$��B��.zN��[w���wl]�C�\���Vrɟ]��D@��12��S�b�q�W���[����ȱ�N�	�H�G��A��:�&���M��Ʈ�o��P^������_:���
�i�&-}��M(�e�����.�!�UJ������7w��:��<F��5S��~0j�'�x�u���y��b�81�A���C�pC�U��*�8)K�3X��]��.��>_l�&�n��,�	��86IV?�D����f�y6����Ra��҉�XV�g^���]	U�|��@��Rô���I ���m4b�2�T%�ڛ��y��}�~6�\��u�yc��T��ۗ+)>�iW�",�9�pJa�\l7�ӫ�В�V�!�Ԓ#��̡.�br�#t�(s6 [�ܿ����+�Ծ��wM�zh8�ܗ�hNӭ�QMx-	,��<OM�j1�uar7M���=�����Ȃ�eB<]��Jm|�9��5?#h���=���hK~�4�I
W&=!�I,��PMF�w���Hz�u���������t��)]�5���} ^���C�� H���Vz���[��;��gՂۋZ�x�gv\kT�Q�YP]4mZ���L:ɪu\ ��"	�\�^u��gC��Vob��F�a����xyi؛���#��`���n�W�d0M�_w3	����u��n	�p����tL����A�Ίa��:��`Q颈��0����?��Q�{;kV^G$ؘ$6�M.��,����V�e#Y�����#��E�꨹�Ca���!Ԏ����\�Z�i�P0:�B/�}z��B��'.������q�t,Qϖ"X�Ȉ�M-���KW�\"��R��˚���K��p�rC+*�G�Y���K\�c��uɻ+r<�pH���4�.�99T�C��+�,��p�:��� ��g�D��\���A�׬�r9�����HM.�]+:I�{cg���&�Y�8~�a���"y�����i]�}�ެ@��:9`,w�L��/#����$_� �[��gV���)E��~�/M�]��Í[4���GJ��8�j��*��Bqgrb(U8���_G�!��9��E�/��P��&������ksʷz4Q��	~4TWsL�@C�拊���b1F���[�,�$I�IM�Q�XN�e?	���&��|����>��;"�]�)]y������Pif=���S��#��bLg=����G�V�̽a)[�̱<�}��^���0`=��$����޺�GVDp�3(w��pZt�+�$����z����2����x�s[}A!��@�45	"@�{�d�2�{S����#
�@�ZH�r,kG�!�cl����}��}W���k�1 ٱF��kWJ�!(fw~����Yt�FciH�<"X悎��DVT�0�_ڈ�Д,����ށ5�3��"W<�5:�ĭ{c�)��fcݱ�.���)t'6���[����6|�Ji�(�A�y0V��ճ�叮��YK�{"0��s�/Љ�����LG��5g���йl&b�W�������$[~�SuF*���"�oX�Xm8�}D�I��5�3�,U"���$����6m<r-�k�?�d��v�@ORY���� ���I�f��OD��8�V�y�FVI�=�֥�Ґ��54A�#<_�rx�+����e$��]����_Tc��/�ᡫ�;%�"���Ƭ�i(��!�m���96
g����fl�v{r	d*��h~~(G�+���*�V,dDY��q����)U@>����������̰�{��-�N�����%�!��F2�WcI���A,�p:�T�)=Z.��C����;�Ф����bJ�����6��9�#���eZ��=��Q�J2�k�ͫ,��>�m�F��BF��pf�s��FExG�f�s����S8	iy�0 � �j>��z�p��׳���OW8�9��`}�Ng¨�����˨e\��u���5Ro�Z`p
�)�i��p�G��aߛ�-+�y���	V�����O쮩�'��n�t9�0U��/�K���s�!	[�y��]։��ҋ��7��Q�՛E���aEz�Z�3����}5p&R�6f���昹�8<jD�N]�����N�Q�Qq�n�
���*n5Ͽ�n>�HC����W���{rU]O$"�~�1��+�42���cv��4鄍�r,��7�&98Vi�d�"�I��+��� 6��]�#�#��-�#�B�j�q��"܌jR��Q���0+�f\oGi4�{K�86ɽZ����q������d��D3DkP�%-<W� �jh����wo��.	� I?jӦ����b�_�1&���1{�\�:@:kR`���B̋Y��!D+	28Qg�|�ޝW��<�6�d����+��Nk��h)��[�t��|׻	9H�ӡιMVº~�Oq(c���T�к�oO�1�15�k#]�n�R�g��0yJB��T�O�n��u�}��ȩҪ%�(tжm�/��'4�>딂z6�O�ڰ}�;�y�q����,�
�Q���K��D��jF�mf���:��+����$��B�&��٤����Z�:�p�5B=�>
�x
D��n�c-�+��bu�]��?=`x0=�=$a��2)���2
�RM��)D�`�*�Z��)VC�������=�
��E5�z1*e?�g���k�ރ�z/]�����>�V��ҩb���,;<E �<{�W��ܺ�iw%_�٢��D���Sg��]�J�,g���t(�tz���7�e�c����(�5�u�XE��G2�3��cڋ���2�����u���c�ᡭ�m�6ZAo�_�b+��_e�R��kG$�e4�=q_�(uv2��L��J��*���6�үT�%���I���=F�L�Ά΍-1+r(�F�?֝b�4��92
j���CF�1w�C�Ul,��D~Xh§�:� ������ �q�����y���4�2̍ś
8]�F�f��_p�k��)�U�2�wH`<�P�<}�d���nL����ϧ ��r+H�5�}�����[hJ���玺<��J�Dg�y!�4e��]��Q�ÎPPݐ�t�_-�=�����@|>��*���W�YA���<j�'L����x��ٔt�������u'm���d\g��9I]/7��|6. �����_+"=Fې��qp}͇�h���x���ew��B@�=3Mv��A�ߖ��6M!�s��c'6X �C' &��GS]�ͼ�n�Q6S
aP�^�_�?9;/��V��5�=�a�ׯ�:2�w�.���̹�uJ�v^Z��f9]��i>����r�]=T�#���*�GDE�����n�P؛���8��W�Ҿ�m���A~����ۆ�2<�I��!az��^$�%��5-O�t^��i���m��WZN':�*H�^f��K���C'�'RM�טp�dAƈ4b�wT.^q1]��ey�o�cJ\�� �0:��5h�W�+�`��\�,����Wk��f/��<�EnӼ��<p�،��L�jj'�&C�w��풼*,��YRL��c~B��;Qt�R��nI�V��@w�����B����:H_� aK�W����rĔ�4�	�q���1�n�?I({����9h�)tLg�Ռav���ӒQ�O1eϮ��`=g�M�z�[E�'�e�R���FYX�NHl���R�����7�q΀7�gH�w�g���vI�	k�v�R�o��}�� �-ʇo�S�5�f���j��1� ��cX��c�<=r/Vë�3�,�)q��l*U�/8�����]H�5���V����d�ɞwb�nJ�j�!��b�����ZRZ��|�O��8b��XmH��nN�B��ů�Z$�:(t�\o0S�$�a�����>��{�̸1&+U;drh�{�����Ԯ�U$[����"�9�u�qਙ��9�@��Aof
��L;p�|�(�U6������9�jV��N��y�����g@��z�I��0mG�n��X���
Ԭ�էkZ�-B�RD�;NL�%͵��u�V�R�u)\�K?6\��f-�H�wB��.1l��m�es�at�U��\�+r,��s!����S�u�4�t�C�J�N�FܚE-��gyM�6�R��h��_�:�,��ej��R�CQYs����FC�T`OK�<0�i��m���%Ԃ^.ZbT{��zOR�I=K�+wQ�	l�bE3xle��P>���,),h��a����ЈC�	�{g$א�)��2[x.���G����������2����-��$������ns�E_!{��}�0'M������[�k��M�r�!u�7�F!�3I`��
�'TU�IVU��#f�t걷���9������%�[wЦ+���M��_��R���Uś�1��fW����@�\uۘ7(,-�G�_qs�g�̏d��qX���ɝ��/k�NZ>���G����Kј��E��x̪pH��2��ob�����Eg�/a��%�7^]��\��B���H<6t$P�ێi�X�zc�[�@�c���g�?H��ѧT�I���}NX���Iŭ��+b�;���[F!4�j&2�!�&�+��Ό9yK����%]o݌� �Q��z���srA�*�����T�$b.6�Ug+��4�`��OU`�D?����B�q$�/��k�&�0oPu$m >�`����@e�3�#�"�w��#���V�8�$�x�����ẽ���V�0㇨ş�X��{}��
V�]����"�It�[��Ztʦ!�f����x�}cN憩	YLUy�Gn�M(��wr��S�Oc��{�]��q'L>3:��A��d5��ˢ���L
���m9����jM ��J�Ͼ�پf��k�ţ�Dl��a^k�_�OU; ik���-�A��|f[�=��N���u��	�V6ư}۶���X�h�m��7E�q&[g���&���H�͕�=d��!��+($��g��iy�]�;� �]������4��Iq�]g�X�%���WXC��;j�dDv<�@͟�M]����q	��`�޹I���n�jw% F�c�]���+�@)�I�e���P�@�PR�d&�oW@7XTGl����Ԥyk>u�7�d��F�W������#L��`�g_{�P�U�vc�;�]R�량�1+����o��{^]��\Hb��׷Q�!0��H8���y�и�$%%1ٿ��"V�%�[�R������l�qM�Ǧ��G?*x�r��I2V�LU<����N��}��4���Ob��� �����{�Op��ewVڿ�����8^�6��s�>�/?-��d���}�k�;��׮t�ӿ�uh��i��a �p��� ~#�',/_��l2*�d�BS�>��ns��~���|{\�š1�̉Uov레�(�#��6o��p���L/��Z-�_l$D7h���UOp�� z�`I-�7���t�����&��ik��^O1:}4Yh�^6���9O-'7NFԅ>/�C6/���t�����r;���h�5m�9�����{V.��}��D�J�ǯ/��������>���.���T/��!��yW�R���Ayd[�v���D7�s.�XQ�0����D�H���w-l3J�Y��)����8e�E[."�A��_���kTݧ�<���ٷ&��Pp�#7�a��V�E����|~$�_sS
E BJf�Δ�D���;m0��y�z�ָ��6{�W��q�	O(2�/4=�k�ͅ�E���%9m�n|ܭ�����5�^�I� 5�>ܿ���َv��}^)| w���Z-�9֯�]�T� v�%_�������XZ��S���y�v� ��=����O[���DLGwJJ�a�wݼ,0��)U��xqW���pN�]׵� �N�L&|��?%3�-��L.9(\ii��Ȩ	��I8L8�����htL��V15\76ya������3��e��d��>��>�T0�����n7<��D��U���ǚ�6_p���|����#Ũ���^s`���Se>��5R����Z�``�p)�x^]Q�̭�1�R���>�ѩS�#6�tP�N��*7��ݜI<�4ku�оYIG����iҼ�rm����Gqc�R��^���'B?������/(Y9\A>9�֝�n	���6�Xq���-�YD�U�=0�c�[���%�l �5�'ܿ��Q_C�����a\ؑ��bѸ��H�M�=Jw/tZ��E���e�Z�0��Ƈ�W��X�ԅ��m����,B�U��j{o�����}q�X�1���%�'�u4��l�G��_�O�S��4��w}���y�������J��:&iY���r0B��t�T�IK��^5H��t,C�忟;$�C �N)��S�li�%m�-��H�����m5�Q��q� ��
�	~��z��_���*�3`���L�h�٪�]�'��3�҄D��_�#�z��$�L�2� �n����(��|���ô!:d�x���ѵ��Z�oL�b(�K��x;�8�Ѧ��ƣ����xbR���N�<Rp��ˑy=�_{�&q���8�
0K�p�����M(-���7g�^�ͤ�mGh9����=���w�X��\�*)�A2�=����@{h�"c�T��c��K5+1`����6�p&����0�k�n3#x �l���8���I}�Ol�Ծ��y��Ϳ͐RM{��}�-�'�w���� $���_��9�;��D��*[iK���  <΢!�[��O��/u-)��9'����?8|�̰��`vO��f9ڲ C��^�p�^V�k%�l"vs�o�7�d�i�Pv� ���c� �p$n���{I�����K���6LSw�Y�����#�2I�%,C!Tw�L�?0"�TK~�66�"n�ؘ�s}�Q\^EK�A��E6� ��O�O�ߩ�v
	S4�f�&�S������!Axt�	�4D��(�Q�5\c�"#��s����h�:�dR��B���!y>]�F��5�{��\9�R�4{gA�9H�,hP൒�p���P��Z��H�b-h�y\?+rv�c��L8���J"�a��K�o/?4.��/�^��*ԇ�Y����򧍖�u�\���Ќ���>�N� �/1͞�P17�P�5��W)���݈�
'�z�F�.4����7��T�:#}��r�ı��L6�1�1��9�7!�����{�tI8�ZYͮ����K�P������eo��f/���jT\���b�9*9��He5��-��쨟)%C�W��q�C��M�������P=5�R��3��٣�8���
-��)�͕ �֕o�7!7T��tT5�	D��/(�Z�3H	��'3-�\��h��̓uKyv{R[�[[C�'�ׇqƚ���DR��Hq9Jm��~�Y�lPb����&�/��"�+3JV�a!�W2��9}<,y�~�����p�^3�C8�B;�W��	���CyWR�8K�v+���s�K�J<t=��Ps�@���?��?�@L��N����-��ʥ*��K�1W��
v��XN��0҆S�f 꽈���ecB�o�j��>>�j�g��K��"�L�V���ô���_��s`��8�!9۩C���D|gI�IIɶO��Pd��M��eYy�s����V�����OGCԠ<'���٘���%�@V�`���Z�&C_t�V�D+��u�����IZ��o��W��ǂ!�a�(7f�����$�����d�j~z���O���H,,i��[)j8����F��OǭN�Q�x�Z"˅��j��g�dJ�m�x�� ho�7O�r�㐊���n\>%�^umҐo�T��H� �9 �����~�p����|q�TI�ҳ�S
�D~�<yG��㱿�K�2e-�_�^����je,�╓���(e\t�V�V�h���q�LW}���a'd�Om�>�*.p*���H
p:b�*�"�]C�u���}�#�I6 ��l
~�u����m���I+��t
�gձV+p���z
SC��+D"��G�Z<C&�a,�����^iѝ8��$[>δٮ���ܟ�KS����|��s[-s0��b��h�)�k���i۱�Z�"3��v���h���bui��h�I5k�Wf�H^?�������ّ�jiD�TD_�!�X\�������am�Ǧ���x<��Y�
���MWU�i�-9��<�R��)��U
Q�+�G��F/b��|:L��J��^!�t���ʸHԂ�o0��[Q�l�-�W����i���l��W�+#:Nā̖����ǧ��U�
��9���j0_o �9��̻W1�0��@�ω��LU�|��>�^W�&a�-��)���ԫ����xc��S���6��IJ�2
Z0 ����E����t��1	���K��h�$��qK����-D���'��p����g�a��(V�\6�<�n�<���,w:~7�x�5t(�Q�DS<�r5?�i#�R��h#2��'��W�Oc�
s��7�}��|���c�AU�ʙ��m�\��:�Ͷ>���ئr�#��l5�&�������c�݄��#�ip�α'(�w�@2L.�Z����<C��A�d�}S�������˔��ߝp��zֽ����!���5ya,�c�A,+�&#��p�;�.v�#�P\3�Ɠ66�=�o��	���y�6��n$�ζh�-"yN��-��:�=�8�G�s{p���&t�]�r��WP�f[��=XfO�@G�����y�+�8i���ɶk�5�Gȃ4��.=)��K�U���YU�7K
�J���[��'�,�6�芜H"����Ϯ��I���t���k����=�z����H��H�̎ۮu*��~�'5�L��ȩ��(��C�5�%���%��@����:B�rm�=��&E��{�3�3�Ԯ�_�a1����s���PE�⤎S�2!G�*��@N��h���cx.��:�L�Ȕ��J�笓Wם���0*O�X�4�	�	�����f5s&������������3akJ�
�����ʃ$��86uQ!꿱V�tǷߠ5�����H~�Z�[�ԙ{��T�NB+%��KJm�}|A�ϣ�5��$Ǒ�-�s�����T�5��zx�TM� 5��L�K��R��+N)���tŘ3��OQT0"r�����c�TxE�; ��_퉁d����A5[(��g=��5Y�_��r�M|$�c��)KX`�wOa{���^"�	�6�z۟��֞�=�h�;�Od�Vei�i��-T�� b��4IVmdeي��AL,�8Q�uD'�8�!�]�Z�f(&�8L���T唛�Uʘ/��ua��*��C����3oɾZ|`B��Y>�b|���!�bߕy����ؚxN�U�,��ܐV:���T�/�TlΥ|���SV܉��Z�/v�wq�|��yHSk�ݜq �X*tnL �F6�HzcI|3۫�a�c4�@�@���M���o�O ��/C}��:�T-�rӦNG��vt��mJ�4/�0�����w��7D`o�ɡ(X#�\,���5ۡ��0x���Kԫ�E2�\��X8l����ag��:�,��b��i/)����A��<��V�߱���@����E.�ȩ�S�BM���rds3/�Ckf(�f�*�7�Z��/6f�T>�Y�;�ML4O��;ν��v��v�r�Ŏm��[�)���j5)���#c��K��g}��Z��9��=��{��������'� T \��N���M`Z�lw=�`8C�Mbu
�X�Jc_�H�}��t�p�v��� ;Db�M��X�4qw���t<�Pf+�A7Q�k��iC�:��&��CVp#}U#��5��+Q��u�qY�^�L����^}}q�nu�*~L�����0	�tf͂�&G�n:Q�),�9=1-����s	���@^p�AS�u��1�	Qm�5��t�k��Ɓӿ��&2
>�b�ED	O,H�	�e����I��tχQ����&�M�,5���p&x�M���k�~߀����[�>T, �f�H�V�e���N&��n�e-�"K��m�jԁ\���1���y�FH��%7=�17�c������\���.��-r
'��r��nwO�_�pJ �ɈBӟ\Z�u���qPE�W����f"<�Y'�lT��;�^)��W�9�����@����k-��4㠨�6)���Xe�WƂk;Y�}���0���f ��*U�(��VdU���6}�ZR\��D��E	i�iq�u+��5)��w�\�>�C	2{m��p9l���K���h��`���^��%C}�׍�Ȅ�`��#�G�	3�dDi;�#��JoqGO�`[V��S��$�{U��{Y�^�I{������e�T�O�Ks`&�~f�#^lri�J�l2)o��f.�"�q9�B;������m^M
���l3��NtF�恴��	%l�^��# �g/P�k������4ϛ��8�,m�w�5�ګ-$�y/\A���8�%�$R=�z�g̮;���{�K3��_��+U`�{U�Q�7Y'���x�lY��h��*��T�ڮ ���X�j=�qw��60>��g��_���%��4=�)�׮G�F�Z�<<�I�����f!+��˞� s$�!��r��@:P������0̋�c������-�r߭�Ԡ5�G�bj��X�j�l�35�i#a��C��FP�2��I��0;~D��x^׆�.���f�����c#b4����t]K��(�A��uܤʰ��n��J�l`����p#˒����L	��R�������Fg��%��0��F-)g�;��	���A� ���x��̘����</��;��Z��mA4lt�q�D� 1���E��_y�9�u��.�m���@fj���.�w�O��V����0 �H�PB�q}I.Y;#D�m��Aɋ�A��9�M�(e�.?��_�����Y�H��=ё9[@'U���I�3r�7���*4�48Q�+�c
B����n�F�	8{no۰LՉŷ���t���2�[D��m,�����)4N/B<��Cf�~�����U��9Dm��D��3�>�GH�8	NW�~�G�
�_Y"�Z_1@�,d��ty�	�2@Z�j�/U�~'H���,!�8�(�	�&T[�� J�:��T��~]|Š���m����^�S��{Ո��(
*�v�"A+�Cy����[�u�`���ɽMYR�\�VX�����Z�B/r�#}X�@=��F�劁��QZ�����3{*x�t��ő�`�I���E��^oXi���I%��r���^6��١5Za��7���2�P�u��M��0N�x��^��0 ��3�b+#P5M��d�P�[�XV��9U�qG��U>�)Jgy��>�X�[�ٍ�
K��	靓Aś��)Ϸ�pv7�����k���G�����[s7��"�d���m�n��>|3r�޴��;w��mp���s`�2*�9���:~���d�s��_�N����-����׻�0�t��l�tLA��2	�M�q#w(e��A����v������H:ũ[ə	dpd��6y����k�]]����R]�+8�w�	��ɀIʍd��mPUL���s�o	��	��)o�گ�\����C��2W2İ�^�c7u���4!��������4���D�X7`U���bB��j��s�T��p@�w��nH��r.$m�O3�P"��T<*��"TL�ŘP�	rˑ�H���T#_�p(\k�30�X+���A�Y:���mp{�,��R�E5e��'.�y�}�}��nmr����,��$�r!R=����J7Eq^�����W�t�L�._P;����ht����+4�Tלv*���=i�b��~�n��z2}�J�4�n	�������Ρ �T5d	R����	�L��}��AWM�4▏�G�8��3�[Z���k���N�¸��WSv�V|U���"ة?��A�*(�SZ����{
D��4�ְ[��N�L�n�X�JU����	!�+�6��w~��C��PwG�r�FUC>�T)�� ��|�A|�1w�KJ��[�ۇX�z����t��bQE.;�����'v���N��+�	`�YQ�-GO�ph��V��\ z�8�x	��� �I���Rd�]�����9�%�?Q��q�s��9�G2����7ۅ���\A��L��\0��E� P�P�T<r�������5L}����%0
�Ñ��*ѷ��\�+����{�����^UY���3t�?=j�OJgaW1�;����Ab�5"AP�Go���8l8���d���~k��,
�i���(�����y�>�3�<|��-����ci����T�9�h��`M�2yl�ۭ��=ܸ��順K/݁��O�2-�Ov�3�A�����؈Q���� �qW��/�,�Ц�U��Mw���麼�S�Ǿ��	` 7l�oQ���iok)��5\@wZ`�҇I`@�G7*��y���m��M���Jx�}IJC�� ?�fþ1
�D�;�y���r�y����f�"��!�g�ƛضQ1f
�<�I�	����ɛ�Z&�;^U	���rS*��9I���10�d���yeaڦX#��jV����%��FAKn�W��M�ec��������>��}|��`lmխy?�e�)&�-��nTw��tzE��Dk#*��1��+p.'�(X�R��$���"Jl�?~��i�Q}��e��1���{��(B``�hǌ�*U�C��;R�|l�ʥ�N�U�tY��`���b�{+�|����:�3m�P⬀M��2q����^��&�[^NF�W2>Y%��u5��7��X�| �!��1��o�)�٥n�R�0�[����ɦ�31�&̠q��!ʾ�Nq�.&un(�9��.*�8T^bLJT�ʉp�]C{N����x"A�]��'{�T�[ԕ����H�g4\عU���]\1L�
�A�@M?m��Z���0��?�N��2�RTҜ(���?av,�C�ђ��\�^��ƃ/M`���P�ŏ<"�E�x4���2N.4� #p�͡yG|���e2	�k0_)��ifg8W����1q�Ļw�fߕ�B �T�$?}bp#5��	��-�pvR��w	'Js��p�i���>)�=���"�ط���u��}������\�95�j*�<=yi�Jc	�qJ��/�
12G�1/���&��=��n^u�
>S�9aיV�j��A)m�Kt����?�D�����I���D�lK�X&�sx�$^�/���0�+��rl�Q�A���ů!G_��}����oY�u���6����;�,�zؼ�g`��nB���HZE7Ԫ}���d�}�/&5������9ۂ�
�ԑ�@B`�i�Ǉ��*��w��{8P� f��������_��xη4wv�9�Svv�r�P�tӿ�B��U�-͡Rʈal���I�'n�O���)�h�&�^/s���3#ѤR�9Q���}� Ւ�Db���6�Z~�cO�O��C'btG{��"�[��d �@�툵���Ӄ<��05}��n{�S
m�Oqq.��������S��h"���f���[�7���s�&�� ���P�@�:T�csժ�(�]�����?�s�c�`��w&�2�o���7d���()�H����(��RD�RqB�e�^��TO�;>�MH�&/^����8�G��Dl�g��%Xp4���#Y��gwd��]����)��P�ھ�&�w�t��r���],��ștZ��b,�
�5/��ذ!��޲��� ��'�aO�)��L��aƏ����5;Nq��U}���⊼R�F��Ku�'�P7��7�C68��[�jW����/�b�/hXЮ��a#���ZaPwtI�Ăa��Jr��|���
%9h�ݺ�C���?��V@^z6)o��Y(�&Y���&>�IS�����9څ�@<#(�Ρ��٦p���R$F����:S[k��dj.
�mE�8=`3�u�i��]S�=�_���Qh�+�p:�.�9u��t_M�(�u�c�Q�3��4/�T�m��E��}�{�>�Q��*���Ȁ���?ᔍGM>c2��(��4`6i[#њ�`��8��i>	B���3����d6B���:e]�����DX�z�.M�}�KI��<�Jqn��;"9#� P9��u5{����&8��&�Pm������)՞��
)�I��q���n�S!m�:��]��N�Z��Gq)�r*[�{��`������9���3�*o`��ʚ�#��N��;SFRjQ�(��o��C�w��r�(ϔޝ�G8�eQ?/��SIc�X�z�vS�C�Ɓws??�����^�k@S<"�@5��y:�y�eR� C�O�A��
����J�X-u���EG�Xmy*cxJ��.&�On1�l��|�w�6���߭�7�o���es;�i����7�e�cV�Z��(�t�=!r�<�>t�������m>˭"DL�p��̛Z��v��V�58��>� X�"ʧ�C`3k�,(���ü�4��H�2�W�$����'�"��ߦ���pj���1�F�y��hH835O�:h�5��%�7�k�"����Ͻ�)	Gۉ�,���Y����|l13v�x�c�R2�Y'��?2�?k��軾�����p\*�
����4�����������fǶ�tc�������A@ƞwG��ԄF]������J
�H�����Y��w�Je�s/� ܅Z�@I4���HXO��ú@����w��z�{rZʴ�\vu���0Ըc�S����?����P'�p�T+���u8b�S��� >߱]�*��Bi4ȸ��|�7N ���G+G�����~m�$%�4�_>��h>H8�o��w*�d)��kJt
�h�|3�u��M��#ܝ��bQ�YؚQ͏ ��xK�@{�V�o�)p��>n� tS�o����5���dI��Q�p2�5�,/岊�Ũ36M�H+y�w��P�������tYA��YӛQ3\a�G~��4pU�:'X�.H�Ě�Eb��nx�����&Oc�S>� 1�6�$�;�����|���*�1�ј��-������zL�,_�{&�D�1����g�g3��/b?˅�H�>)lq��8���PZ�6��@N^�Y1��ԣ��!�؈mq���%I z�ԡE=��ו���d���Eٝ	)c=C�Cg9%e�_�����&a���}z@7Vw�""�FGq��:���s��ҟ����tsV���3�w?+�?r[|B�Z�}����:Q4,?�e��x�� �K���@9���Sg��<v_�V�c9�Wz2Z$0����{\����;��a+9�Q
�sݻ�Mͽ��}��yC[d��Qn�Է��%c�$��Eִ��%�d@���J���Ś�y� �u��J��-��WL�ͷ��X��\,��\|3���+����&~ip$��TڟD@�l]p��l��6�߬�}�{@��
��gh���Oa�b�Ύ�s�)�g#먼�zg�n�(� v�M���N�M�"W�M(�RK���y���u��쌹�����Q�	�`d'��a���!��e�Hp��Q��!�I���ś������t|=��']f��J�N��&��~箽�l����D��X�sR����qT^`p-��k���3[ɼ�l�?��4�[��Lyd@I����?!H	{�~B����&�OJ�
����A�~ٺ=�1��Ϝ�V���FP�	�qȗ;�z���������7�d�K�����P"w�	B]p�oKA]�}�@+���7��i%�/d�����F{���IpD��!���^V�`�衧��=i&F%� ��CD�`..έ��AW\A�[���� v�}����NvrT��ܻN�Xt���n2��anY�7S{7��pH�]z���'�L�_�Rxx]����ǈ�k�̿�U:!��Ȫh,���������nsp\�@�[%,�4E��}Ș���M�%�T�W���>sb3yi0�Ί�aoG��R��8s��=o�Nb >(?S�Z%��2������4�P����I��L��QϮ�(��0�8�!��������B,���"�	�Q����B&ԫ�:8�w�3��=����R���T��(�.C��[�R��K{e�p��zOʲf8�~�(~y�$R\õP)�����+�KW.�=�vG3�����Aĸ�&ui��`c�9�ݑ�i~���V#_����I����9�AQ!^��@G���<� p��e
<ޒ[�yE�_le��J!��z���IA`���bL�o�z
��\��4'�-�4��$�迹8�i�� ���m�&�X�<�����ZRe�0�#S�_��ϱ��I{�q_m�C�%����f4���φg�v!��_N�;Sŕ�LO��v�5����'OYT���'�_�����c��:��L�z��79�?�l����ئ]�Z��,E�y�1�U�i2J��7
�@D�N�~/:���  ���f��R:4��w(�s�Ȍ�����^~�T)=/$%:�v��:���{�m��Rq�k���1��l�am���+�ǭ&��ӱ��K	Lp����I��֬]���eR̉�n꺀K�*<�ʨz�:]�S��x�P*�����:c��
H5J�z��hl��u	�2��3vP�d�������6�]��Y>�hQxG�.�]6�O���)�5:�+����:0���qC_u��/�gɬ���[e:�OaI�vz��xQ2��l�[�z��㰼;������V]�<)bPzz�^����w+���:n�h�^w�.[��v�wM�C\F��b*�����.�i�T��HvpM���ee*���l�")N�]p"�4�K�WT%�����u  ��14�*���^}]�љb�V&[Z�6��]��p}ՐC8au��X=�!��B�`++� {?�THe1���-����&�z0z���*Ң��a�t�c�z�8�KA��٨z�e��;T	z�@w�����d�-6���o�Z��N��ǶH�ȫ�IS�2a]�*����7~w���D<��ćEܾbt�m=��_Q�V�Y��du�S�BU�u�%T�a�M#&N4GVrBw�t����f�A�R_h��g�� �f������x����z��J�n�ِ����>8���d��k5��������y��R:**���o� 8P�5d�$?������q��])�2���s�"T����m���Շ5�P�n%��Ŧ6�
�\�jqu�����#v)�b��.��v�����|�tq2�/��~�C�6�dn�L��t�P��1E0Up�+��D^J�`���W?�ͭ ��t�iĪJ�u�̈��,+lEOH�v�P"W>�q"��A��K؂A'2a�Z�^%�R~��U$�>��)M�q�V�����/�J~����kb����	��
(���eŲ�|�z���7V>����U�SVB����²��r�S��|�`��V�`��8�jq�V��o�k�Tk�	�PU����i#ߎ�}����ST{����a�Rb�h�v`����ik����_>��j�D����8�d�v�،�n9y�i�,q����_������K9�0���f{���sc"�{��	f[Q�M}[i���Tf������_��"���B�L�<)l�*s���nc��zt���[�
��N���NWt�A�m�)_����.���f��zа��j���\���6���Иz㟆����6�!���;�p���aO4���,�л��|bQY���{ۺ�B��	�ϤzVM�
h�0hYĹ��������p퀑n��d��d B��{�
9�v1Uq�̠J��E��M�.&��1�F'*Q~}�{���l����?(`牔'��֘�"8'ڝ�*��Ih}��t��h��^�Ó�z�Zf�J1<��m��(~�R夐���8N���[���e��0��F-��r+y����s��:�va������vT��,��Q\ׅ�] (D�z��,\���c�疪�������2����M�;L�	$mG���Ub��G�u'��B��T��F��;��\_�ֵ�k:���P
y�Q�	�%6�"y�B��L~�u�$~�Y8X�0mI�]b �U��5���yz��#b�v�|��s!%�Ԡ���4�1`|�8�4ΐŚ@���9o����X7q��?T`Jc��{����U��d�U��;3�8�&
��E��-�³�oN�WC��'���a�A�ܤ��w����|��A�T�@�gc�rvT�L�,;*0�ʢ�����yK�����U�8� *d?6c�X����I֔�f�v���M�N��r�*G�h3�#%��S�i鵲"Q��пm�`'W�Ϫ]�R��2�G�������W��"8(G���cY��]�yn�~���~$�#IsH��mo$~��|F��y}C0��W���~�������Z��� *X���h	`Կ�d�7�@��S���_"^>nL*���F�q�pt�Vt�����[��&-��%�T���b�ZZ�P$�����mC=�I���Ь�	#�.��a�(�z^���u5K�5; a9d�3�����t�S��V;8����P8�l��n�(���h�Y3mz�����r�,%�{8���= �8n`[.�T����f��u� $5,.w���o��!Y'D85���x�����b&Fg��2X V1J*�FK�#&��5e�(p^O��>�-�f2Nn|6
��L�1Qj,<k`;�3��iå�Tn���WC�(L(��:C2�����Pp���4�Y�F�<�D�Ky�2ɯ��*$$Hض�1�k���".?�%H���	�a�0S���|-@�Z���������s{�:�8��L��e�G���F,͇Tm�a{��:R�y�nKt� _)h���@��{2�ӵ����U�Q#3!����=���s�eqRV"��L:��� ava�~��g�-�\;j�)�^e������]�%��q�Z�#�Fb2'�\��Y4n�{�?T����8!����K�n���|V�]8�g�m�n��ѥ� �vT�S��C~`=���&�Q Ε�d1X�'L|�4o�O���k��lz��J	_���%=��#��:+��Z0#i�ku�"��'0���q8�M����Vo��:��LՑ�x]����n��b 0�tw�/���Vb�/f6k���Gm	����'�|]zvQR�G�kN���/���XQ����	�)&�kJ��.�����P��@0����=o��8�A��
���W�6�Ԛ��,eL��>4�R��Wa^*�EBR��#s�^�\���r�V�@��+?BP��)�	�c��O�|�*��nӽ�]�N$�5���+[�����O��_��T�\.���4�Du�g��Mll��66�c\tJ@��*�93mn���? �ڎ�8����@��%��B1�������(χ(�֝����@���Y�y�d d�e��Բ�f�]��Ѣ���Hǭ� �
�a���hB�El�Y���:��-��N��BSKNB_������:�<8����C�mN�|���j�<��Y�=+%��A��l[m�L�qݰ�m�]�-���a���ft��u��y�P���a������iw@O�=S�@V&j�5�x�nQ*�&:N�6��뮬�5uVx5��B;���cĹ�g��K��#�����0��h�.uy�)��y���MVb��c�g��5Y$����>!`�p�ݗ��������`N��.V�{�l�6���?�F��;�Y+�u�/�.>~�&2)v?�耓N�5	��	�ɡY�.������Q#�_�����[i!�5y�
�Ӫ�9-ߜ�O
es����U��V]�u�lb�*�\���~qk�6(`�l+Ѿ�:x��Gx��}8�'[�N��IQ"]�x{a ���Ώv���qZ��6�L3�pȧ�������A�-��g�2�Y��D�ō��z�F"��|,� ��DF��q���fQ����Hr��V��4���Me�J@rQ��e�g��(H�tB�W��}�*yNf��RSÌj"��EZk���ǛA���џ��eK��Kv� SJ��L����7��:������˦fx� �����]���$�#��}$���݃�X�zD���氍
7���9_�͆����T�a^�y�����;��9�,�`�����4�k����W�ygo�l;�����^cv���͐Q]^ �p-��ǈ�p�1���l�t����o�>u�� 5j�4��r��Z��%5Xr�MV,����%l}���}��� �|x	w(
�^C��r�x��"�`�.��
`-�b��(*��?pGb���/��8��_�f��_�|�4�RA�$فqZu0��B�-��\؝����"�� � �@�����e���"�j�	�ԧ��V,OrR1&����� ՁVN͌S�b����X��t��(�����R�ذf/�LR�0���S�j����Zg"��3(�^u����z���t�ls��?�|�?�w2�`�����7��2q��%��C`�q=� ��ȳg��
܋9�5�v�T0��;k�#��K�睼gTG${0�o?ЅK�!@e rz%QI<��;d��읹}�������HZiIm��nר�:��S(�~Z�d��)��ᯞ�����)�T�����Ag�=Ҙ��0ڝl�Y�� s�&��: ݚ[�� `3l�iz`G����(O�������Do�_w!������l�3�@��+���g��`f3�ەH�[4�P�q�n�\�z}
䳌w�g��{��Vm���HMRjH���8]���@���5 �'Vl�L�}�<d�����z��'կ��ʩ]�������:�<��H��7��1ï�(AL���FLB1|�AM�~��{�<���|���KB���5Jo��O^���d���������ކ�Q>a�=�Œc�������Nf�ח�C'z|E�T������ �^�z[�]X�Q��@I'��EH9*����8�M��ᕐ��+�^5G�L��^��ĕ��"Y�"}`��f�]��ѐ�]������_��`C�=��7����m��8\�=l�����J��>�� v�p>��ܵ��O�%�1���i�Xf�t����qP�a1�j���S��X�lJV��Lh�SI���ڲ3�����/Ty�r֪�����2�����$3��@W�0^��kpbx�$��q�Q/���;{s&�P�FC2�~��}�H�i�f��e��z��1�S3�-CSJ���tm��Uw���5�[�9w��3K*O�����D�%�{D��jwo'���T��"`E���b��眲1����7y�D*��65O��'7rϨt� ��O��B�Zv�`����j
3B��jc����N�L�K�v��E\6�P2�V�#잾����D��ȶ��Gq�@��D��w���ndl굺`{DL�7�y\'�yǔ�]�y܃�J�!��US�-�t��vI������<���՝
@`�a)[� �ue]��w�2����t�$0ǳ\y�H�B��:��ifkmS=���L����[��m�@!Ԍ�C�C`�Rʈ�q���E�W�{_��KN�K��u{Α��2�E<����װ>N1�����R
�Lt��G�Iƀxs��Rm�_�*�F���z��W�\��fJ��O�$7R���u�7��ф>���*������0�Nj�kS��$���ک�G�M�9tt�7#������gj��}�^�F��y�<��L���uC��!$�8��w$�+���Вx*�[͐N_��c^��#��B��4�TN�W[N_t�Ew����j�[����	�(�/��n��y?Ug~X:��@o]���V�[�K���`�ҋ��A���Oh�7'n�r�-�eE;�@�7��g��OI�s4Tw�ة��d�J���x=�?Qq�Lr��JQP`,��C׃�]�kx4�G�&O�b��s(���#�����f=(oC��p��d��z�bi�a��n�]�2w[S^�� wڿ��F/~h@9y|�� T�0�	�f�MEѭve���0�ƭ���!�=���HEw �;1�3���4$3�x�l� ~�}�F��?�{f3S�|T�M4��A`����b.A�f�%�d�Fl�H��V�J��c3Oyk�G6�Ӹ��TN<� �X�&��?��F2��/�Mq��/��2t(�S?�F�W�a�"%_ky������l#��� )���do���BGQ֧��*uwʨ[�,0ݨ�v�R�V`!�?��B ��c=J�F'GIz��V\iDXf�ৰF��bٻ=�hRg�c�m-4�D�T��M��9�8L�$�T�����7�	k�muU�h;\$J��Y_����d� ���(}��Q_�G�����
R�G�B����e��������vd�?�SQ}����8�z�:_��Q��:WL�� �6VB��{B��3�ӞaͰ6+��Z���$�@��#�tp��`���c��ILD+*��Zt-�HT�����ӏ�[��ζ7
�V��%�,3D����X�ܶ�/IR�r����=}Ugd���c֗Z��0b����-_K��o�jeOdD6Q{$I�A!Ekޜ]����%W ��^��2�[9*	@�l$����\ ������_N�V�J�d�F7�:Z����ʠ;S����M��~�` �m0�I�a([{�c:�����r;�c=��[�D��'a�ku��R��0^�9%��f�'����R)㏎���v�
�����ǁJ�gL�@�`v��u�Q�t6��=��.�1U]���\ߋ;I�� n쥤� ��/ �ܸ��J�����g�!-�b����S�w�D/
f�_i�b�jf���h��úO�&�.��K���E���k�#!��u!����8��k�v��o.<�@��D[�m�P�{��)�[�tLS��x�C,��*�h@��P��_6��d��Q�Y�J#<b��d���kL0G:f�T�Vm���c%;��R�%W�o��~�<�Bm�4J�3x������v��'x�/ձ/�?�*��:W��9�TY(�f;���#�^=Z���C�i|�v�S�m���'cWJ��&0$"�}3�����t�z�wG�lAX�Ó�9���gX�)G�d-n=�I����M�!`W��n�)�)]�Lz�b{x�-+%;sZ��߽$���k���_|�E��JGp�
��t6o
��Q��׌a[7�-m@=����ݽ�R�Z�o�f��GS������VVן�pWZ|�v�����z-� ��׫UR�p���aQ{x��)�1W��.D�Fj��]�������Bi�.����x2k(7a>�����)���3��mg[��Ǎl';�˗_n~�3ez|���GBD�{���\A/?�q�O���wHG����r7��jU9�������{���|w�>7�d��mU;����Zv�b��q�BO���4��o2��l�f{(�f=��'8 Vۡ��S�<P
��J���g����;��l|ӣ��:	��/U�.^��0�n,����D�UB��|e����r��zB3*�����W����v�O�[�d��^֮���WJ����_�+�;��R.��oץƳ�Tq }J\���J`�-�h)��Sn6��oBz����V��Ƿn��!As�o�y�s�_���W�q�UAeN��jN��F_�H|����/d��̬�AP��ewJAKܾ4�]���q��`����W�0��*��"I�A ����]����^%�6��뇑���Be�w�Á� ژ��e�E'����G%	m|
�G���iD&���[X�]����n�O�ɫ�������`O��4�>�-md�ؾ�ng���#�ΏMI[�پV�O����D��>�	����.��d�_�Y�xp���L�;[C���"D�]�H-����}���0�;�����f�7�02wg��թ4(��85,��Ρ����6W+0�n�C�v�p���@�=�5�J� =��8˿��S��}�w�q��wdzC\#�ͽD����A�S�ES'��@ǛL�����6y�SlA7-�/�3��-*|�71�xJ��lB��S=Juֈ�A��`��|�8z�aP0���\u!t��L�ڻ�4��<��h�;��K_\G�e�(���5��x�3~"����*���a<�N),�ǰQ�>��_px\����xa���E���O�h�R�aS�bw0�W5�	}�2�<O��p�\g��RX
y�w��Y_H��RM�$Vm��V�ю��� ����W9!���6P�{G}aç�ʻ�M���yX� �]��&=�g_�K�`F��＿E��-����^���d4�/z���L0��C�ى&�]�4r�G7vVEq�5e�5�,͖15����!���Q�h�i��4Aau_������ bZQ�b�ݓ����?.ܞϫO�H�V��ϙH}��b4Խ�2���`[�LSXd5����UsV3�w@�,�7��iE��X:�ڶs��Z�}c��v��I�E���	�J�b��o�C�s
��;�0�����[�����~i��P��<+��~���0��CGm�Y��OL[�4�5�]��lkQ�%9�%�[&D;Vv�\����IO�~*��ٲnê꿣��I�����jXVI������+��Þ���M��w�%����q��(��ZDNka���1�0GjX�q��ϊ5s��l4I�A����N�Q1��L�ctJ�h�:���&y?��B݇�e���ܨq��Q�!b %���g�N 
3�I#@.��O�tw/iPj��(��.E�[On�	TI-՗��r@���K�޷�L�����^Ҋ�n���kC#mI��Pa��K=�k,�$���C=o������]!�����p�g��7��Ġv���i;�U��T����1O3��� ��U9ڞ� ��!^v���I�\4�7Z�� �Z�[ �7�W�J�.�`�z�Z�G�\�~x��͢^Yʁgk��irsT�4Ds(���Y$\`UYŰ��cM�y[H����f�5F��ė�v'��U���k�m��|ˉ�0��T���0(����'-]b�rb�*����
����}��6F[� .��*OsB�{rev0,�!�җ�r��Q��A8IT�����Tz�k�4�D�pD�<�I�+v3>��3��TA��V���z�M}c�3�Cê���) KG���C��Y�^牸�����es$sM-�9v���[���6�:��*7W4�P��F��Zif �r��8&��5�L8�4�h��4e�5Z�$;�!@�;�����X�wA�ߥ����8O�iJ.��h��"�7��	�z~p�B�L���m�v��)
 �"��9�A�З�����^j0k�$Aqw�O�H��	���ϸ�f��㒳�m�L�t�(c����~��dXU�-1��*#&�SN
S�� -ʤ����:B�}�#Io���T3K�E��-�qAT#|@���*53��|sq�`��)N	�,y)e�f���9��W�E��36�==.IDh�ն�7����ߨ6��^�9<w����>�y	�8������!ڪ�Lz«@X`��I{���J)-6v�?�QH����"9K����������`g�s1�,�$�]�>�eG��,ff��%t��P	�;����D#��	�ϛ����������w4ݘ��ᛶ�0NfOզ�4C�K��E�$^�R^�À���"�D�NH������yg㝇�nu.��Os?e�o/�ŵ����z�ޝA�����i���_w��fm%Y��9�:|��e����l&g�	���V�r�B(�Y	I���	�yZSb�K�$�!w��ªP�Z3�&���$�!�4��� 㸍���i�;ܤ3;��V��$J&�}�3g�H#�0ă�^zvR�J�v��5w������"v��8��l�txp9�A�wq���=���jH�Ht�v�&�Ȑap:	`�@�V���_�a��ݩQ.�ߛ�]Ju�p�f#n�]ބc�a.S�ܢ`7]Iٛ�	h)�
Û1��y��ͺ䎝R{�I�q��<�*�b�i��� !!"��rx��L��7�il0I���"4}�b4�k������J>���i�)�-�>� �+������/��(�,�d0�����#8��d�;읜v F�k1�'�R�'Zy�`g���`���0�]�ըԻR�z#�!,@��-��k���	��iE��ȝ�8���kA��j<&�1 �󜄸���2-T.EO:�2����ۀ�J1|�V�������fZ�SS�/�W�����\�<�X��?�}��KmOr
Xв�_a�&5b{,=�6�9V*]1�y���õ��걶"�j<�2$R����8YR���+- ,㒩mbBRe�ލs�Oؽ� �Rk���d!�:��J�{���'��<~f�Oz[�����	ڽ��_�r��Ψ����B|C͚���}\B�'h�h��9y2�'��B:z�͔虖��fu��>NTw�-�*��6.���b���\Y�fn$'�e����{�=�&,k�w�9q 2��ڂ��o:��/�my}%.����Kŵ��՝��4�� �8,cB['������Dg��.�G wp�ޭZQ_�m������.�z��]�K�"6����ͦA��6I,�N��GI��M;>�[���6����l⹮�p����_��g��R���#V5���]��v�s���&�4�� !p7�M�Li�Ωz�rH-���6�@J����J�P���Th�H���~��<�X��>й�ʜ���pq}�ȯ+N�.zX��*�J�Z��P�`Pfgq�0����ؓ��݋5O�k�-�N7���n 2�h�٩�
����=]�0�}r�"C�l\�B�l����!,I�)�k`�`�h�H��i����A�Uؒ��o���� K-yo��s=X�kV�o.���g�J����,��4�&�-[�л+׫Bh(�Z��{�sLԬ-�;x8��������r6�8�ل�ha9�(iJ�e�>��_j�.�x�C F�t�:��+'z�����|,�n�M�7$ύ�XI��g�0�Gɻ�-�w+Ył��%����O�ֻRB������xG����n�,�(�s�Gr���I����q���P�(������`%2��_�`v�� SP&�qdtsd��/�٘=jZg\�ޠx�և{4�O��2Z|T5�����B߇����)5�^T_��i����Y�4 KX�姎��y �z�S��>�?@�~��dN{d*.��̪��m�ep��a	9t�szn|T�
�-���Bނ��T�akXJ=r)K2��ݤ5�c�4���us��Oꡢ��/J��~L��M����%w˶�1�~���_�M"��[�z��Z�u'��J��ռ/�D/?����|�\y�x�ca�
����M���2��h����\}Ҝd65�2��b��(�gw�3L���W�;�K�����	��2�M�tQ�yɠL�D���@�;B���u�TE(�7:�x��(HKE������%�Kq��(�	3}+<CLɄVņAJ��9�mQ� �&Xϥ:�h���e����ҌN��1U����.H�H���F1�������c��3kRxi]f������Rea*<�}E���Ch2��nd�r:�n�F=���8��_�c�_Ӆ��'�Zrsc+F]���JYq<c1J�ڗ�LQ�嶟�Z�������zσ:�[�v�*�gŸCR����[d�ف��&]?~�EZ�����7Ɏ� F���X |[6MNqƉ�q�M�SAL9GX��ʟ��C�!yMmkz	Hc��ڪ�n�A���'�zD�� J~D��\�辎0PhU��E�A�9��I��COc�QyQj;����N�v�7�1�C���-����j[��g����,�9�Q�`�䢢\�+~�n��9�4S4D�p�����ތi�MT���MQ�ܦ�g��y�x%�?����r�_@��X���NeO��޸���p#���)LaC�-�M��B\%H�G�n�`l�QX�XԸk&<'�茔�U�4tl��I-N%a{�mV�/���"3ǚ�&{ؽ�+��h��/x�_j�"��G-���.��'bK���7���q7bFZ�52�<ǗqV�9��E8��Z�?D���
 [E��py���z����v��H����ي�Uc�H�Ҿw�T��|��#�Q��T۟Qb������0���d	Nk�SdLO߹퓂Cw:�K�H�GF J�BrG�G�x�o�9�VP����Bҩ�+MLe"�?�~"3������D�W�iP���/4�������,YR�]���w�D��F�H	�E���-`�׹Z,o��d*:� �PH�#z�0�����kK��	96�����
T֡&i|���C^^��y���Y8܍{I���{������(��zi�L��.$����͚�v'�-H�\�Lfw���N�9�L>3�,�vj�i��8q����ˌ��ԇ��"F�я�l�Mv=*%a"v^��S�{��2�R��fR��,�:�,}�a`����]-���l,S�:����j]�M�w��t�UM8�|��42[IyY��_�yE���۱;ӹ��A�!��A��JvsT�$j� 	�Y�/�<a��tK�ϓ�j��<�l�B�I�z߉�R��cx����Bn0Cݕ	�h�O�)�8:b�U�+$'?֧��k4"�-S�:j��I�
D�c�\��~�y.�Ը�1�S�@�����c�°�w2[pN"�)�HR[n�Llv3\_�X�g���_��d]������X��/5���~YRӡ�%���?������l���Xc�E��.���o䯣1�!=��
�s��QŪ¹V��G0ۿd�ԬnF��Ӏ@K�0���d��D���?�՝�uf�.}"�)�z)�O�%R/G~�Τ�_�|�W	�w�d�z�m��-A�,8L�-v�2�;��*�)�\9��66�,�~IJFi=��ǅ�YF!�Ŧ�D�AH�1ʻCӉ��(sz]�0��),;�x�]g�c/An9b/���kO�C����x8�g��H���R@���e���G^���U�7
��C�'i�"j�=j^���+�%��E ��2I7�H/��)ַpy� ����p���R���z��,/�Kw4xu�g=�a��Dx-��Y�S���_ýDB��sԭ�5�黬�7b������T��^χ]fB2���'撍�����10���@���|�o����Y�ĬӋ�Vv��m��9���n*�ɥ?V�4��Nl����ppf�u�ax0C�"ʴ�0;�N��~�Z'�p�{����?�d�f�x5D[��S��`���^��FU��[�ٸt��h� I&	b@�ܵ���O��y6�)�Yf��˜ �V�D4��ˌ�4��ͷ��k�x��src������4�k�,�蕹�oW|����+�b����u{׿r�%x��v_{���Wƽxu]�`�F��h�3>�9���a����V�go������ 	��P�P��#o�(�fW}���c�IM>��ބ�Y����y��p�EB���r�=�'��ǵ3��`~>!�mײEh�D��"���� 8�_ڏ���=ɧ�^�c�Y�Ǔ��.VS)Z���p�)7��]WXH���`qFO�:�y���'�E�q:����SpX�m�bx�L
��J�2P]�@�"�t4�a3�?��֓�h���#?�EQ�D�������:8�}O]��3r!]�W���&�υ�鋑$ƫr�z@6�vW�������d(���)��s���B]#�1�$�{������An7��=w� ��"�ZR�^��k�Пx�Q<lwae�_t%���}J���[4���o�U"0V����9}�������#�?���S�s���$i��O����Y��;��%o.�;�i�x�ɕ�/TW!�F�դ�{���ԝ���]���[�^!8�[w����v]���	�[�:��P�NC�V S8&���kG��4�'�,��v����9��9���uk9P8'PL���<`%�(�DG�9�N�j79&`XE��.At�j6��l-�nc�2�/b��l\Q��0��p��$g��:���rv�a�(���5��|��kn[�����JCm3{��������θ��U&Ѳ	
��mg���q����媜��)��n���z����;���ȃG��v�5%��mt�G��3N���@
����J�T�Il+A��x(?��?+S%R ^�����߅���K�MPw� 1i���l[p� �Bi�cjy($��q�5C�;��ޙ�&a+��O&*E>����������x<�|��F��R����T=H�*~ِ�a*0���@�R��� ��r�]�=L:��")�Js��֨��{X�&�<J�bVʥqem��ڞ�g���_-,'���/͟�[��ICPK���p4ZԪx�<.���z�ٴ�p����ȸnwbj܄̋�b��ϰ@I�����SVT�a�qss�Y����/r]�dM�:vy�;��G2Ӫn0���`�,a��6�#�VG-u	��࢈y�Zi�f��tZM���QqΜ���m1H�8w8�oî*�E>��sXJB�ݲ�kU�2�h��m�C���Un���I�.s�45��/�1/��<�Al�2Y�0�н�I�5Q�z����������"~c�]BH�Aj��߹lխ���'c��:kp����������vs���O��l9��fӓX�/ݍ�gm��W}`4,�e�������ʇ��I�'��wԝ�d��S?��I��c���PB��!���<~�o�^�6$V���Nh�_p�-Sx�l�R���G7o�{��|$[b}]1��Z��\��1V���߅XZ���T��<��D�|���w<�4������Jϊ!�i��_	���ޥ����%����7�2a����K�B�̀��XZqO�@y~o��et�l��H(�Y���kw�j���Iʘ��F�)Y��p]��tw�"C?��l�{�ګa��Ka`⒣I���o�7�j�C&%�A��A�`C	��#��q�
&ջ7#��`[g�H�����<�n��?�z��m��aK���a��3��2D{��������x���j^q�ΈT.W}���r�׶�0v�5�u��u~������� ���?r�ݎ�ҏ��|�����0��\&��LuJǴЈ���c�H_}��=��` �1�S$�[��,���'lv�8��`���"�g�e���4"P�W��'$��§mM�*Nύ��O0�V|�jX�dK��~���į�'%�4�^B�Y�sH�1��4��U��5"p��=m��C>_)��J���������B��=Wz��̔V�!�WE�g!�fYŰxޱ�?��z�2���p4;��s�}� 	=�I��A�7���ct�bSŠ�y.�V<QbL#	-D�+xRJ�w
K)H=q��_��:B�׷2��L��(�^Rz�W��*X���s
1w��g\�W�Z���4r�W�n��-=ݍdz;����.D�O�k��sQ(���MQ�]�F�&��!�r;�x����F���̩\��<D��-:L%	lB8]�o�j��<�bbr��$x��A�?��!��|�߅�8�ӷO�
�R�����Y�k�Y���Rl4{p�C������P�"�I�h72�nz���Z���_�L
g��i�NJ#`���	�����-���<�'5��y@S�����R�jԓ~Jԋ2�'��O\��O��m1=;���b7Jۇ�w��NpZ�N����n&q��s���3���wu$��������k
H0T%�#"g�����ߧ�gG�myNb��V�4��UM�j�N����^�ʴI�M���'�0�r#@� �TB+\R	gY
Ϟ8�^��ɦ��Mz�&���^��vϕ�R�o�TF��f�H��C��r[�9���˪��-�� ���E[��fo���;�)h���D�.��6h�x�]�`	Ks�_��#%nҖU&e`L�歡��z5�/m�5�Am��R��	C3=ۉ����n����jG帋�z�a��~���¶1B%��D��,��hIؿ
���T᜽%��y�**i`Ph��F",�£���e�����<�Ƈ��?��� j6���m��l���H�ʊ�����(��W���D���������'�_�2;�,��dJ�	>)����J�h3��S�ֵz#��"�dN���J�|y��4&�5r�N���+z�iC@����p�R�N;�t��M�U��$���c����n�Hu^��j��[^>.��a���'���o��W��Rf���3�j5���.2�M�9����ۿ���7B���3��H�q��q�yI���ֻ�Y��N0<�4�d�R�G�j� �o��7����=K~��t� L���C�-	r&�s�FY�ί�ױZmb�8Y&I4�D�o��n�W�s&=����ͣ�{�x�ݭ���?_�X�eA��Q�?1l����A��
��B��%=�k�M�\�E�z����g�y�t�\�X�J��a��Vg��N&>�e/��	�jС���'�M��O- Kȧ�5|%>�&Lۢ��gPrz���x1�3?{���68�#y$=y!cr��N�U5kAh3�gfk$
�Ǔ�S�wm7�eE"����
��3ku�d�-л.�~a�˛�������+]��b�e�r���mDL�W4B��΀�Y���j+�Z��L��k�<B�B���w��/��p��@�9a������lO'�KJa�=��r��1�|��x��.��a������B�k���p�;:�X�/Pc�U��<'NT+��Jmp� �/U��#��q
���Іk�K���?����B�)��� �����Q
j&�Ш�d.���[�, X�Ⱥ#��P4N���Y\��� l� ������P3H���@!�߳'�Q��̟��Ɓ��=�/�p�H�T�%�����Q�������7���M9�)�(v����Ņ#�'�v�sz��;kg�'PJ}򠬰��͊�*����=��|PY<Ɯ�_c��{�ĵ&�_u@�r�3������+|�qm�;3�S�Z���9�Y�6��&M��BiMO�Z<�$3�����i�|����2�NU!4b����/�b��*Z��b��E�#a\:� *��rX'ge�Cp��b�Y�(9u����H�ݩ����8&Ir�V\�x6�G'���G���'f��e��9v8(58���G��<�ٜ�|����B�~ǜv��3��$�E
s��$R]�$rk7�D�tJ=���V�a�!����+�;�k���^p��<�a���5�Q��aԛ�G3?@^�����4��v�`'D�N	;%5~��,G��,^��n(M�:p��7���ujn����������pM&�����ޅ�-�������]J Ao<��vp�1�$�_�%L�~\�&�LJ��N�L�٧�Q?�2�CP;���)��=�%+�UM$�D��>�Ց�wX����!�u�er���0�Qib�]�Z�&��K�;X ��B
Fx\A�XS�.邊}D�Z����bN�W�z�6/ �����q���d�{���s-�[���i��M��R�cf��o���*�(�k}�CyN���[�=�p$�@��fo�Ҫ�,}^�7�G��WRLuQ��)ƬQ�d�N<�tI������h$e|�q��FH�T�8�
؄@�{q�d�vb�F���(�����Dx�7�[����R��V�/�Wy:N���PLrB��ç]��3��ߢ	c�'<�͡�U����=b{��F�l��[i<��H<���qZO�(�Hύ:UK
�.��ܮO���Ăx��6M��]�+j�5�Ȏd.��w�<*��u-�F# ,|�tE8i�P�-����5k����D5!S���h�M�K�L�W@o����	n����S�u%|V�Y����̚L��jY`�?"x����4�E��|���5;7�'����l/\���� [T�B��T2��$M��5�����q��1<̙ ���L�?.5\��{�y�Mnm_�ˇ*c�VM���=K}�{�d����m����]�K�����˷N�(�_������IIDpe�c�ުٮ��*�7�Q��2�U���h�zmz`�͵p���ɍe��I�!�lG���}7L0�~b�,�Χ�&���	��R�\�'��.��Dۺ%ZJ`o@�JZ�=Gؙ����k�i�	�:�]�Q�uU=L�,���E�_��K,�Mw�=�'V�����M¦	f����7�����f��I$���(nėpu�"<�������$��-K��#�Aξ����	)|���k���@� O�������Q�BH��f�bHn�ڞC���#`}�~�IN�f��*�=��Hy��c:�=�7���ފn뀽J
�~!� ��ĩ7/,A��9���C�F`.>� ����"?�z.�!����x]������*�YHSں�՗�Ăz����,=:I�rN�懼{�9m�4,��۷�gR�y��Ib�d�����QV��$!���5\v�kcs��.��l���OЂ�#��m��6B,{Π^��-������N0+�4���"����6�$���4�4�������o)	H���\q�i��~r?�\��R����6�Ny� P�w���2"{�s�X�c��P+�I���� �3��@��l�d�^��#�3w�#�[�V+�Iv|�Iy%*�ɗUH�[v��y?Q���S�	4 ��K����<�`�BXt�����MI�� ��]�G�D�|�3?�[_W���t�-<:ꛖwq��u�x�q��!�	H`����{C+��:���a�yFn�zQ@��>dh�z��R��w_!f�xM�ЬL�[�ٯ���jPş�Mt@�&�hZ��m.��NS� ��ُy�A���#���:��@t�����j�虇��u��c�^6��J	W}�J-�-GcWS�Ƈ��Kk� �r/���"N?�PL�M��k�1��KLn��@�Ug�ϱ��߀��I\�v�KJD�Fa�qu58Gf���} f�ί_�VT	�-(U��p"Bj \� ���Y�@����j)͋ �zS�p�q�n��a�$%�ٌ��G����8+P��p��ʶ��K5O��%�D�/�S� l!���.����R�IST���S�l�y��<�|H(�P�5+-탨��<�;�sX��u�2z#l������^�3%m�\Iš|�	����J��
���/���}OS��XdSkTps���+2��[�SU������F�i�*���0�>o'V��7�+��O�Eu؏s+��6|��t���8��U����y��� ��S�?|��bd6��9
��_\L��ʂ'.=�"����xv��Z��Z�����w�*���i7C��0��"��@O�Y�}y������R��{�8�۾ ���@hv�D�x��Zd���v��8M�	89�-A~����?H�k�s��=y�mY������)$��
&#14hXRg��q�ٔ��)[��M�D�,�|H|����L�����=0#W���������f�A���\�n�N��e|��WbEuv��<��S���V@��`:c�Ě;מ�py��#n���c��îJF7���gr����?�?���5j(n�����;:���F�]�.��;�!�˓$l����E�ǀA�S8�5<���w(O�ci-�b%��'/�o��+�+а�=ɞ��"�R�X� ��d�e����L������%h���M�WT�1��	d���؉r��f�q��'�m�ר@۫����K8�4��¼�y�P�Z���)�J�Yn�q���P����vō�!��1�jr���Q�9r�q�gJl��c҅�ew*�Q؈^S4�_������hD�h5�Nf���x�94~Ay^� ^�������qj���`�J*]�PA{cY���YPH[PU $`?�(��N��"îؓ���H��jZN�':�G��Wݮ��h;�#�%	3�8����M6 haA��A*�u��w�g�r������[�����t���D�������gsKӢ�H�;�-X�C�Qu�}b��%�q!�	(�AI�%�$�����p`�0�Vg'�쯶]W��+r�7��QL�J�� �3���@E�q��?�3M���4f�US�dM(
�f���s������VZ���^6�a�L�U$�q��cp�@NL�
�V] m?aj6yZ*���Q�y'Q�l�e������Y��4㜃rӁz���G4M�	Sr�հ�j�WyL<1���:�2�e��&y�:�ǯ��u�O��hN�p��KY���>����~:��w�Q��ʱU�6�J.^T�ʶ�;k��(q��O��p����R�#�&��v����m!��l�[壀D�Ll�s���ۛ�<����eP�)xk�ɀ^7���+-�V�ғ�b�]�����ۻ!�<�i�K��^��^n����7 �2ujC�8m�H�}�	�ק���PH|�ٖ����(kZ(+5�g2�,���Z��L�!$�<�Aݣ�:Q��+Al�݃0D�5j��T�H+�$�_P=�� @h;�Y���ȭ�x�O���F`�j�b�ʜ�w��`��|�[�UP���Jq�> �)��������-��H櫯�]s�?$f�p�z��񮢳S��Sc�w1��D~�ڕ�����m*Q�1-�;��\V^����0"b��xP��n3� G�y8=mL������5��~�ԓ�܎���-J`�s�ߴ����TT�7����<حO�DыȲ
�hfY���t?�Z0^6���n�zb���*��D�zEA��! cp�iG�ڰ�%��~i���'xd(`�K.�g���}P����k3�^&sm�r+�J�ƵҶN3Y����@mϝ�z!xf �Q��@mt���*�� L�ȿ�ж���~MT�c�P���o���Q�
��>�e0�=���aa*s�BRG;�˓:}y�K��çT���(a�_��0���>��4
.�k.�7��멛��F��y��No��=�)y��J���l����Ot�?������z�.9���= ���^��2��8��]P�]ac�dC���a�o �b	��ծ�oӉ�b[��c���9	��`�`ݝ}|��[�K�ŜT�݊;;.��=l~�sJG��"@j����8;���$nǘ��G�3��e�-C��|F�}������o���ϒ��j�8p�TQ2,�D
���g)*��0��<��˽>F�$!�@��J��Vem߁�<~|^AHX��%�K���r$����Z�V����k=U�r�&�
��Zm)Φ�[��̔��ʪ.���a��L�L��6�wϕe6)`�����0�|0=�.>� t�C&�,��ag�y��@�u����o��t�q&��M��y���c�c�<�YK(��!Q�7`���Y���VMd��;O�Ʈ+�b�Q�LU�ȉ�d)���S�I�� Cȿ��s��δ��(���?�M��4�o)�3�%s����1��WcL奎-ݟK(���P9Y�d���v69݊X�~}&�[8��%�c^���"��p�������h@�F�h�f�R� ����8ky䜗5Q t���C-�zj��l���?s�g��hŔyL��7�ͤu7�ʧz�!�9HӤ]Ezj��b��{���ۜ9FSw���Y�M�,��TM�pQ�ztc��=�/�,J��������+̃\�T��˰�_(w6���3�w�b$�o'I���R�=p���:Ԏ��<n!�Q���dPT���i9��yVqtS� l*#5���;&yU~]�����ql=+��Ԥ[J#��4ր�煰���sH �����=i���+q����������O��KmT����(C���rN;V�e���̰��ہX��{0�@6���>���f�D#�քjO�:J՗f+|���$%Q�$�i?DŚd��������M��?S�#ȡ�k��s^<l���+�x��k��ܻ��'���1�:���0���xA%@���|�HB�ӛ�U������Q����4��S��.��X�Ĵ7�ĝ5�ݦ>d$m�T{��0���^�����剘�Yk�}j}f�.���pe�V������iW�lZ�B���u>�$�ڠK��5�� Gח�}���%�SE^��uR"��H-_��&���,��8i��j�4�V��{BCB;o������k����� -j
FT�9rj���v������DTT*8ZP��m�Ti���G�!sH��vg���~�0*#S����C��_XJr½ �B���y�zӳ #,�D4�I���K� �C䗛��vj��N�C	o#P��x&�S�ַ8�ht(��
ũ�+�o� ^_	�5q�<��6��S��,D|�l�
��n��`e�x����퉳>���-qz�H����ы���C��E���>��# �L��FF?߹�6A:i�Pr�V`^��Li�"e[ƃl
�e:��Cb1De�rK�G+4ܵ�܊\�M��x��~��%^��$59�����N���EZN�<zS�L�̦e���v�X�k%�rN2W�	�f��K��k�55[b
���7�O�(�ϳ�V(w|���~z�|�c5�5ϴ3P\��"\��]�NY�=�}l�|a8sj�%*��;��ۜ�j�y�3I�NO���<��AG���. �Q�T�a[uE"`�Q���ŋ*��_�ic��w��uڻ�ǃ"C�~�=C�9޵�fT^��_l4�{���n���R޶�̹����}�fS}����!my4��h�+�ڠ���Ȳ�S��L��.���M�la�Z}e.~��P��D�W(�|6-zfk��&���1B�l^�y/6qC>M��(p����3�jz5�B\0_�(�8�ˮ#������>XC"�n�Ĭ��Mw9���y�F'����k@��zs�[�t\�6K����Ԙ7j��]�X�����F��W����Y���[&`xgQ�>�Žz#~�uf���3�"�%��2�;��c^��W]��պ�%>����i͌�e�@;o�`��3�1X��[SBl"�3���Mv�3@��}�9�5P
x�YE�T�c�f�s�:�$&p���Sٙ���|!=��l���P��ϙFI�+ "�u�*+����{��ɛ�׀n��ܪ�1߶����`w����OF?�a���ǻH+=柛�?� �2s�M���E��1ި���^.?���5~�e,�Qo4��N����Gb�i�hNN���4����A�c�9�#��A~I�1���JN�2��9�o0��q�ØU�Ղ�J#�]�L�Dޠ�i��1�኶�b��*�]��	_��⩓�Q�w����5�pG�lD�����D4��"tj�l��ޖ��C�[1��ѶF�[v���2�z;8[��c�Z�92���J�#v��Q`�ܕR��7CnaZڿ��ʺf�]����c�d*o��xP�P6�c�(HT/��V�a��d�\�W_O�����qX#Gԭ���p�J�4�nʜbx����G2Ƒʃ������g6��$�]$�� ��\ ������$�1�ۼg��;h�V�Qn	0��.���V��%D��E�z|k�����|��,L�#��؞�;����9��o'pP���Z(9xIM��|O}G[�	��jYh����N�w6ّ��Wƨmc?�n�UaM�Z^%-��tG/>*��,�������f�P��(�h�si�����j��Xߏ�+���@v�	�+�ݑ�)Z�VaC�C�N�<]O�i:���� ҭy�E�[�.;.Hw�[�gSG@!y����(�q/�x���ۢ���p=tVf	�sھDﲬ>
���7���O�C)��������*r�Q`c�"�8j�-�0�O���ȿ��C�ȁ��5@���q��6)p�{+�=�L�U��K�[�	tImƸ�w>E�8i��Z���b��i�@;>��/1����z��]Z�k���N�D}Y�Iv׊e0[H��r{/�ƜF�� ��6��33��J��T+�'�R�u�L���D.����I�P�8��J��:B����/�J�������.ŧ<�a����,��!ד��Q��8+6,H����W�+�$w��E��s��O:�v����"�&��ʓ�t�腽����J�n�$��S cG��T����p}-_�($Vk�v����}���Uac(�P<�f�Y��[���@I	y��`���Aޠф�?�C]߸�v�	L l��5;ȱ%�Ʈ3[���V��-&Gz�Vʹ,��F�t�uկ��#.�O�%ܧ�]뤓��*�	'�ۺ7dW�{����&�۹_�'nУL���_w��
�$��y���@ý��k�(	ǹ�y[z������哖� GIK۳���9ͬ~��]e(�1�$��λ=ĳ� ��v�*JFذ����00������	*ć=wõ%_�lDz�GX=׾Ca0��{��N���n>�Z��{�u�i�� �ׁ=MҊJ�#j� 
����� ��d���&�0��r�g�U��y?(�鐮��<���l0(I3�j���������0��]���D�_WHKF�|��z� ӂ^�s�����`��o
�P#�J�LĈ=�_f`��������{-o�Ux��@�"���VCE$��\u�#���8�p�](���@ίA���L[��A��pCɎ��Z/(�\߮�����m�)�a��b�ꛐ��3�IZ�y�,Tj�άo�ޫ����}������C�I_Y���}l��� ��A�Db\����T��~�tlp
��>_]H�|�.1�X6�12�Wǹ8}����hs�A�m+�?\z��s8�����c�@$"��k��24�+�7�P��l���%)>���e[}�c%��jw�Z򑌔�z��H�);�K$� �l�=f-�N�6� �������!�N9�$�����i��`!��]�Y5z����%�l���jI�v��7���tH���  A�^9����K�V���7�^[�ya��Ʉ��B�����ؽ~��:���i�oUMZY��[���hS���D$���&��J|OY��Iksu�y�^U[8�5��z6CeW�d��uV��;Fx�/T4v3@��/&5�K�s3��I��@4_�vm��RJ޵.���p>�-��ְ��K�N���xL�/�t�ɏ�hM
�������e�#�V���B��aGd�a�`�ld�~^�Ö(QWKG<��sj� .���}��7%���"8�hJ�4�G��K/���zv曓ʽ�4�՜��yZ�b����-�[���[��������\��P���G*ڼt���j쀙�1�Y��駃��^3�I�_\&U��Z�Rh7�����8���=s�,,�[ �B�e	�.&�
�{nL�Jis�l���Y��Hڸ��r<8�h�~�6
��h��X��G�Ӏl�Y�i���+9��Z4�!r�տL����m�^c��ʠ}���
�~`?YO��|:���7� $Ѓ�������I���j;�0�������c�ڈ����L�ٝpl��NXO�j�������Q=����su�U���a�;dT��O�ӬEҎ!�K(V�C�nӻ�۵о?N�oBA��%�x��y�[�g�t�m)���ɾ���[���i��y�2�]��Ml��ō\��d���M��s��_��;R�6p?��}����S��.4�;�8_@!z9�g��B���kYu��C��<���]��U����&�~WG>n&�-��dp �ߡ�s�e�YF�a#D,�mrg艒}D�G`�/_9����L��1�2� �o����>I~(䬢��S?�� ��@7u��)8�����n䭾�ְ��4t�8�N�O#�� qa�rU��=�§��&��v�7z��������]�����Q��\W(��V��_Izt76)5RYbC�|�(��<��fE7 �F�o?v���%����6	�E.�P	��ܒ0.3�K�4���Ӌ]�a>Bo3�d
J�����HG�AN�m����;\h�a�J��+�q9\�����B[�_�B����l|yu�M��T��:@���7����Qu �	S�qe������	A��r}��'nRmcn���8�ؚ)�!����u)H��*���ٱr�2��4O��(�2�'����P^�7��y 2Ƀ\��D��������q�����igu���r^�h�"���jdz1�^����ey)�K�vZ��+aI�tԟӇ���y~�:7���'M�H��@�|w���:�� �y��ۆ�>�H2+E�b�-�s��&��젊�i|�z^*�u��������l�0 ���$��7W��YGk[MPV�c��Ӓ�`�����������З._k��3����)�Ҵ�ϋ5[_�� W�ʘ�T��J4�ГNN{���%�/�]"삽s�����a�DO�@ ����|+��)ͤ���p7<;ɩ��� ތV�ǣmLԉ4�=_��L��80;}�-�x��y�)V3�pR�}eb���dn��g�b��C�L �1D��YP?�W�씿�1ڜk&c�GG{������Nm�g�a��wc����$�(�Cރk�3z�^�%�Е�<Ն� �-8�h� ��������k�(��^����8�G#&x��dQ�B e�W��7`������PY-��v�	�nT��.�<�\H��|G�N�O��P�N��Dt�i�])b��eq������ C�I	���5�q�d�U�O$[d;���go�*1���q�p��n;�J�Qԭ��d�?�v`�����L����P�l�0?�T՗9��;MB��n�24m����!�#"�EK1���$Na���8c�r�t����d�&$:��7�a��\1p�5�l��k6l���p�AP*֍�W6�aS�F�N��jB*[�4|J�A���N͜C/&��#OçpoYdl����Ԓ 3�{���}RwYi��}{k�t�n5&��'�B �.goz֞��u�E	����2F�:-���]I^��{�ap)�y��]Ż����9��� �Ci5�1u�%��~CP�3f��܁�s�0�@3�j��yݙ+ax�	s>_�!Y����˂^X�µX�
쯁�L�\�$ITvB�W�'F1=��	�$lC8ɱ���%��Ӛ*�B픬�n5���`�l]�\i&�7y������/�ǻL��k*�c��`�	DNu-���'�~d��c��gt���w��J<��Uk ����Mռ�I0d5��A)�s�[]�ˉs#�[!��pm��6�.��)6=��^�i1��z8O���HIܐ%E2ŜU<�ʷ*u�S����%m�E[T��\����KP����79o�#b��mx�6�̛�E�<e>��H�a��-��=�fF�q,dd]kw����l�gZCL�d���-�Y�!|��	#F	��CĖ)UX�V��]�ө-Z�7��sZ�E���}U��<Zo�9|S�?�T2�$��v&�mf����H���1s�H H�q��9#ѿ��������׊m��j��	���#�e$q,�c?��	2ܐ[o$t�z���C��quؐ��%py:�_���8sH��wm�H�J�3�P�#��6���p�{�x��
�:|����5�,�� o��<�,�tޖ�������7�Nˉj>��?�QQ����J϶]�g�&�Bf�#�r5]P���y�)�s���iۛ8��E)t�.�sڥ���X1�M)���x~�a��݋'�$8�r���:�o1#�3]۰.�������4�k�#�J{(�b;�}*�ܻ�6I���YA��~���>������]#.X�5�ld��d�p�n� |<r��/P��2hw�&��̣�F>ݝ(!�Z:�1Θv�`�]:SV�$�iL�������t�7C����nV
��֚)$�S9e��Q5W����� �(8=۟��dXx��|;y#)E�դt�!�b�ϭ�=�R9��b唱�Mp3�<?��Z�ʣ$MpH�6A\ס8Dj��<A�=(=*����E;k3�$��ʞ�lA��i�)�^zn<,ӚwbZ^�_f�6�~tH2�^�`8p7ykc9'���y	һ2������V��3R�'��g�b	)zS[;��`�����:D+x5H2��?��ƫ�T9�#��X$��*�?t!f���0��_>�S���,��-���/z�i��m��Ԁ�]4�ɟ�,7ę=N�׵���s���%S�_M�S2R�8ې ~-�Ldü����H�s0�Y���~m[!(ƍ����Hd�ێ������N�i��t�J��^�۩��	֞���j�߾���� �F��d���_��3�1� �&M)�kQ�X�9�R' ]~:aSi��"�ᲄ��G�L��%�Y�G��!JhMg���vDvZ�3��u!yѴ�Bϰ��N�U�4KT	��?����d���hB5��x��֧t��ؠ�B:ݜ�Yձ�U*b�-���K�-�f���{�t�S)΋%4.�*��s��TN����-^��Ix��3�:kM(]J�OO��Q����U��bR�ȵ�0)��z����	e�RK,��)�6d'��*Vv�M�S���\Ј&#ݼqJ��P]��;x�CAC�"9x�
Omm��/���p�2����F����n���x��H�
������ϋ�~�-L��7��6�5Q���l������e��6$,�'�}M�L�s:.f���D�8�Ψ`6]�)
G�]�q&�<F��,N��s���:���u���x�Q����5�پ>tc9��ו*Q��Tx��	��QzN6����<Kɉ*�B��6<+"'E*�ٜ8ә(_�ׯ���$���F��� �F!��(ǃ�Z��= �K��W����gn�q?�I��{(�b�������=���f�(@7������g�a��)�E#�=0�y��0�����+?
;�\цe��և7�%���3Q�����c��y@dlaE��=��X��rV~b�T�r>��0��s��8��	�I�e�h�3��[�Q%3b���(6��zϡ�HE�,Mы�(8��1�W*N��ysމ����!��������Q�H0e٪�M
�ZZ��7hS̞x�	x��wi�����xyG`Hr�!�[��?�� ��@]�����Hځ
��#�o���}�n;[m�� �\�>Bt����5]�6��fP��q���~Z��}ȍq��A��TL1i��)�I��
��72�2�M/��2�u�oh��1f��֢Z|��eB�4������2w.XaR�����8�I���?HB���Ȇk��U�&ۤ(ض��Խ��_��Ґ���v�?��l��zL����J�U>�r��Fax�H5�-��"�o�� �'Mv�"zY�]~��Q�$��P%�V�����"���-�������H��,�d�Q�<ْ�đQ��D�S@y� É !�I�h�h)�@|���}����j:�[��`A>�g��\��g��erĤ����uև>�h$�l�? �������F��P9?2ҕϺ�V>/`J���Æ�W���>$��c(���
�S��'�`Ӿ��a�S(<j;�!�iY���/�D�I����Y����ሼ�M��-�u���a<�#�
���+5�T�W�_vPJ*��,�ƿs]��n����E�������c�9X�7�����p�"��D�	�@��}&���>���/p��5�TML������?�a-� G�5a��!mPW8?%�-��E7%ʐ��M�N�&�}�)�$�b� ��� ��D����]������~MPa[0��-���K3����-����a�#�
�T���G��HΈ~Z��ҶT�2 �ԅ�;�E�J��A֌�U�t}tn��j������Oya���5�D��v�] T����􀰏�r��������0��U�OM���U��
2d�i2�Jn1n�r�s3(�[�m�e���SET�	aHSI�q4������'Y=x�7�)�jy��I�F��j�.+�Yތh�=�k!��[Es���P�|���v"������ZWѬ �Cz��U��tɌo�#f,4)�ae�a,���,ޠoM�h��+Kݻ 
(���/�8z��^lX0϶���� )O�����f �=����ORЮR�{�Ä�]~�5�J������Y�Y�{q��f� wGa�Ԗ�^/Uc��Dp} ��M��?�,bw��u�d��vMW7˨��Z)��SD�8G͡����r�������trI�Lʚ|�q<w;������bm3y��B:?�j����x{A����!A�Lk�.�A�{ dd����I���e���z�QAz! �CvS2-_�v���n��E�w�M�	�-ۨ�c'fTc;��̙VAp�O��X<I��<*7j!T�ln����L_�q=�XH� �:�W^r7�g����t �]�7���l�*��u;��W��T��&
�PiO �7h�@�bE�O�j,jtyN�'�"%�k'5�`-�An aݪ��f�`�Z��J����g
�qO�������l��&�=�Ĭ?�g�!���p��!LU^�����_��$*y�X�r16���o�cų��gU�G���~^��f+-b7�o�Ս�G ,j:\���F���^
��&��U ��]Az�b���u^=�n�����+w��}@J�˃Pc������!���2­w�����Q�c�&cj�h�Pd�+��u��.���E�Lb�26�'��2�+)�}��x�2�o�b�Csԕ��A�
m�#���D'F%rF_�uxok�]�FŎ�#�o� I�g�I"�,����Nh�~7����2b�V�
���F9�I�SL��2��< ������ӱ���R�}uĨ���Uɻ͞Q�̒FR�p�;4�D��u�K�wb��s�������bɕo����P���
����EJ_r$%A�>�w�>��p@���W�ɉ�X`�@����b�K � �Z�)����4�JDR�����n�-��R���eL�!4����#���-�l37��t�=K
���-���� �6�~��\���H��x�+:X�Yb]h֘*c"n��E@�2� �(@�
8껵4�/�Y�g^X�S���w3{:bѭg�y�iP��n���_��.cO���s"ҷ쬅�%�}��C������H'�5$�O)�'l��� �v��g���׌m@������0ĈH�^�ח.����E�*��Q�C1O��l�\�-ȎZ�:K��~(67O��]�P�[���U� _��]�*�h�ґ�f�o!V��w�7��E����c9D���BTJ6�<fӝq������9�A1!�X��8U�M(��"��/N0sx3�y�57S�]8��W|���!��\�&�U�Tɦ��tl/ң���������Ymv%�}{H%J�O�ҽ?}SC�&�Y�m0>�f�FC� J������"{X�Q.s~T��V�K��n��ӯ�`	��n+V�t��-R�"D��Bv���Q����t8w�}5�E'C�&�$XGW��xO(��fE*�,Yv��~��R3���l���qu���
�����q����������8�x�r�����9�(��iPKH�"���ۧ�6��6F�?Dm1��FA��o�p��-bY�7r�ܣ̱V�*!�;����R��������B)�^���3������]��G�*�Z4���=t�� ��zEI1B�:맰�c̗_���D��Fܴ�Ť�ˌ{Z��D���l���7*%���/5��t������E�0O�:��E$��c'�9[��`)ݏ��렼F"ͤ�9�1���׫cԚ��H�=�w�c]�s�6~���S�^�tڵD���GJS����N�����W���r٭�R��ð��~U��4ѣ[st\+�b�d��T�?�?�8`� ����-�/��l�?20Jq��c*��O�ލ)���;{�68�z�ovƇ�"o�7e_ �R��l$W���w٧z��Ծm��"�X`&�:�i�Ous�k?oL�z�>�dB��- �o���b������n��澪@i}�suZ>��=�k@)�t-�1G	-?�+�!����9�]11쥯e9��_�9�k�B�K��q�< �o�̕Sz1�~2�\�����rƴ|[I�	w�B	�Ɖ����I��⸥���R�.Ǚ
aV�q)�^���Mw�C�$�w�=9E�p��'*��D׆�h����	�>��a��Vg#�Q��-?	��B��2��>Mj4L���eJ8~�����^	��g�p>7"���'����>��������h��d=�O���V]D�[�
�U
�Q�}v��HPCUOՌjAr1G�h*#o]�a�m��d���,x��B���_�hl� �EA��ℼ��?�=���P;�������_u�0�aN=��דW���j�VZk0��3T���3��8��,��F�%N����UzY�s�
�[����W���([�ݒ
���>�`+<��c���l�Ah�f�2��v%��eS�?��\���Q�2z �vU?t���e��f�̲�-+�`uI7���o�H�>�Mڙȍِ��J�+���W��M&_�)mY���J�+��:@c`k�s_�xKB�q�	�����@7��^��@b��U$��Gݖ��ͥP$N�O9�d��|}����n�⿚ZI��^��8�K�ؚ��s��y��{�	�(�L�~?�W?1�SX��9R��a�LR|���<�P��}5�R�bF��J�6M����!?.��.���Q ���y�T����Fr�����suנϢ�ѥ�0��Ri���xvY����>P���D�#�s����k��47�u���#&�6�PQ#����y)�oD��e�|�u���\,�^����a���y��ڰ�b���Ȫ��Xt�g�7��e����m���5m�n}( Ż�
x��8c6�Z��ʎ�j��n�j<�)��)�sW�Db΂���{��Q�B���Q(�zT`�����D��Z��s�pA[�wi �)���\9�\�G1�� '���t݄���:��E��yl��ښ2M��/�Ҋ�S��a���.Zl8n��m|���4ک�Z�\3jjM�W����q�0�oCB`e���x�%O�-w����@���Kݐ���5γ7~�El,��Ry�8���|���sx��B�KN�B�C��V'��2S��y��{P�|U!-�'�}��Iҷ����-9�'���n�G)�j�	�-b�\�����9c�@��C_;��;C����#z�LzḶӋ�=(�?uGx=�7EE).�@����Z�Mf����o��H�`�B�%7/u�b_�aA8mg�U(0�fȷ6c�F��C�J����MBP4gkB��G��l�ȇ-R�?;2��Gp"�Bqx�-��r%�Cc�D\���x��W@��2�p`��)}XW6���K'�g��ќԋv*t�vzI��E����r���	@A]-=q��P��!ܫ��@�_�;��+���@+�k��9fص�{��~T���	#�&� C~;,�lӀ~��5��.c«���Lu�������������f�-fPd�BР`���̈^eʱ��Ͷv&�t� ō��hǏ�Ǎ���Qt�R!��Z
�MLz��>����d��tqzoͯ<r���
٧����_�ۧ��i�3n�1��o[�)�c�I��&���j���oE�h��ޕ$�h��w�0����L�ID#�/DpE�_PM\Q�:�R�������i҂+��!�g��������a��_Y:�Y��"k���&+EG"�4EZ ;G�`Ք^G��������|��GY�_�%����;�R/2���S}*@d5�
��=�39��E�կjhM�^��A��l�g�V��������@��1E}�}_�p.g/#���TC�u��hS���i$�Kg�����c�/0k��W0b�͠c�{AF��$QF��=��|�R(�w�`Ζ��LZ���!�34h�
�y�����{ΙZ')�λ<5772�V�Ey���N��=l���,b�Յl�k�~kث�u����kT"����5�a.	ZJA{�G��K�9�]�&���Fd�������'�)U�"�g�=��bsf�-��F�&4.=��O]\�i	'�;#vx�
N��C'��8ʹ@ p5�efׇ����Ŕ~���8��#~�C���]����d����f%��̘�Rg��H-��1�΂N�t�s��	�Lʑ�������P���s��Cbm6-2oSl�G)_���V_%�1��n�|��|�qd��'h���0'����^�IBoU��� %^�Q�2�kʲD
8�����kp�
m���#& ^��u���5�)`o�`�����#�B�5�	�q2����󏠉G�L�NC�CE"��R��a��m~�L�_ۋ-�Z� �$����0�Z���F.�7��0�
v���6�=�i��{�4ɷ"����P���M�'���m_�%���g+sH�k����R
��جs���2��K0�t�������ܼM^�(ў�)�R�u/�쉛*�P_!kkj���&�˫���!DIc�!m�A�t�+��x�fsA~B�<�2�?{��SF���w��=��:$�IR��l����;C=>
_Մ�I�Q*�HbY
��X��y�h!�hu��Ɉ�Bk!s�,��[�ﳔ ���8�m�Ra��Dr\����� *�����y=Us:5���Y�W�ŕ���A�~�8F���x���>C���P��� �.;������ER��B��ͬB�Ǳ(������˫��=NHbbM�r�y�����{�f���ܽyF���{�c�e%R%�ʪ����\���a0Nނ�A�}$��P0n��u( ܡDZ~��ʷSpbW>Yɂ!Pp��\MB�Ά|�?.w�.�:8�ֳ��{���p&�hOZ�	4�4����]�	мm�f�I�b�����K>�pa�	�"�hz,
��;��u";�Թm�wݞ.1�y�O�W��=,P�7ūm�MN
	+��6�9s*�y��g]�$�'�U|R�Dz\�-Ɉ�c�ŏi2z����3ۓ-m(����F��`������1��6*v���R���f��.�45^�ء��p~@`x��Oo{�Fu��=y��5�Lԝ��Yp�%v��/X�h{
��T��k^H��񚉺h�����+��O��(|�S&��ǀ��몽t�~=�+�Ee�ex.����1$���7=��K{ûXv(�|�e��_��ﻬ��w!�R���C+����SY�h#�zV��.���D-�m?�>�5���C��g����/���e���G�1��R�\
��wTb�쬇e�=@��#J��(�K\v������R�_��:L���C��oK��p������*+��K���2��Doe8eg��]ܵei)$U���1A��G��1j��~�&�!d;�tS�g�r�ƥ��I�9��f��|���P�t2kQϴ�=����rAQw8'?*�l}�u�oa=��/6*� ��N�n�!�Tm�Q(��U��j�k�ѐB�L�l�òu �7��̉�싟s��@�K\��F�$�2}��r��	�k5��Rs.�C?�pYu�^!�|�-��y�$��)=�m
��vϚ�+!�BY��u���1ޟ4�D~AcD��8����&`#�@�n��P�o���z؈�)�-χ/:|��U�E�dX׳?�����;������£��(���-�����(����9�P�C`���Zw�n����ë�k
���;�8o���H1wa�q9$�h��8���j..�,���/������dAB��W>?�3��b�]y��'t�>���B_���y�Q�����;�N8Ʉ�9��5���o��ύ\�B���5��rp��%�a�C�:7�dV|���Ǧ��7wA��+ϑ3b�㌇���޻�s ��ʽ��N듔�`��\w�K2� k�^�~����a�s8f�0�������R��=�3���X�w�f���uS�1��!���)���r�t���Њd�>!f����wI�xwjj.�\D����T�L�s��-5V��,ٶO��m�7���>>�IA�x��'\�H��J���lꗄ+��F�/v�k�������j�)0R�g�=j�a�x�]���U��\�a����(�/�Q���׆cT�A��p��Ҷ)ĺ����;���t%kQ��b��r#�R���TwQ�rX���>@3�@y����q��L��&�dn��:��Ƞ�<���4Q�$pV/�S�׵�f����̰�0�
���TO���Շ���7��ʈC1� 7س>�0ձ��7[����DBTc?���cz
Z�� ���rD/���;�T�SV�iːՓ����#f$�X!����C`������ځ�V�p3-Õ6dx���f�MVk�]=�ݪ��>����5�&*�æ<���7cΌ�Z?�"o�t	�!�z�XK�Sv0v��&�PP��}V�?�!����p65������j�dfq�Ժ��Y_��Hx\ˤ�:�i�QMj��@����[ȣ�Ċ��ٶ*��p��GE��+V��c�_@��<�uo�0L��l��������K�-KB;����+m�����q�^���� 7���S��q�%��T �+�h?�!����<VJ5���&%z��w�腑�4-9q[-Z�1�R���A�B���f�b*r�F��;��꺤 .h�~���5��O�>*,r�E���nRQ��ʷi��.#ئ����[2X
���)��n�.A�eIH54�%���VfU��Pb��U��Eb�_��5�*|~��pĻ��S�Zμ��/$*h�~J�t�V�*�d�悍�'�^!���&�3��M	9S����-ϤW�2�K1�+�8��sbVɛ���Gc]����Ay�ㄶ�����zgB8;	��K���,�I�p�mHR�&�-�w��]�k��R�}Bh��,`aY����Asɯ����29
�^A�ڹ���f?�
�g8)��Mo�QD�c�y!,�8�������5�_�J���
�kx=������]��TP�y���b���y�Ä�`_�{i����G��������;-j��}1�fUA�:�|S�����F.ޣ��-Y�e��==Ќ�O;|+w��QXJ��t��giJ{5��#��!C����h��}��/h�ƈ� �R�LVsUG,�DK� ��3\7�J,sBE'�=��
F��� �[��(�J�d�P	�b�T�f�φ��j�6!�����]���Eps��TG� �������a�Ǫ�g�p���́�b��U��w,�!���:Q�ŝ%���5ŹM�"A?�o�f0R?4`#N����Ҝ�۴6�}Ԏ/f6���q��G,񂧮4Ӻp�lq�Q�nn�j�|��%�w��z�Ң�H���h�S�^7@ʥPh'�7Z��6�GH��������!/ ��딺�G�����.[ ԿI��TlIf`(K��Mq�>�W��b_�	U�0&YZ�����N�c�"5Z������}!�:+�L>mR�m�6�c�H8�\���t�@a��ktS�}��D�&�^<��?�~��ū&�r��%����e�A��g��d	��Z��z�2�"�� "����:��r�K��l��%��J܁竓��*���D���q��؈���!n�&�������5�̾�Op���!+}�&���0�%A!?�Pg�E��4�
�mć�3��"�=�&�&aB���_J�����Ĺ�({8��t����}�#=!�B��)�>iԘ�҈�r:X~3���1��U�4�R�#fXi��S/Wz[p#&�"�2�Y�t���>I���7*�����҅?�<[�r-�e��1�A^��?tZ;��,���1�]X�puh+"'zq����v��o�*
�f^�s/��,��u�6De0����#����zO�B�h UL�9y��^]�P��1�S�Qu~or��M����}�  A��^e�o�������7/ /�"禙�;Bئ�R�Oq}�Vfʫ�rw�~k�0�l(��,�G�}H���>
�(]�x�_��$�����]�ԇ���Ҏ�&��7�=�"��]��>4E\֋��H+��UB�����q�y��س��G�O����*��kX�d㌜�H���.����12�"a4�@B6��'�+�n�Sl��fUfvK@��������9]��1�����8G�RJ�T̛�k~�����C8�ő���˺��!��,�ov��-����q"���q8P%��$��9�7_��%��x����	m��>��~_܁��v����NR�2Z��`uT��68�l���Y^޴�ep�c�&ÇG��N��0��oL�hצ�ɖ�pѲ~�>�;K/��N���y�.�28wD�{��)P�%����̺��	�(��y�����ҩ����%���42��l�J��/I���.�ɽ����E�K���	%�G��쑀i�w�H��G֘�e�DO-��͊�g�	��e�r6��1ڏ�gL��a��l���
#���|>(��ZM� ��A��-�=��A Y�I�J�0����o����){:�S���g	�x������o~�(�@����^~i�A/H���c�8�'k�%y&ƅ'd�u��"(7u/t���I�bvD�� %kҀN�a��u3p(���Dp��!ʞEǒ۰�8�Ƴ�+�mЀ��f#�6���NRٕ0ߘ@��0�`a}t��K�3���X���[�`i�Y1zA�;gc���O2zz�^>U��E*fb����}n����r�!a*�hfy)U��V}ֽєPa=���m�N�K�4isZ}ieE��}X4�.ɘkސ����g�J~�%��/���aA��nN��v���L���W�3��H��X=�r05,/���:����O��F?��8��f#౨z
1�ef
L���]���F�(S���Ѭ�������`�zbiI�_�K�h�_����o�t9x��W�DR-^n��Ε2`��U�E��TLֿ/M/�����
չ��p��c��9�O��=��
t���8�Z&��7�F唚I5ܷ���Xx������W������"���="�y�K����QV��#��b(3�1���>�U��y�~g��?�d G�����fKF"*(�����.&�dU"!qMyaf�B�����)O	n��4�e��UjSb�F�RDx3"og��#,�a�b��h�{X����<3[�Qcm�X�^[����޴�w�h�{8��(��?5ӸJQc�֧yc|G]�}=�~c����S�>Z4>���tID���� ���pu�5��n�i����2�fGV�}�����`a� CT��Z���b9f3vǙ�0n�(|ט�v,�X�2R=r�[T!:a�6���ad��'<��Z��Tj17IN�?d)���>֜QϠ;ề��:К�NI(�Ƿv���������?>3�NDx�78�2v�Ζ����A�J��@/W_����tr��+�e�+�������wL 6�`��o���D"\5�e���^:)Y�W|��6��9^���%e��Jk�����[ʏ�Ry�4�o��ԍ��u�s�Vm��3���8�-4�b�B�<�� V��l#���^���"8���ǭ�"�y�e�uo�ȥI]�i���
	���:��d��þ�}�/-���t��3�鰉�P��z=ۮ[[w�������y9�}�g��)�{��!:5^T���|^,����;%j~klG��
�uKZ�@��5�㐷������n�����6I�p��+����N%��NϷύ4�V��(�Z��7	�LM�^���U����Ձ���)j�ha�Tx@�Lz��]�n��ĩ^o|��<����{C�\��c��aL�YoJ^2���{<m &m�1<Ȋ%�r`/���u��q�H\�VJ���+,����6`O�?�&{iF��52>�y@��a��ab�6�*:O�s�6<Q��r�ܦ��+�3
�q
l���{��\������X�<�;�[�w��5ܑ����7�R����L2,����+ݹ��a��ELJ]��٩�N-q�o���8�L��!uib�'�v�I�Q���9x��?+�'<D����sH�hg���N�8ݵĭM�f>(�AKF�ң0A⇞HG�D�c��D����lU8@�����ĩg5� Q�|�o�<0y%%1�3�q���IO�J�Ѕ��!�y�6^t�;U�;��:����z�\9b��I�A]P�8���C!�ܞ猬'���C��=T�ʲ�$���H�8���\�7p��*�F列_%Z �c?FFOkR�����)���"l���Ud���K�W�J­i���}��=F?[�O��~ p��v���(���6M���w�a�3�lo�sV��Z�@�Tg�2�à��W���٧��Y-!�d��By��9�J�u$�'\}��Z�6��鋼��ėQY���.p]���9�_:�+�M�ܡđ!�v�'А�[v�v�v�������j%�]�q���"�+kV��b�
�W�E`M�GF�9�_[�����Zw��^7���M\����X ��&��@�a�vJd��Z��ٸ��Q�6(�'���@-��=� j�N�^�~�U��=}�M�_����2��I�`hP�ʢ:�E�\����ȃ3Fw�M"�B�e��}��'x�U���.gR��W?ן���c��&����6ap̣�.�?̮�b5��R9X��G} CA��=2���+���YBH01���:lHo���j�O1�N�*��;r{g(���̬#;���£�����8\.����8}�= ����#잊�WT,�<j{���/��}H�%b(���"�&��{��#و��bߩ^3_��>��QM���!&~-��c�L�Fjn��ؿ&j:R�-r�HnSj������dL�st�Ɉ���AW=����EI�_�'�#�%ՕDb'��yj
�
{���������>�V�O���B�e�W����q`�S��I�z!�0���tj'hhK)GU�f�C���}oX�[#�첥a;��A�'���<�F��AL�*(����'��:���Y��cK��R�Wj�Z���Ǥ�z��S>���T`ݢ-�:bƑI8�S��Q��A�9twx��oz��B�%�UZ t��G�Y2�����8�Li/�r ��=��f{�_�+��3�%|���Is�-=|T��%O��և@Gw�! ��#�v09]�W����!7h��*	">t$����B�,M�\ѧG�e��E��1�OI���9��/���gFo�[��}�nj҄�B)������Ob��K��l���{]w�_�;�u^��v����-��|��xEt�t��>����KG�R
p�P6g�� ��b�mJ+��H�ur���>vx�g�l��7 �P�}#�
����f`�4}�J)�A��n�T���yn�g�Ƕ%���ԕu�9{<�w�ߘ�lFW�Hӡ��v���$^��$S�Gvŋ�Vvj|�hr[�n.�G��E|���SY����!�1˭=��&T���()��t+�B����ݶf���V����7��K��4y��L�(�%��]�"���PSh◝D�h�N��9��J?��b � @��F��k����K
�LS*@H*v�o�!��7�Zן�-�z^iQ�T ���	��>Q�bpYa��N�!�y��ʨ3�g�)yd[O=Б��b�A.�ɜ��7�w�O�~K����#�Y��^��p>���^��'��G�Q~_����k�v�����;��|D��P�}@�_8�LJc"�htb��{Ü�M䑕��:�+¸��s�L��`S��S�I���eqb�Xx��c���y+��EY��W�ge5��er>����vI�4�S�{o��9����ay�����̫���`��/c@KB�K8���	c>�h��GK����3�h��桦CS?e�џ���/�V4���{U'�5�����"�
��7}������"�F VIOg����-g�/��:��P�(��ztO'K%��eJ�p�X�_1�v�A@����Q�s���#�!+F��	L�(��de'Iϗ=��2=���|ݜ5�t_�(
���3_w����<��b�Q��!\�ձ�HEp�Q[\Xۣ;��k`��[����Sd��~�6��8��&2[z&LpY��^��v��&P��zC�rogG|�
�7�`s���|X�U�h:d�!�VǶ=W��j?f9y�RE��D����=�|�d5���:譹��<�����V8+�#��N�?�T��_�O���}��,��A�7����`���fBH{��}��MqҤ$���9>F�'.6�fL���!�3�HƼ��:��ʱ�K�t�V�^!�>,bKd�r�ǒe!����wzĞyx�J���2� ��.C�L=Dք��>�Ƙ���k2��7�"̈́>���Y*F{G7U*���&�;4����i�^N�+�k(���><w9�-?�Ҋa�U]��7��݆n�ơu�\8+$0�� ��Q8���]�MT�ۿ�gWpvk�����r�$��T�G������W�W̽�5�C����C�����_�z�\Y��gW�o�%%5�Ĉ��̀�����C�����D�{%G�-�KJf`v8V��!�dK� �q�:f�T��\[;��ѯN�Ԏ@�\Օ	Z
���zN���'Rn��XGG������Ɣ��#O)	����l�i;d�w=��N��屹�����B%f��n���a7vyl2�-��lQi�	��f1���UO�d]��M��WpǠ���5�ɅG	��?����U�l���0�BOH�_�Ym�(�6��
F�J�G��+��,r5|����?i���b���Bm��")��w��	���>"^pa���(���ш��%=Ng&���r�/5��O/bJy�(C(�m�q���bS���"��B��:��=�rN�gq��kʗ�����j���=�[�Y6X�&1�8
�H����K��6� �o�����ZV�UԹ<�ꙋ��C��B����C�S��^"h�%������雁���0=G:l2��U��;�>,z�m< վ���u2�t >>C~ȳ��*���X��D��{x�lj�������r6?���'�w^<Q.\U}	�RW�s�|�����3�����fX���Q���b�������f��e���m޹����cW&n-��V�A�:��{�2�ʃ��z�y�� �%�Dl��< ̼GG���p��� X��L�+yKa?�R�ƅ���Y�LSd��)�+J4Z��:�J+�^Ӥ�~Ұ���ⷻ>m�N�����G��Q z�ޓ�e�C��P�.���g�yLZ�gDD�Y��Ġ��_	�<�b��ǝ`~t�眲I�:�K��єKv�p�a2���n�>�xl��z��a�}�Yb�Tk�Y'�/."TKǤ�\��'�	���q�R���u��)�t[��=��`{��W��9��u��z�s��:��9��'���j���?�:9�75�LA�hm��4K -�3����%0�������jpN̟7�+M=o�i�oV��{M3����m]x�}����oT{x<��^`����T��O�:/6�09�)> c�JR`�+6��t����p��9z?�"5�m�;!R�y6>_A#Ց�a\���|q����+V+�1�ά���7(2P�80��B_���R�xQ2�рՉ�q�g{��������ߘ���C���;��d|ܷ��*Ǆ���`��8�g��T�I��b#���Y����q`gІ���v��021Ο��n��%��F���Z�@ݔ7K�]@����U7�#�I#O�C�����r��!�g��h���uR[H���K��A�O���@O�W�$|c�E \��>�8��~=����`^���pT/�FN"�[�U�5g���0�m��&�S�O�x`F�&2����
w�@���o�`Y �;�3-��-}��&����9�j�� ��+�똕+���[e3�j5�E�X�/e�=�����&��i��{�� ���w?
X���9��:��(_��v��{	g��y/��|��؉��a�����R/f͉;TF�U��1_�T/�܉bX���7��#ھ�COo��T� �7�kf�C$��
�u�y'�@����к62n��*��h�e��E,�@T�&90Ɋ�/��6�r(� 3'��� *��"��^$�4��bn͟M)��X_n�ԟ�k_S4y�>��sW{�ݝ"t+R9�=dvlt�Ҿȏm�ڟ��Ȉ�>�ʟ�4��6C���މs�g�i�`j�#�W��|�""6l:�[���nn�%�x0)#	J�Qg�?~��
��1�	�'Q6fՉ�]�\
9��$w���r�%��a�F�!Ia<��k�?��R�\��}�u���p�X'F�{���y�{)� F�޷b#�*|����;��a�u;�����mE
!j���W�����S�nZ'T�*MJF�Ѥ��EL,�'Y��ߠ/��{?��3�fn@��K����8b��.��|��+jrtd���gJ*���R)M�P<;�qvCz��G^��x@������Khg��D՟�T.�Y����X���#�E����P#���(/�3'�3 �j�l�A�:���1�!Hz.����EK�*��R��"C༉��fcj�L$��N�#\iu
k!
��[��-��lڅ���M��,9�������-�Í�!lƹ��_�M4zu�Ag(�A���k�����[톞$P���2�~(:�c�[��n����W��#뎞���  �
Pѥ�3ږ�  �9j2�_��%',-Co��hE�r�p3#fb k��|�)r=Qp\�6�j~�b�*���<Q�#�"M�+ca=����{}o�)�I� ��]��ј�Y���1-����K3)$(��4v�z	$4�\�ޞC�~����S����h$����{�'A��/�d�Mڮ�}0��ק�O.��7�b��۶�]\T���JЌ�TK� �.��~�.8!���:���e��(�nI9o	vFn�J����'��*��&�X�����+\���:���;���J�Qld�%oLpj}�����x��P��1���2�0}0���@>��mm!���L��ߞ��6�]� o���;D	b�*	}3K2����"�{]��!����l[˸�Ub�HCX��[��Xc'��p�p�tְL������J�\�������U0��K��(��E:\��o�B��`'���X�[��7`��	XC�4yHl�K��G24B]pp 0���Cq�N����V"1n5(ў���R%��+;��	��t'�]��w�In�'���8�,�X�T��B~�-�j�/P#���w�a�]Ż��:`�X��Ѷ`��@8w^e��E�"qG��ϭ�J�C�@� �2x�nY�� �F_L*��^�3����L��?�dbY��H6��"�^J)����_d:�IڀX�-
;�孞΃�4p�%(G5��Ѵ����`疎\ͩ��ə�J ��zg\�]�Rh%"&*sA�)&^�`��o�t5�WO���H�3�%�`q�=Z;��D8�� �R(�Ͷдh^X:"<�и���+�X :H����>��X��M����6���	ਠ�Xz���
29�|1��5B�Zϫ*,
��=xOÄ0B���~���,��?��;�m�E�!-p�E��H@{R�bg8�:nf�k�x�����y���Y7*6���������w ��<e�\��~B��cR�[|K�DD������g�أ]z�f��޶��	��Ҥ�!��г�I����䈰$4MR�����`�/�{D�\T{��2�+In~���ͧ�AW�4!��É�rBF�;��R �~ �R��^���GQ,���k��f�5M�H�$��6@h���=Ŵ-��� �o;�(�@]tx�L='�m�����=v��`�~m�_c��!#NC��n�*���]7`�^S�Y����xLg{��+�\��x%�MS�0�k��o��Ә�27>��K�c�p����C��*o�ǾK��'1�
����K���W��#m�&��-bd�˟��0�S���i��/+�hj��PF�yf=a�%��G!h�m�N��[�>a}�1���@���H��*��,�������h�8gX��B@Z����=Š��3�S����� 1����|���t�����rq�s퓽��z3�nB+�y!����T{C���`)�s	�������J�f5���8�OGߐ�N`vB�R\6��:�˞h�d��.t@�s��fΆ�[�'�?��t�e���rWZ;Y-o_U����>����R�����\��4Ҳn��i�0��pt��!9��/�i�+�a���2X}׭�$;�h��q��U w��k�}���Z�4=��lA�V�'�7	�I��ǚ�0Z�Z2y1�
�h��;��y�D�lV3M�i�/�	�;���{ⰨK[���[	מ�9B,�ˑR��I��$O�?�il��C�$�0Ӻ���8�
s�2̚�uD���{��(_�/C�Ci$�ui��t�����p1~�k������"��ޥ�O^	�g� )�!ފ�U��:�'��?2S)��f���~��~�?�Q3��Q�8�\��D��5t��;��܊)��d�%�M�J߱z��#���Xu��
�5�ơe��7���kE˶[���1/��x�}�UR�_�]�����خ�u��u�2{p�q���s�(;dSED9�ub,�i
~h���&}]�P��5.õ���e����wq�q��S���+�~�6Tv�'�A�.9$�����e�3�/�f�L�7�/�{^ɰyg����ģ��~��i�~��p�L�[�*a�Vk�"M{	�3�޳�ʡ*��p�^mF��n��o뵆�ΡvjtD�)&ݷ���~C�p����ߐ��R�I��g�-�O��p��$���"j&mP�f�Yhѯ���3�#5�1Ѹp~�A8K��Wlcu���ę�?�_�לlR7�
��I�˖d��m<�h$�QIH�iA�p <�8�d^K�!$�b؜���:���쾡|�
=L��F/��B���Ň��?#^��xߝ
�Հ�]�������'� J��*���Z�V�Ư+�34��M�����&WG�V�ff���h	!�7����e�K߄�]+�p����&A�!z�u��U���_��9)�51�K�"�VY�E��<ݣPPh�xC˗�2�zF���_��PL���Ю`�`)!�a&���<�x��.Z���|ÃA_A찷��~��;��2=���Ю{O�#������Z�B8߼��L�����o�^�j+1H��a��O��,-���Q�f�wg�sAԼ���8�e��z`����q��� �؁�.��E�g�3H4Ry�gz	��<���5{R��n�5��r��\Xr��>f$<�t+��6tx�
��C��,9|&�Z(������_q��C�k�*v�k=t�R�̈��D�}����sJ�b@IxGZ�R��&<:$�ֱ0S^��¸U�b�QF�����WtM�W�@ _7X����f�����rdt��3�릒���L���2��#Z6Q���� �D/�j76?���+$:u�e�C�Ј�G�&���h���ۜRJ�f"���&t�ϖS���B�@j��g�������L��~�.R/�By�{�a������v�K+cc�#}t�1bH)P<I#ϋ]��;I���u��|�'����_� F��\��m�Z��T��F�	{FZ��	�"��׼��5�f�%9�v%�G�t�s���ɃWK�iQ^��=�n�\N�\�N����r@7�Q)�{�ݪ��dWz�y�g��:��.V%�l��x��0�By�%&�ě-䏮85��ϯ���OȒ��V�WM_g`�윽���u��'C���H(��ru��#�Y���=+��u{�
YȘ��@�=�]�ҍ���L��K�U��n$,�[�_��&�1h��ҵ�ۻeů+.��EwQ�Y5��" ��gGf���ȣ��54�h^�gzf�P ��lFn�N�?Εc�o�[q��V��+)�R�bs	�Ea�,p�7�+)�JNBB�,W�u�*��:g��p{�g6�/�|���d�B��F�'7&�M� �pǛ�J��E��M��꣫�`������pZ�j��wri[eI��`3V1[3��}e���=ou=�[*���UݤC�[���T:�I��델�K�bIP��>h�c���!��8�\m�7l��� j�f�2y/]0��z�Ik���v�o�$ҲtYY��N�`����&���&�"Z�N��O��.7'ѫ6�@�'Up���߈k�JĂ;�R[��V�1���kp�»~�E�v��9�!��̆B�~3p�C49Fd��h�n̔�FY*K�6-�H��,S��W��_I(w���tǐ��b��c6�)v0v�i	�9S�#�:b�G+�v�p�
P4̔�S�(꫃��G"ӈi�<H�ky�P�P}��.���F����x33?�Һ �T!��N�� q�=.T�{� �x]j�3�lF�
=-֔	/'W%�;=Wi����)'�~ȑ����~�&y�dV�'����(����G���HmK���(<�~��fY������O 9)�w�������!N@a(.|xu�R���"��� E������7� �E�'��-�V�ɖ������!�)8�tU�[ˈ>����>h�OB۾��}2�#D�yuQ�]�g�=��#l3A�X6`��F �	��,� ��d�O�'�SE�]�;T=�^]�L�3�O��)���mk��|��rX7WQߎ�i��-<��Xxj<ű�/���5�b�!�R�,�䟦�W��"��(Apy�T}h@ɇrE�`$X7N����<7%�B/O�L�QrxĎ�H}�����hB7\�`��fjW��|���
�sOO�.�[6�z�J!-����̷�Ћbq�!��VUB��)F�9�X,�����Qh���|����EݘM2a��8����Q�8&j\�?S��R[,U1�X�
}d�n)epPI���>�7,�aTB�jHY|e8V��׃�Eƾ���� J�d��W��	�)^��rm%�C2�sڄPB�k`* �`�Q��	�?�}l\��F]U;�#���u(���7?l7�S�b �')J����!�̓c����At�~[�T�1rH,�bd���닕�}K�ڱ��-OA6P��:�;��N�_X�"]��Fͦ*<͞��Y/��K��e�[�,�3�K�M'on��"�3����H�jX9����ھ/z[���T�^�Oo3*5�� �*=9w7��Wz�M�3�� �8��ҽD}��
;h����a�B|�X|�3)�@�*ם�;O�r��8�bX�ah�{�`$js�s�����*���n�b��ui�gv6�-τ�'��e���1�+�40���fdx$d�ӄ$ܜ�˟��	g�����Z��  dY<���-�#$tZ+�q�(��8X� ����>΍Q:�q.��_J��6��(ujw�X�a�	��]���i�3Ls�ı"T�=N*�����b���p#���B�Ph�nbn�7�t��hL�:R�Q��1/�|.��ԏ0�3H\
���?L{6"�b���2��ԹК/:D<�F��FЃN�Y�v��r`�a'H��P��	Ӌ���x�w�?���]����c뮺�bY[�О���}	+�/f�G�L},"�^���ɻ�g�n���;IF�'�^��#���P�CDu,�D+��h�_�0p8�>��u�{7dx��2 �4��)�m�����Lv:Z�4&�Mݻ��c�L�ǰb!PU��ˤm?��9C�ɜ���^�_9�j.}r)]����R���0��="�^�&����r���Å�tc���3ˡsHEbv1v�!92"̓mM�I2[ 2�")�a��a
�z�}�8d��@x�ۻ���>/s"���ԯ���{ڎ��p�I�N�>`�~���y���t�j�ϊ�N{K��� ���*J�e߳�zkKz���Nd�2�t���G���������W
K��d!�t{(�i�	,�6ꫨ�:[61�t�'���������ɫ4�j$-�Lb�̡MU��>]�� _
E�.\X�2l��b\8t������k�B�OB�g����P�pߤPőI�&�	}�ң�</O�}�OnV�N3.oh5�r���Dx��q�8�
�C�Fhl�t�$\�&��Y�B�ʀ��c�y�8�0�ȝ�)�ZsL;�\��W巏(����@=�ǥ������R�Z�$����yV4�C��/�Z���C�?n�1h�-`��,>^�<T��4��ӓ9�*�z�ҽg4�Q��κ��w��3��z��M1���g�F�C�εU�����򕛭����rf&z�"k���w:S���y��'�Mj���q�TJ"ƪD����0guR�=�.�E?��F�λ�� �k)�l	���C�\�g�v��P�ԭ8S0�
�5�4�ѫ��y�9�B}2߿�?а3ިx���x)$�(�#!�Ė=~��"�~�9Y��]V�|�A�i�.Ţ2-m���OYO��4I��e��?	{ۋ
��C�Z�[.hO"}_
\a ?��6�J)�4˴�T=O����ԇ9G���Cp�W:�y����!�Z�� VЈ[t�}�]��:�0��K�#ķ�dt�h�6�%+S��6c�|�����?����P�ϙ��� F���q��zY]��ˈY�B~�)艝P��J�Q$T�c����F) ?I֚��y�C�g�C�������z�9Nb��|=y؈Q�g�}
��'Eέ���p�$2:�Y=���*�d?��n��V�=��s���>��&���_T#=k$e�o���� �Ɵ��7��~�~�'�VNLV4������� �xoH�k2�`����ղ�46T\���$Cqs�
� դ˪��"�tE��;ZX�~�,u���U�����z�����	1(�v��9J��&%�ŔE���3 S�i���*}��ׂ�ۄ)�Q��heϸoc�����(b[��B|:Sd��XB���M�VJ���
�����pA)I����Lhܯ<����|�=�x��xb,N��=4��q9S=�e��߱��{-wK3]���gO��7ꅃ��9��_c��$��I5�MW��^k���G��\���a�g�*���~���Z��fƽ�9._��5I2it�k�Í��u���mj'����!�F�*�ފ����H4���|	��]~��)��ꯍ#�{�"b]݋�:7H�Gwz�y7�Yt�O��q��8 1dw��(Qz�ŋя�3���f�=^�j�B����P�Fv$A��O9��a�}
�������1�G�Jܧ%�a8�C�^4k���7}~�3[�����8&�6L���K��K�_`7��8���%��%ȋ���ޠA�*i{���[s@�ϚK0�M��o�1 �"CT�<D��P�����u���~�^�yc]{��@�j/�r�<�X 8�����7���(���:���ze\���v*5�)޸�1��إW�l�B��EThe�0�L\��M�#�O�k��d,?ya��΂� s���W��7)��-���N��0��Y���P~+I�8�w��q!^�M��D�y�k��ߨ����r%�Ӝ_��!t⿓v� ��i5�rv�_���^��{��]R�JZ�� q�(��NFbEz�͙D"���,�]�������*�oγAhɵN��o<k^��=�ϫ���C����q|�1�j�F��ah����6����\�遬o	��6��x޺�+�ز�Z�`(n2v˻37'��I�8S�Z.�ݘId�u�EFć䒜�֎9%�H����t�,a�[�!>!��9�3�M��W/��M/��ȯ>�'�־�P�fy�cOt%��Ƿ��m�6������7����E�`X�v~2�!B�Y4��hBn-�)����ԃ�T��.���E���x�����FZ� �:�������~O��O]�����jhX��c���hʰGD�"W~!���gO��H��ܛ��ۈ���,�L0v�E2�y���HX�2�/���B�P���qBmO2�P��i*�3�n2�&ջ7���&�B�����T@��CR�W-7
�"���m�i�����Jt��õ��K����|!���g��|t��C�d������ڃs|��gjߠ:�iu6��_�Ѝw3�D��T�C]��!���'�`�y!b�>��,������Zb͗���;��r!���@�@�w;FL�8�m<�W�I/F� �j{��շ�;�YH�*��(kC+MX�*�X/�^����g�[g^��	������F�K�HF�<U��َ���p2�'�.���˧���t_��ٓ)����x�i,������u�h��ܔf_=."��6���j��k���ײc����R�?��3{��mޤ�p?�h��	Z+�<�������\�yn]&�o���IK�#p="~H�4*«��´	���
i�U�ү�Hˈ:�-�d74 {�!�&ٱ���:��P��-����`�]�����D�7.xWզ�̩'�[�w"w+�̪;*|W��?c��e��������~-�mA��Ts����<z��=���);{�w3���O�W�T���P��w1��lGķ��0�w��0?��sqy��1�������c�g,o��2^7�4_j-Z��& ��k��-B�$�&-V�����UsO�.c5����<,���>��&�7��s�h3�E�QQ{�d=�KBeA8k�����	b����d ^$6s��N�m��9��ۑ�D6ׅD"�;����\��Ie�Aо�$n�+�O .�i�u֎þ
���Z.�=95c���B��潖�9��Ԗ�I�\-��k��S5O�����Z.���L-k$�]�O!���@�8�����|cY�ۓ��T�ms@%�8���+$�/�^n���-�h��H94��l�W�Ah���)6�=��`�=��	�@�}E���6��Ã	B�$:m���*'S�0/prI�f���;�~�?��A��=Q�m���A�!,T2���"As�4#W�ݡ�c`1`������ă�c��[�y��<�*ܳ"��KTB�os?t��ܒC�`�;vH����mp���w6��ޒ�FD̅|�Q%\I�4'@hג}�%7�8�р��2G�F�a'7����N[�ə�A���;p�%�Ir�6f�(C)>�Vl�"�\wLįV:hB�k�M�x� �J�jJ�ϱm�z�W�����W.�a�P==gL~N��l]�P��� bE%���3V9*�fB6�Ko,��QNb�U`��P<��xi�j^�Ӄ�/t� VQ[����:F�$¬U��Zb
����V��8E4��Zu@q��C@����'u�������������A�ڶ\jq2d:���,'�{�q�Q��f~i`���^�㍁
4��+�v�<�>yVY��#s���^��#�/��h��N5寓��� �r�62�EZ/�P�����Gt��1V_fKmr�_�ޥ��~�V�ז��q �r������?SNd6���! B3Ld�PX��b>�<�=5�z�sU�ޕ�7��|�n�K��XQ(��iUN�2c�v�ߠ?�����>�$�����~��4%ɼ"���[����P����^ƓR�}�`l��~���� ����ح�IpE��7}]���E��طu����2��u�,����ɯzzvc�>fI�s�/J��q���<�6�%���#�7Rƞ~�W���*��<��SL�o����/�
ﱴ���\1�Z��)�C9wN7��,�O���s�s��MO}�mO|�"n�������!�����!�*5����H�z�oZl��w�T���NͶ�3��n�²�������B�G���3y]n�m���s.�Z&����V'q�8�2�Ǎ!L�G��p�Dd� su�UT�qScv �8e��\_��P���S�dOJg[��[NG����.���b-3���� �ǝ��B��O��&�H�C9k�/Gh�d�:_�.P��5�^��2h*��jN���� �2�5���+�V�M#��V=R��z��3�Q�J���-u��8���{��m�Q���"_���n��3�C9ŕtz܌�UK$�uQ6��`�~T�JP�U��<�2?�G��G8'��	�7����2@}�!�i4b"���)����M:�Zz34���:ޱ6d��b���+}�߉h�}�U ��2��/�C�zq��^x.��q�e+/�cH?\�)w����r���w���Nyb��R�6����˺I㣝=Q���pj&��8��й���i������+�� qB̽0Q�{�W0�(G�*��Pzx"���{4��V6�^�[�Z�O�=a����`C�}}�+�Q���-�+�!�C�[ ��t��pf>�YȔe�I���`]ɣ�RO�����H�5^"`���vϓ�b����<D�?o2V��oЌ�o�|]�5��j�b�邠\�r4۴)MS|�Y�h��i�s���{�`��hΔ=`����f/C$뎋�M<����/f�be��/Wk���s赒�嬏�侽�>&p����#_^�H#��G�7nu�{3��pdz��
�Ԇ���D�<I��6ci�~٘b/e���#���6G��|�Ϝ\���/80�V�_�qR��~M+z�j#�h�@�������Rv�B5��b����[Q��8��JɄN��$���@2,�[F��78:P���7��`��A	��g}'��Ҿx�"ū�՘ b�_k�B9�)Z"+�]��=0]��:Q}���H���!�������eV.DG�؋��Dm�ӄ>v#��1�f���U�ZP'��3�N�0-n�V��_����O�{�?��4n�Β%H�/nx�w�Ú�
A��i���Ђ�ȁ�m���� �Ɩ�����y���Mǲ�n��y�Xl�X�"U>\��	R����k�d7jU�B� &��c-o�BH&�a�lc~�5i]�+Vr�ȸ�ʋ���:�X����<d��Ef�'��&P[�,��v����)�`�o{:O�m�;��P�W_�2l>� ��x����3F̣�����QL|ץ�~Ӧ7jkqn��/�����<��($�˰hS�4$z�"d'���4��k6�IU�'�Æ�_pR.�*tU�|���ks">#�*a�ݧV*������in�$=��b}��Ԁ��2aC��g"E%�[EO����Z��-�3T͵ͤ��_-tI!�]��?��i;�@j�7�2t
~��	=sC��M��2��NwN�n�0[����R�54W������x� ���+�BAߐĖ	�q�ZC(V��/�@]��vT:��b�}�����������"��}q���Yq��}�e-�	!�+���+Y�P]��|&a?��GH��࢞�%lW��d����ը8��^(2��n�I���t0�Q��N��*]��^��	�/��?�?܋�5�����16���5���GB\���R~ͬmG	�s�88_�b�arA�\]�Qk;I9��^�qJ��*oa��6���`��╿金(��M�<*���~���n#��P�H�! A����?|$�t�𪴾؜�N׊���G�)�m���^M�лK����>;�B��>b���}(�JL�v��y����.���<dJ��ۦYB�f
��I�o�`�":�t~+���	��6>A���T2}j�r.p�������A��7]Hz{�]?]xf�s�Ť��DR}JE�|�L�������p���|
����uytR��~�~�&��d+�8|�?���.�����Đ���!VK2v�YB��ں�p�)���`��! l1��/�D�b�_���#[B����č|ߐ��p>)��F����\1���	+	��c��}���Bid�����T��2r ������8 �F$!��Yf�*�`��/&N_�1[K������u�O�=���_n��xE�a�����y�l���%�.��X��?^#�*t!��M�A�� ����-+�-�Kw�;��E��+��帉��4ђ����R�q���jv7@2*����`���*�.����i ���4H��C�N �V�`�b�� �9��Z],�ؼ����v���l)��ƙX�U���$d`bA��0��5�BT� 	�|� ��Z�qq��_��Eȓ��=��(�;��8�=�
�W�(��l��z�ưTL��,�9�����Q%k�Ό��k�$r<՘�骢q���X�A3<���d7ީ��r���7��"����/n��awT�d]!Z�Q�|���4���n^lhdM�&4�ٖǵh)(�h<t��TI�hk C3�Ő�pD�!�#�w(�J	36�m�n����5�������"��P����<ߒR�s��I~_1Z�v�(���MU��2Y�5
fk���cNP�����Q�s��t�c#'��=�%wz������L��a�8?��t��*O�Y�@�6��'�n�n~&�	2���Om�\�k=|�lj'~h	������[��t=��&. �!@}����9"�ؾ�{�*U{����1@����P�>`������R��M+w��P��A��KnQ��C�Aב�I�t��e��S	^����.��P���I��������+��M3�K��DZ��Kf����s'�wP��.�S�C��P�K2�5F���TN��p��[k(+� ���ȝ�S��ⳃ�d���4�B.��M���!�	��ybjx�ʕ����b@`��+�寮��J0�����@kٜ޴�׾�6���90�nMu-�f���^�0��5σUvt �r��|wL����x\�,ؾ�~g2\�f��$k�a�z��+�����ŻU�z"���i�G؎#�����FԔ��Dt%��kH"�D$��K�M��Fpё�n���.�Ǚ�ع�忿hP�3�rheSZv�MU*
$�q�6��+m:p��\%����l}�� o���@�s�(0!��H�}�$�`ӂ?3̒S�����@����t��<�8�\K/�X�.�^&1Ι���or�z��߅(��Wd[^�䷴�Zj��쌸5�RNƖ6GI�2�J����X8�;st��u��V�Ӄ��)0}�/0�����b��[F3S��������#dv�� L������p��#�,��4��ٕը�7�vBI0m&Ϣy���FI�
7�V.��'�Lꑴ>y��dÚ�(d��8�,޸���[)A9�`����^�*v�"IU��'�&�nY(�|G�`{V*V���pG��cpN �W=��{��t�CI���uV��L`�7������܀����Rx��#��^ů��m�i$q��������]�Kɒc^{<�E���������jڻSgX���1��E�IIhS��;Y����>�I�	^�胦�j���Ff7�C�b%0�ڄ�\����L,���E�'B@x^Y�Y	�*%�#�l�Y��8�e%)��G�*u���`<��)s��8��o�# ��6�v����2��>+�K�lI������sYD�d�O��ً�����9 F��=��8Ǫ�>U���0l�[n�����7m Ѩ�f�&>�V1$���6éwH��v9�ƪ�=1����1뜈V�L����˼����M�׸�Y��(����Y_��b�H�F|�j1��G�4%R��
�^�iR���&�d�_�� ^(�fn�ѧn��I�>����;gkB䨕?<�m��ç�>D�����3��J;w�rW^�TQ��_G��{��0�j���̵cd��6��
� �;�c#g%��<�'bڹ%����0L�֋-kԹ�'��2�l��w��=e�W��k�пm�(&�u�=�I����9����5�?�V���(�0ZuTC
����ڣ�8�����z萏L�i�R�W�e���Y]�m�f-T�h���*�0a�Z�2�M�3���<�+�Z�s
:&������X
���u<�F���v�]�{Ғ�,��9�EVE��({H�M�nVJ��I��O';��;K]������IX������U�8���m �.ʈ����7��Kv�J�X���Cv���BB"���.�ڹ$�o#4���(Z(�R4�j��йJ��э�|`ՑY ��W��/`���I�������#�`�-��@�S� Im+ڷ�@���Q�U��r̋����~{�.]S\c�4}�������Ј���Ch3���
��K4%"���!P��n�5p�44/�8��RG/'����m���MQ5�˳����yDぎM�@ͺ�q�Ϲ���ٯ̚0:�Yƙ��Y�6��C���B�����wƶ�_b���i�Pu� ~4�K��S�"����#��z6{���%�#	"���лn�=s��(�����D��\s΁���n��`yl1N���"��^�z���k��l��YGG&gOoY��4��]��m��z���B����5�f�oRX�s&l4��/J��>#�}����P5�/1<]R�� �05�un���@AN"|�2�`�$���|@��z\�$�1.�U�|2��}K��q�L�1+pe��������de�"����y�f�yjH�)M�qq�2W��)�$�ғ��������sD(Ce3K?d���	��#��3��t�!M��;X��hm�H�E�{���@i�lk\���yLDs�,��^0�}��o"[��?Ѝ�RJ���.V~�V��Z���L�h+�%�|���b:�[�ae<�����7�E@�
�S���B������+,9��\S�n�'�"x����Zq�} �S��6�T|;�X�
�<��Y*���,K�=�Yb�i��^�;aS��2�ʴ�|m"U/�p���3 N+���d)��l@(]�@2@^H��Qb�ךj�s��Y&�G~O$����x&�F
<���2�%D�z5a�G��ч<�s�,��;?��&)���ћ��e_�}\�u�q�e�B2�ý:�ۀB2�+��G[>�O�UW�����O��r�Y�� �C��f'��x�v���c�|���:�-�v޻�>С9uR��q?�5I�ȣ���Q*;M{@��/:6SV?}�?�|g��vj�+)��G4��L�v���i`%��7���3C�M�y�C���1��/���3ԁ/ƼK��؟�Wp��
]��T���:� H��4�:�AĵY%�65����q�Z�&8`�����nyiX2*䩯(����]Odo��F>�(�J�>c�}����(��j���* �H��j~�����x��f�g�B�x�=�XθY�^�f��-�?��tx�#	�����v�~�o�4!��ϐ�?$�<���#u1�P'z��u������UjP� �o��G\�g�g�9p��u�zDVl$Ԣ���^��p�zv������Vn>U�#�*������ʭ���js�=�g���v�=�ى2�-��螇��,x����g���~B6��Q7�"-����4� �So��ϛ2uƦ�	Ra�yJ�#�2�� <(�)�o=oSL#d�P�Y��*�ԋ�9MO�惺�/F�B��J��A�P��� y���:��6ˬ����p��\ޏ�L�+0�xd:!��e}^{n{��Cl��"�cIE���B�ß��P�R	���ŀ@��h@� K�7�]>��2b��ڭ���?x_[.�O�ܨ-.���H5���߻�m~����'@J]��z�81s�h����
&G�_���W7`�c���_�y,����8JK_��� Iw
�R|�����e���Uc����ɣ��G���;t��0=]�ӌ�;��q�I�Fyc�X���cI�<Y��� ?BI�Q��;N7�����2�?�O��"G97��ܿ4�2�?mFa�a�͇7���/�t"-lIAf�?�N�l@�BC��@�/��s�%��ׂ?L��}Y:��G��=s&��K���r\�E���\�
M�kt�k�'_P�UtWt���\*l��ɜ�F!�ґ�E<2�Qu�x��V_']��c�ȒK���Ӓ��z����)��n������}�,�;����P��Iyy辔�+h�z�b	��
rw)"�E��P5���I�%6:G4;Z[@��)SCXI�H�<�0U'6�@P��uc�!�/(jSR�|:w�~�h��2�A�fE��N|{������!�] N����W��`jf�@1�O�u\0���Ay�U�����Jj��b G�u*��OS�~�� :�s���Q��a�[�`LTd�V����u���Va�q��+}p��*l�´8 �������:K!�l?v=Q��s��%߯�R���$&<�Hݶ�h��-@�&<�M����Ue�r|92%eso�-q�e~��j�Ȳ�"?4�8��4�)�rm����M�}��q`�D)���l����w�Ec��P���x���W@\'�M�L���@�-8A*%�6 `f1 W�GQF
=��`��b9a&��Z�/�l��#0f��'J�� ����J��#�"�+/��r:�@�h�:?��Ԁ[���Rw�{��.5���H��O�&x��w_��&-C��!\�7�i�3��w�dx�ȟ1�E8j8�4�|(H�E�{��I��C��VOe��H�ep���Dȟ�x�-�����Zv�iZ g��_�]�B�@���V��sfJ�*VĸKu���y��XGe��Z����7"��8T�-+ី�I�N�|pM����A�b�`F`3.�5�V�TE�|�
5����,t��}��	>� �k�.�n,��Z�ݞ�#��W��
�.2��1qw\AP!A��e�x���JF��-HLe��P���g���8�(���2}�ؠ�o�l�LE�8��]?ۂ��3�h�G��C,����	 �� @��ѠĈΩ�zoSq���4�ऩ�QI;۶\��K�&�=�Ǐ�+�$�/-�WO��]/��K��y����u�Ês.�S6*�?
�	A�O9����%����8Hi[`X��s�K�KG��l�|eƦB�c��=�@�RuS��%�%[�V%؍-���9�Z����;#���;� �Ɨ�l��c�
!H�)��z���-T�5��Ay��w�aj�9~7���n1�J�4%鬝��U3�A�=h"t��ܝL��網���ޑ�W;��^o�j@���-6*ٓ���Tg���mm�h��L�r16}��=�7ܣ��|�P�u)�-6K9�rI鎸��@Ƭ�ם�����#K;~��Ώ�K;R���� xj���$xs���^$Fa�^�ϔ��N3}��(G�$�r����+��?�Oy�k��H�ϧ�~��?P;�g��A1�����,:6�k�ͱ���lC�(���0�.j�/"vS,7�����q槌E�˒{�������]�̎vb4�G4>z=���W��\!�Y��e�����3��zVb-ķ�����W����4T�iY.�8UnM��Հx��g�b(25���W�
�ҫ!V�S@�<�,�L��՝��L��T�c��i���U�~ʭ=<�ʂr�������c?�-Q�M�}�<���',G#g��Pt��H��_(���Ģ����%������-�R�q��ë+��
�~eBw�� �1t�]@��y�/D	�&�[��f4�%�f=^(p߾�}�,ƍ�rN����mS�vBH J$���Mk�,^��|Okm�Şr�%1���"�Ө�e��M�8�W�	H}��C\�T`)<�B��+�-�/�rVcO%2%����(��WQ-Aif�▊]Lᆌ�5ŏ�%At�x7p�o�i|�"d�@|2a3B��aF��%��V��B�fҲ=�1�#o)A}>�f~�����b�����Ův�SJʥYe
no��d��Č���:$
z�m�&8ZL?�>�=��6�ݿpI,��Sa��Ul�B�#{���lB�E�I�>wό��ܦ��y.�Bi�a98��Q�Q�D�7r��!b���KM�k���k���|�uEY��m�M���,�@��!E �J��������D��Ux,���P�n`��s��I��s��_xXY0E�]ki���U�D��RC�uL��(�����𑐖p�Ÿ��$�=3����*>`Gl�҆`��!f�>Lp�b}T��V��ރth�6o�a����߱&�Ն���&�]f[5�j�O�
���U�oc#�lHa�׆��B�Dvaʎ�A�z��P�EB��^je��2|�	��X`��h"�Z=�/��u�n�y�Z������}yh�Q����A!�P���e�gq���X�5&���nE=�b��D>��G��� 0�U\�)H5n6�^��]wV�vF8k$�<1ڍ!96�_H��EW��$�J��jq��Lı�����wm5!�e%����(ՅEXC%�#�U���!B.��y 9�n	�4�c�����.4��X����fÐ+9�Y���4�_��7�o�<ʚĎ۝Ђ��!{�ۘ�}8��_F��Rr$�p̺�=`ϐj�T�3�Wd'�|���G�xA��D8�m�֐� J�<U����`�13��m2�  $V�}����FrI2�m[b��0�.���T*3w&̈́��]u�R��T���=�Z۟���A��_d���{�[�m��)��"nL���P�"4�{��u�-�;�[�Xn!��p����͑�1koB/Ӣ��G��=7���d��,�+�Ѯn��$����uE�Ֆ��,��GbH#��r��D	�0��S�DN��:V�D:+g���E���׀�#~�Օ���;��,Y:Fz��G��(�E�	[:p�+쳸��=}�����k� �.����mFY��M����.�c��g�=I�֊�����I����y�i�e+����>�#�cCБ�w��w��j�Xc��K]�F��:����rI��r|c����d��O�ꘊ�ʊ�7TS�Z�65�W8�ު��tp�4t�\�܈I�,��.�0{���P:�
��[�Yӹg��T{;ߟ��?���%o�蕈1�I{|�:%��K{!��;��u�vG[3���e��µ|֓�jm�j���٪	�w��ƹhy��a�ƺƚ�����A�	`�SӓU����
�D"z]_Sǽ�p����������"�*��������vi2�Cp^O��':��M܍;�v�aQ�F��3�da�����>��b�i�����E��S��k�`2�����¥�ș�)#�p��������NVد������@?�1����,ʱk�L��(�����s����Ȕ�Q�I��Ƣ�����ܧ����d	%�
�[��h����^�6�XYՍ��Ҥ|=*�I�Nk�O]��0��;$��Ocʒ���6��-,��O��]���x����\+$M^Qpr�i��V}x����]��8s�d7>8��@�D�o���0�r�2d���`EWi�4-W�?uj��1*��"MZQ�$���~�����m��/�Ë���x��p9,� �6F3)�2qЯ�kkr3C�X�{Dܾ�h3�cNn��8:S$R+se嘧�0��P���֑$.� ��ɵ>�ό�QOd�m���b8��l��7��Ae�+itTT�I�CX*If�f��-:��枋�����	��j��D�|kh��N�Š�	?/
Z(����K�HU��`6�q,����L&�_X-�E�~S��+�C�0�a^��N���c�%��A��G�G�((G<�&-i�~�Y�W;�qԟv��mGkxq�	�,Xo�i��&��@�;��f/��ӹ�0UCG��}:D�%y�9�Q#���<��KiO	.�i�cx�������Z�YZ�\%f�e��-o5r�>��X��D��QzP��dۅa�Y�+�z��{܀3��*��Eo��e��f��SS�ߖ���x��&�k�Н�-�x�K�L۾9�kG�4�̈́K�_�Oڽ��&��
|;c�8L����-�����(r��+-�#dZ���X�R�ȵe~�deG�+z-~�}�$q����s��2�\\�j�2� /
{T��*�����6�u�O>��(	�8.9u�Ͷ<�#�������0\'`Wʛ'h�?�����HT��zP�'y}Ք9H�5�'8?%U�+8��6�nT����N��@☷���K����NR8��Lotw�?��{7I�2�e�����N(�v7����zP�^p��
�Sy�\�Z ���ն�k��Ԓ�g�S�E(���t�_��}�B�ҶL2(�V�Z5�;�k/\A�����^����@�$Gc�g�7q��pF������}�'d�̑h��$)?/�O�Bw��]�c�d�Ѱ.��FX�Ο[��������1�N���~���9�t�R���V��?���nM�bL�^ٙ��p�`�!.�n���U[�̈́h��($gh�y4�<��#����/s�>�b���L�c�a�a�cT�~O�&�(�:��X>kS��,m�W�3J$Ԓ��Xu+�j�w����1&�]�����;��f��ܛ�r ��X��[�ϞN�om\������m0n�N%O6�� ؈"����nV僀W8�jP�]��f&�®��s|*�4�W��fl��!�����7���]B9� L2�l����<Lc�(�n�h-;�,!�I�9}�+%Y|�-�H�����r��K����|#�Y�p?�:���;���a[C�9��J����$lK|�Y�uW�n9���x;�/��ʜ�"�u�>
�/�ɍ�=�_i�|�6���?���#����x��*�P�p��B�ر���W=ш�������ds[��9�x���%cEM���n��)�c��r&���qm3��ME9�����fx=��#�����3�=�T6S���\?���|a7�g���t�vv�.|:�Ũ�����!lK��"�;&�1�]8�+�����I�ħAk��~�C��MVO*��
Zt:zBٍ`֘�Ċ��"��1/(�'�\�}�~@�z�����7W�,I�ugt���	.��{ċ%�N[;��A����S����/D�4��V�]<'�PG�'+�!�75	8�v�;g��f���7���h�7ץ�r1��}l 2,���&����{�@�j�)7�u�p��[�S��]�?�K+�������
���>�&R@�/����H3|�]�A�܂yH��Bμ��?n��x����Q���_F�y�3��~H�Ԟ��7I6�H-�k��="h���+�x���;<s���+�c�~�Lh� 2JQ@���{ũ�T�2ʊ�.��D}��L�nz;�^��GS��ܪ�O����Sv	�Z$�s5Y���/Af�c	h�����+�e;������-r�*T�)�=o�>?�ޡf��{����y\�G�����+�y�����JH8N�3��Xu��N�G��uDk��ɤ���c�����P.��-B���<������H�.kr�*
����5��nml��W�^�L�d�u�� �]!�������
�K�/�P	���?~Q�D(�9��:�xL����od,��3[�sڇ�@�<�_�Z�D�:P����!c(�J���A�6�f�*_AA�g�\X�2-��ж"v�0~Г�`-����M�kH6�2�Νw�
BG}Ђ��ʚG-�#؈�Y��R���� ����ԯ�i|j�>THv9Y�sԨ����g����2lu5���ˊ=���+`�����'������r�9d�&�.�x(/4����j��u��C#�e\�]��2��5?��Dk�F,�>�fW�<�9{/b	������Cwû�	�$!V�`���x�[��'��R�A\,����� � ,�F�K�d��� �|��ӭ���l+@���5#���煸���2�V}�����������a�ɂ� �͞�L`�9�������K;��*��'��ۘ�q��ah�~&�f�e.�
�2��ܨ�O�.,:���S�Y�!�A���ioٙ@����*������ъl9���ew�z@��f���fdHt�˝`'۞�6��~�P�t���[tT�|0E�^�J�nuT�K�Vm%OP���h���^ְZ�5/��'�tZY�1�轲a�fJ�A����P(V4i����G�+��*�7��k�f����p����}�fc�cyƤԩ3�P�+�)��6&R*��mW�Cy�����-0ؠ�ف/=�ɮ�o[HKƋ��R9��;����E6�qkne�G#� ���Xz�X&�GbB0Zt�b��%���s/F 53��t��"�)��I.�p��i�����-봠	1��z�߮�@/�N>.�11*����6�6���$[%f���Wsj������o�6�CŬ��E��#ꆀ��\) &��U�V����4R
T�I��e�]��4��t�I<̪���K�1�c cQ�zz���ddwGs)�&�]ǣ^q��䇦|�A�]ݯ�0�;9k�
��pW��_6x�[�e�	Е{H��O^�'n�B�L�bI���kp0 �>�3���*�:�G2j��L 0�,Cܤ!I;��֫=TkI��^��ќ��9(�� ^�|�� �F��T]׹�����5��������:��>bP����	p �ٻ��2M1�y?�*��ܮ5��;{��6���S%c3.Z�x�~�Z�vh\�h�ؖZ��O�@ܰC�tp�-d��&&yT�;��"ܣq�����T�i��Q$=L�O"`�Y#�������Zfp4֣2��� 5����Z��^�������V��X^N��-q���ƻ�$q%���[I�#����nGS}��-:q��桄`���ζt�pʋ�K{2�k�A���C��J)�]1���V\\�'�0)|��d������Y���ಭ�V/#`� g�7���O?�p	a��_��+�j��VOs��zt���m�SV��������4��E�k�L�����A4[r��zZG�:l0�U��t���ѴĞ 3#C�ʋ����ޗ��� o��Cw�q�5U�)�(������8b�r����7��ǚRẼ����,�p��� ^��@�$w�%���H	���fb*�����܈؟�'�h}�˰y�p����M��ѫ�8%]e�~�|.8t�y�/6�b*�X-5�	)��&����m4���{!�e�t�~z���Ɔ(��� ��ى��r���nwGa�����cS�Bp8��r���u����*y|�E̅���
⮽�z	^��0��v$�ǲ�u��Kċ!c�E7��	��ZӖ����4�r��h�J�{k����Y;.��ބ>��/�M\���� z�L��H_��b_�҅�cGҡF�>k/�ؿ�\A�4��|F�Bk�B�����*�siN��q9�yB�����/��<2 �_�6��:�Z����p":��?Mm�eEk�"��4..\+�d��r���H���z�<��
ª���8#��S����Y�/Z���W=�Jk�jDt?��lSn!���B5*�����m�
��B���v`t�}{��r�4�;n6�i�mRg.H�$�ˣ���gMf��t'���o��>Z=ն�gZ�Xg���5�/��-�ǙGk)NI>*��2�}��D�+U�	߯�9nŸ�+ ��!揻փ�+jlA� }���c��v����	����$�Q4s3�|P�%D���2�&u�Хè5���l��҈��|���i�|�8WSwˇ��q�o^YN$���r��MN-�'�iH�]�a��L�]{ 7&N]�,�+FBm�u�.���x�n��a#Xd2�P���"͙��ƈ%d�Q�E��Я*ߪSO�{���+�Uy����^�	",o�4d�:��w~o�B����̤e���\�|�^���]�:zQ�Y-nQw�[��`x-��H�_�������quT+l2�\�TX�ʘ^�=�J��X@���l]᭘{�k����}�hP8Q��jir�]�x^��t+�o�~Q�=H�n�*�!=W�f`V�'0�X�����+$7j�8��5��_FB���E�>hC���[����� �����|��tʹ��i�3�z�m�̳~��D��2����^]t6g?p@�<��v��m�XS�Ԧ��|${7���-��~l��a�?����_�-{��U�(�7�4[���s��^�m55C�2��~I�iC��H�jj)m�vd�{mN��7Js��g?Ɲ#�O��t?�]O��&��#�j
�)� A�6%�)�¬���\uS�j���j�����Z*�<k���&�o�qS�G���ͱ�B��+��G鍴X�R��Ȋ5�p�B0�lᑅ&tUe[JW���
�b�q۬#2��ۯT��U�+ֲ~���lŰ�P>n慾���T�$-�ߟ6\�.`����`�B�wϑnw���ܩ��(5'w�@��4�#N�h�G5^��@B��#p_�IDW�\��ᝫ�F�ޞ' �x+�>ǁK�����@J��!��0ٽ�d#��v�tC��޷��-����T�^�a6���>i~P��y���fr��?س�K�۪$��f?����y����E�����ښi�z��P=�ѐI�%JL��Tܽ���S6�7�2��Wx���+WMȦ�0�L������%�k��BU��/�����'gd-�t�9=�

!{�:��S6�3}@:����7���F��ԟ�e�+P�-h8�y���/gG��2�8lC�{bi��(}��K����'!V������c��o��Zⓥ��2j���)Q!-7�4�A*����A�JI�{������(|�)-�v0,�A��5�mv��c	C����0��#G�c�~�^��D�'�A=p���RQ�b��Ov`[����1�T�2��sO=�g=����N�kq7ދ��ЎN�!�������w�E�oz�-u��V�����G��>��%������b1V��R)�Z[뒜��7�:��~$73�7��r������ض�ģ��t]���Huu�B��*���ܝ;i���e%![j�*��S�[/hњ���;�\ ��&&�*���� 5�� "�b��_%��!��Dku� <N�.
h0E�ʰӶeW��SGd��L�;�L��e���o��<\�\�G���Di��-�w�E��ɲ��Rm���7�- �����O���#?���:if���d�BR�|�}v�4+�c%ҟcz��7�2y�D[���I! ���P�"����Nz�ĸ�=����4�j����'����r�A��{;X]�#Վ����u��:O��B���a�9*�����VR�ZN?|3�+9�A X�;!���[ȱv��`��8���a���!�dչH�5k�K���B0���\@�m�1v%���0���������"�d�y���y5����X	i���v��_ls9}�G@O<��%e��|Il�$�S�ݨ�Q.(�vf�꧸�;��F�����r��,�<�񎱷�F�J�h��G
�%F��uAA�Jn�"'i��2؄f���O��������26cXת���u�4�$��]Iǔ��HA0���"7�M�q���=[ޭXc�3�(	�
�{) ��;�"\9t�&����e������'�Y ���vu�떠Ú}
���1����0�y�k���&�[b�A�[��k.-��Cw�Ɓ�7�	O5�����?BC�5�U-"�X�R�����l;�Nȩq���4L��d���O{�{���$�G��8++��`�%�˶ّ�(r��`@T��}b~1�n�U���/a��mG����4�?'q����.��ҳD�A���i�:��4���O}�z��ΫX��x'��ޣ,m{�f��x�Eboia.>7�"��N﮷���۠�5���]I���X!fCS59[jY��aq�B������4�J��w$���\8��'3f�q�Onځ'�[�ۇ
�,�=7�*]�x&ѻ0�87q�#�E����#�q�B�TT#E�=
�����eB��kE�t�K��&�[X���S�U1�^��m<u����`�SO<�"���,��n��̦���ր�m�-�ҹ���5i��C�^��Z�K�`��8Eae� ������
W&=#�Q��O=��鿣��;Vx���� ����!���m�ޔ`�=��%����ЅA�9�M@�a?���i�E�CqA�x
>P��zxx���Aʒ�؇&���P��(�Pg��Vȱx���_Yh�����싌y�
A$V�����$b�l�B>#���A;!���,������t!�^91_M-֎�WQml֍8;�lk�0�,ъ�.({��2��b�-�(��b�����AK?���5��o%Zޡ��+�i'�rj�Z嚏��/	���H����:��ǜ�l����~�Vq�,eh+���կ��3�E���{�Rt>]?+�j�*���б���)���ǽ���~�<���NV�|���4_������!�/��g�+��A��o`��	�`C:�'@�Y�5�jv�N$ǧ�=���NҊ���LO�>���v5~����캆2Hi�_�'ӧ����_Kx/�����vP� ���~�E"!:��3IF�V{��N���h�1,:ה�E�%fK]p��F~ky?����\`�6�2X�1	�	��+� ��йo�M8��$M���m9î��-�J�Ol�r]:#/���x��E,�M�+j��6����``J��1-?6U���;v��E᎐��63l���|��N���|��k�1�첣z����!dS��B����͸�Y�N�O�f%��)�2�V��������`ݎ� �VH��4�L�,H��2B�L�Ea�}�<Q����?C��]{����xw`R���ݨ�r��o���B�.�"1�����=)@���k��u���?ƙS�"��z�i�X�7��z�X,�]�!��B��;�zKZ���⪫E����MMċ%b�Sj&	ɻ��h���5tu�Hw<��}�L�^�-G�+ўB�*?�G�]�r*[��Zg�*)����	��&��}�v�	����I_<��q���ίۭ�=��$.�ژ�y��T��n^�EJs3�-�w�P��(T�rI�%�.V�U��X��3�cW�C���'�c��"�A@|9pow-�l��I�j$m|	4�ٛ��!r��֌Z:�}� B�7:O�k�pJ�a�sP��vcU�D%�d#��"����! :�#3� Hm�A����^�N��C6P�$�E�ˉǰh��Q��X�t��b�ͮ~�\���í�@A�vMJJC�;�ow]�Y�����ŧb<�I~�ޡV�� .mato�������'��@��-��O����rOd8W�"Gb?�Q��(��d<��i��tAk�v�/܆Q�\C
���J׎���}��3e[�����qIH]B^A�!$����q�D ji��B�ǎ�6]���O��ƏY� ��]w��A�Z	OI���I�4ٱR�E�:7^� ���e�Q��;0�l�Lg��i��F~&؞&%n�yY�'i�T�k'���~o���.�_זzZ�snK��VW/�Z*	�9&!��h@�qj/�K�.p��!�������n�`�4�	�	z�(��nw��ܸ�l��^�0�����o���*F	͠���	���e�/.���ަ��"dy��&�`��vc���4!��]�R7����)�G�=�X�b���7�Oq�?�eo��0~�僷~T��ܩ(�6"O�&���i�!�r����#�T%���zr(��&�>�~��h]̈́�γ��͂�z�bV�RW+��f��SҵX�×���ksž�aٻ6K�3��<*̮e����C҉j�N���}�W�M����j�!�S���3�x�])��
��V�����U]��Yvmǟ��="@Sj��b�*�������W�z�2Y�!TM�=��ޤܝ�/#8�0e�����ŚĨP++�+���ed���J����C��b�23�B];�L����0��H�D������x��GXi����"Bi��v�Ytܵ�\�X$$�YR�����lz���L�����fR���������;�@����������~xb]��B.�AB0�@w��\��էD�^Q����˹��i�?Kk�{h\:���2�:(�d5����Ӭ�{W�|F���6V�H�т��D��Qԅw��ّ��3u���2mߝE��>*s��Om������Q���5�����A�,o���!��o�r�mR��N���ͧ�5d���{�m�Tcxb�V�w�Yь�%ڻѰq�(`zx
W���=���ʨ!��C�q�_�a��b�Gu�g�,�,��O�ZV@�U�@v���	qN�E<)Z�J�g�F#�4QMb�i��9��g��oOa����Ư��Wks�.��c��/�\��;j�{*�`���.T����dapJE��%`����(!(�:C��\�
r%���憞�S��?��K�u�_�HQ��-���&�����"n��� �3 d�l}`=�J?c8B���@�=*���?�a�T�]��=_��	��e9�G�R,��f�yp��04�4��}���h��Q�����N�O������d�-�$Leh�ގgJ]�Q�QAa5"��Qe���QA�X��W;V���n��18`lw#�!g����Yg�[u�r$�W�������3/b`v~빅���|��٥d��6�	�?�r��0a3ZXWs�ߐo`'he�U��M���T]���V��;TZ���ًi��P����܍f���PX'\s��*��m��?��4�ɑF'��k�ST��*	�
�H�8��E��˅���Z�a�L�}P���c��8����6�?1� �F��-�@cϋ?���	l���"Ī�����ԑ�6h	�������\!nn6�X��N���ne�Ybj� %�Zy�����8B�$�ާ7b�<G����s� }x{�D`x�K}�b}&���������ԣ�*7"����0V��+)NY��Z��N.��obW-&*=���v'K��4�l�y�k�]4�#HQ_�g��Wr����$�b���n�r��k�`����B� _^y���ӭ�^9�6N�pt+�J�4�.BM�����_�h2�����μ*K��f�f\�/o�7�%�JW�M3�jK���HY�ǂ�?��.ڑ�c'��Z���mݩ��i�^���Cv��Bk/n�J�0�?�����Ndl[���Y%J֑���V��X�}ۨ���(��ĥw$@n��1B������ſ<�=�p����3�Ϥ|�Ō�dƠ����G�=��^���'PVP�B���S;w��U�p�+�B`�o�~�ѥ�8X;���D���<�i0���_�X�E���삌��9��|�fBZ��'�_<���Jg�'˩�:u�p����_�Oo�O�z��y��AH�_��&iA?k�2A/�ȣu��/	��y�+�14���"%;��%J�E^�1���1.�T�)��!A�C������t���5��s����ث�j���e-���+����e�(���j�ݸ��X��3"���4�Q*&�#�SUv !���|�"!���E&� 	0i�N+�H��xP6/�Ć����.Z��%w4F���������_��[o��`bU�'Vd�p�@bEț�L��l�RJc�pOt3���h:y���O(`Z�Kw��o��]&��?6�!��Jqs_���GggJQ�*k���I>Z���P����/�,��
�)ɱbs�n9�H��㟌k�Ե�X@B���"�hjWt�īnF���⃡�٘}o�o^��22M����h~��m���3����FgN�+R���������A{_�(i��C�ML�#�;�������d�Ds�^�� 
��ƴ�8��h������Z	n�KhVO�e��5-"ӊW4P+�9^-�`�*c|S��k"��feU���R�q̽ז3A��bE݃A�N��S�$�5�d��a����;�L1�y�5�-@����,1ƬS)�L6�g0U�8w�U�m�����9�&��M��z}I]U@R�N ��þ��B#���T��ߦPb����&�á(o��,�w�;NT%}���R�	�>��`y&t���K�i~K���n�d�B��,��!Rl�uzܔR��ge�5�D��Ӷ4�1/�ÀEl�R�~��fuU���k�3H�q�[�Q���C.܆<�LX������81����s2�$�R�v�bhEz}��R�vd�ky7��c4(-S�96Cϛ�Lk�������(�U[$5�㶈9	�E�@�y:^�*I�1�#oVi���D�ֵ���Z7���/@-��ٿΠm���%�!Z�=u8�i[��ׯ�y��K��ل.��+lyZ018�*'�h� �oa�7�>�1�bլ\���[:���(��<������4�����k!�'�����J��nK����f2_�򛳡))�8��O�7~� c����tD�{��O,3�J�Y�[�=�j��:#����������2��I�A�����#����x��{Z51�t������^ <���lB��#�5z�fmlt��c���ٹ���%�R�^� �B��v%.�bj�!��.ШY
O<YƯ���>{�ddL�>��JJ�y7�}/d_0*p�+���7(hv�
��~g��;x�"�eL�J,
��kﲰ�O�%�5Iw�"l�s�E'qJ�Z�{qI�����Z�U��f�
�r�m�4︯�os�К��Np�N�*�39����+Q~	v�����Ȕ���� �`7ּ�=�`�+� b���B�<H�K��0Q�M�FR�c'��"�N����@ș4�X��n�Qa�{SU�s2F���(D�~C�C(M���;o~��P�m�3&{\�(�2:����w"2�>����jCN�F)\��g�C�?@
�*%)m,u����ʑjX͆�G�'L[�~�ʤO5�<ڥ���軉�1[o�A@�J+�W�� ���I�5C��uxF�v�^�S���M��}4�!`f4ʹFM�#�R A5�q͟b�Y��Y�+�^x1��N��t�\۵u��O1�"%�!���*�iK��R�.S�O�����)�L-�O�k[؎�n���EN�\��G*Xޥ��%~���ta�@��-�Wi���]��B�!��Q��ޔՌ�V�}��Ӎ�h��[��Ot��!��$5��LHh�䯶�,��#��\�����IA(�	��j�l��$&d��Ss�~_�����B�+ڧ ��<5ٰ���jAqؠ �Qw�*6@U<�t�s��Yv��ڊ���b�>k<V���n�n�7�U[�F�+� ��i��?�ђ�{BR�GzBP4W�W&���s��9�Ŗ!9�K�z�-p�8�QW��Uh'!v�:֛���K�A�t�%���f2BS���Y�}����3R#i��Gϕü�W[&��Wd�hP�`�n
"�2�D�@�m�_��y~
!�1���Kt�2�3��KE�H�p0?Ь��Ŕ�TC���"�4�mW�ķ&̀�(��4����B-��������|u*������8�O��-m��b�����f�I�F��W�^�w' ����X�^�?8P������;7�ɏR�pX&��enϺ�D�>׿��`�fh'� �<����k-�8L8��̸�Z��.���ŗA!�:G�RB.[�w(�0�Ґ!Q�G��~b-y�n{�:�CO,�,�&��=?����[�ƅ<��jWj9���Z@�P:�2xq�,|�����h�6Qgm���{]�V��mL��s7�S!��J��sn���KC �4�DL��k(��©�O�b�z������9$�q�	�Y.ˀM�#��c��l����I�l��ￅ�c��v�B����Pi_�y=�<GZ��������J��5�H�.s-��w̱��3�y�=2@g�aЋB�� �P0�����@�3J��t�AΏg��3��Ҏ*!v�1/��P�j6@_j�,��
n�.,b�]�8��d�7�঩f��RB���~Rü#���E��y���mJ���͂�H���\�Z�j4O���s_�9�є+��) ��dQ��m�{E^X�d\O�"���o�ی�P��f�^ֳ��=58�ާ�cf��j������|̥���C7Nl�K7�<�ֺ>�8�K"��� ���_N��ڸD��y2 ��җ�qc3^	Ob��2���<p`L���~\[��Э�|��VYMޥ������]�%=�tI� {���ٲc"�|�,E�2��_(s�i4u5�
�ȶÍ
�!S�@����Zb�J�{�WA����S@�4>��ժ����wxոm���\h�[5DPDp �ضB���`~[7�p�ѱ{�Ip���Y�\��E�R�-��_�cH�8ƒLD M+�4U&
�;Fq��R\��I��tދ���X��5d�$����%|�qm��&fs.Q���3�Pn;���ti�EiaR�k\�/��?��'3��NExj��`�j��T����;nCD��r�������y�3��; �K�oΔ�p� G��t�'��{��)Qu�յߡL<P��m5+�w��b�7?����/f���+�$A_���\�ߴ�~z��t4}_�0|8)3q�4�g�����QJ�R������u��*��0,+��^*x�yi�)��+�
��Q��ja~Ń�{j׵������9J�8��Kx����f����[����ʤת6[��^�r��09L`�������e�{eR\Ltz��[ѣ���3�yɤ��`�e=]�C��,9�4؍�W�%�p�f����mo�Be�_5,���#�q�q��n�	�\�E0(=�ڞUxQZV�J(�X	Ǽ��+]���d��+v
ߡ/~f���e��w&��H��x�c�Q���<�0�kZ�CKޝ.(Y��Q�X ��t��_*�
��ܷ��M`?��cm�"��Ӆ��-Z���i����S~�:���} lK�6��S��/�JD���,p����%oPwG��Ö��9�7���cj\s���(Y��?m6�8:�*g]��}���Ss����ò���B7K�$�gu���p�@AĲ���rz�ĀOf(���GW��m2~�&_�*Q�=�5~v��U�8b$U%E���3�yr�F% �/	N�ь�EL���K2"�.��Q���\F��7�E�ϰ�|<����X���*DS&1M�3GHi�b��T�Q8���{��ɜ��ꗑOc�O���76���M��6�B�)\sD�|I�[S��|;�j����@�F�W2͇������-T�Em)��1c����@�v*�D�[�0 sc-[�����L���~���ژ�J�?�F��u�����#F��W�]���Zd��@Y|��B���瀈/��*�(�W �`��tѿ�j�;�;A������L��|�"���a���y�fT�ZB��	}�\��q#�c�������O��Y�f��ϑ�ÃLߗ�f�l����p�$]�&{�9��(�]���fXpP茀6��r������-׷�`�����^�h��"�=T�L�[	0���H�$ �~<�������N�i!`�)���͢W<�Xo��u_�j~~`��F�ޝ!�
S�H�u	u ���惻�/�'�u�R-��4IS�~I��W�/���Boo��Ѽ�/�q�/]��4�����H�*@�ذ��xf�G�Bݾ�[b2�4��I<7z��P|��~F��d~5<7~��8�9.�80j�C�ðHh������u���*��J	==�vd��"�n?�Ғ�i�Q�gu6��ɰ�/����&~!ٽ��f��e>ӫ"�X
�Y��*�N	v��Wѵ�����<a��{#D��تf=������d7���P�l(ҷ��X�]�Oܯ��0t\b+��eh�)���"b��B&���bA��[��$6��Nol�ֹ]%����mbW��4V��~��l�ߤsZL��`�f�@a(G!tt���?F�f �\
�{4��ƘY��g��옦j1/T�>c�!�/�~8�azU̐nnB#�x%Bg���x�6��N<��&)�C�fLo����jQ����k�4]���w ����
僩�9;��W��a���!��������p[R5"��+�q������o��y���$�_TU�&�38F�',r��1�������g�Ì�g�f��\�tє���㝛���ȝ��{�����׵-��1����Iٹ���a��)Z�ū���NM��A�j��#J}U��t�`/���Q����ގ 낸K����αM��R{s���P�u����n�L�x�C�k�iEY[!3��)Ӵ7�QAȍ�SI\;��Y��F,B�0����/tH�x�k@����&������~�<��2q�2_d��i���u�)���j��:&C��0(ԫ1?�/f?���rf�� ����q�Ar'�M��Bmy�o�{���^¨z� ��mt��,C����3��L�<�����h��Gԗu����0��}�gF���K,��;��[:�2b�8!��J�FZo՞��uIt}��i�c�(^!z��p�����;v���ך̞N�p=|.ʹ���A���3X 8��ԶXY\�[G�@�Gd#^q�g:3�\oÆ��b��Fv�Pjw����CA������H���#��&&�1yN)nτp8��w�
P��$��3{������C<�T�8uh8�_�Z�<
k7*	_*a������\�6<x�,��w��>?N~�����,)Ӈu-Z��e_yp�t����42z7��bveb��\\rX������Ik�hKj�MG��Q'���"El�s��f�_����{������4�X,��{�!�"�=y�tAf�o���0�k�j=�Q�κ�c�V�h����6w'�P E&���#��w�kz����R7�츆�̲��q�����2I��7̃�@���S>P��ʈ\����2�����1�m���/��Auӧy���Ϻ阔�2!GM��?}���cbq
K����횸6���X#�'�͂|��um܍�+V��S�=��^D�s�l|,��{�$ 1e1�\	��- ���U�6,J���T�~m���`�|�p���rڗ`�<9��7I��M�ݹ�´f^ۧu}&A;�Cxi�C/�]#֚�rIrrr#�|O����OO��?�rp��\zǥ�ex�a��Ң�٬�xׁB�`�֯eh��W��ї��c$��Gh'[��/.!(�(�J�jZ��������q�h��f�� H�.���_�v7gT5�k�m�� ��]����3s�g5�f�YS�3�DY�!�-u>�#[1�h-�N��
Xm��:H-7��"F�4��n�\�+:V��v����#�7ŀ���GYo�D���T��@7���	o56jk�x�j��0{"���8�d�@��k�9w���lY?�L��ebޟ�%B/�y�bPv&S���ܥ6;��H��!���s�*�ao�	�oSGE�H��ϞNt���..�-d����g�ob�lM�w$��}�2L�/��6g�#.c����D�T��^��e<Nx�XU\
-aDW#4�_T\�ohd�t�l��G	OԶj>�T�!�"Y1X:N��{�¶Bn�.�zDMF��dx��&�n�B�F(���#�1z��פ~	�^P�Sՙ͢�G$�����4D�Y��DL���(��M?�QY�~�����'G+ �?B'��K�E����g�}�i�C�Yeׇ���V<��T�H眆��=g�;��Y`J�e�	C�� tAVS޴�����r��Ь�d��1}d%ŉQݍN�::Q�+g�V�|�6��`�W��٪?N�+�K�o�}�<�F@HA����@����*f]���N5�#dw��$`�5�749f��`�#;p����OA�Ȋo�bR1�svڬ>t	��0Z}�U'˔_�#6W�],��m�}Q4P���wC��j ������%��@���/$�ʗ^&[^C�����ҍ��Wӓ�|��w���j���7��.������5�7)��c-�C��e��`�x�Ȱ🤍D�9�*����o@22����^\tz ��Q���z����H�V�-�IN"~���?�;�r�C�w'�2���%a�]!rA�x�i�JH���U��4W��P�>s��������J5y������e"�0d�����Jr_1����W�y��rۙ�ta�D���������G�3�ܽD'�A�Y�L@�/���]�]TM���6!7�U����<kx���-e&�ή��?pvDY:�;V��Q��s7'�'G��:ʄM�Cm��}S��)X*�R��z)$t5�<�K�fJ�����Y<�hRf�Z�b�H*?apv���r�>t4�!6͵Ro%}����CTr1*Bv�7�'`g�ظ���H��� ��`I;M:@�y+��w�q�d�N�g������w�����]��>�^�6Ƨπr'Aڷ�U9P�U������>��r�Y#�a� ��S�r���:W=$~*5�j/������ۿ9T��ϑ�j�|�%Q��8�
K?��b1���}F���~�ɔBZs���С9�.���]E�}3[	xjX�qu�IL8$�?<gXR��O�ue���O~�� ��Eb�N��$��L#�xw�w�����t���c�22�F�2��< .
�`�<�gĥ��jp>Yt-}�h6��?ҙr��$R;�OS��kD"��ftS�%<o�Ҍ[�hcMl��+}�4�����f�1�\��଒��s_�A�ؚ��ݦ\�T�	�z<����P�3��m	$����E4�l��{�ʞˎ0k��P��ڋj���A���i$H��FsW�3�&�7./�E��&e��P��`ʵp�^�.�����ݫ�x���p{S'�Oj%�.|o� �P�>����?�����J�^	&7B	�$B{'��]z6E�74`��sk_��n���#N����V�&ln�����51y8�̮y-`i;�rܠ|4)���rۧ��C��������v��e�5��B.�6s� �-�M��i=&_�,�g�+����g���l����N���k=x)'B��S���~sT�.��;�B݆6�֨~�Ոl���	��[� ����=�X��Љaf8�?S,*DӓV�ƫ�ѣ��!�4Zy�)�Ƣ������Y�V1����3�\�
�@aN�!k���˗��j���0���> S���hL��u'�M�k�$8V�y?��,Bk��3ˆpN�j����X.��P�d6���v~�;$+�&)rD�4�oU�4�t<��i�?�&�S��j�Mw��3�q_�q\:z;�%鄵*:k�����&\z�}�Tv��G����ڧ��)�;/h�t���?�c<GW�*�C?��UKK@L��&^9�G�?SA^
8d�BяC���2��N��ޞ(.*Rf8�Zl_�>�S6�3nT�  �>5ئ�dR P��,*{Y���EиS|�I}��Z�v!�a�|NC��F�<fJ}�$\K�b�C�ܴ����\���J6Mb���:�*��fӰ�t�kRb"��YAK�x��'���¿���*��iC�- n����NEJsT`%4\�����,9���2�J�>5I�G�Z�r���� Y_.o��K.3�8^��]���f�?i\Nt�*���(K�]hZ>Ra�ēZ��&r��+��h�	����֐���A��=˲7s�ݴ�0�i�>;?.'�_r��X%���1�_O����d�V��$��8�Y>��	Q]j��PW�"�!�W�C��vB��&��ĽOMb�	��o�9�C4
�[��Ki��i������P'r�����~lo��4�W��h�H���؞ۻ2�w�]��!D�b�lz��C3%�ab�?Ȫi����]v�D˺���u]8���|��%f����MB�4�������"���6y��:9��v���J-��ڇ��I�	J����';�Ty-g2��]�ÇٰH�	'�6�h������(���9�#���.�T$�Ocp���u]�g��̈�>}��4����HO��Ŝ�8eT�$�#Tn�}�Rz����^�P��yP0�E��j��5i��%#@���p^�	���F� ���ӌ������֑r�)�Dn���NjmU`�4|��O��B�<H��<��"J 5��g������P*Y����mr�_ho����`�0D5$�V�dw�ww��m���}�E�gEϞm���#ۍ�Y�%�M��)3���?v&�<a"� �����7�Q�y�F��Ï[��*�UT5�Ăֈ3e!�@D
�Q]��=މ��=h���O�K���ی����z�i�Z4S5���f{���W��k�E��wDK_��D���=��o&*�ʳ�&�a�?V~��
p�����ȁi�idˆt�H�+si����¢�A{��؇���%ͣ�cD�;]<��@���g��3�gSO��,D �ґ���?�[D�u�R�ooѢ)���v��It/��Z |㦲:;hyV�n�[��6 ^(�����I�������2��AN���*��fD>v�C��R}<G�	ߜ����� Z5\�����������W�æԗKD&{����|���&���;?d�
��<'�U(���q2py퇙�h�9�0�"�+h3{���^-��<��N�!h)�uQ��"(5�]"�x�	2�4Ğ���,�
L'���a7��f���U7W�[��ҭ�í��!�wA�ΗA�BMС���Xk�F��Dﮛ�6�
)�F���`�F�b��[?��t��ؑ�Y�l$�,T�Ew�r=�.�ԙ�K�E~� PV��ΊV&6o���
&FWf���"��*5eК�[�}�����v"��� ӡ3k�}R��w��e⎐4�|��\�bѳ�����đq�#��'1�:��ҍ����.���B�;&1(m��:Ӡ�����M��~�2U�n����(1�겭�O�}t����l����K��+�%]U�<U�[����ký^��8<��6�ٽuq;��ciG��H�hR_?´/�Be�L%۲�z�9s���=Q����p���ۻb�N��7TW�����H�9�a�O62U��M�ky�����@;���U��]r�^��Im`1
� <}b���2IW,�NhF�4��&��Y�p�L	�yaI����[���{���%��1�9YK#Lqa���;��"f����yt�(����\+�G�5i��*������?Pkq�.���B�cY����*|Lo���2�e��G@e����gF�fj�;K�l��CL~N"򆇖�JR����b���׸�&o�^=�ђ`e�Ol�/R�=񨭦}J�SX�`�n�Ѥ�'���q�X�V���"0���i�AF�T�<�P�^��{��%���Eɞ��I��1�^=�I%/������Xҹ����j��:MQq�l��<9�ʹ>�-D����!Eg�Ʒ5���Z�Xx_��}Ӽ8�|+�� ��%�;V=w��ɧ'b���]O�W"d���S2��q������{#,�X�ڏ�파=���]d�ne���w�"h�E��[����,�����m�8�����ff�����s�u%wc�n~�?�P܁�hMq踼�t�a�(g@rW��9��H3�յ�g�6��ӋJQ�%��'.s۬@��s5��6V�E����̏o�_0�4�����D<���{0A�B�����}F�H�E���! �yq7c�#�]� ��_c�6�;=|���/�S�{7�[U�>X	y�x3�Xԙ��|
is�lzZ$�@g��u���l��{
R��Y��X�
:X�lF�P|ar>��kPı�f�V'� 93�Vx���54���
�sr�c�
��q�d���2M�>L�&?#��V��W��Y���;e�HzCpv&$t`T�<o1��x�@��6���3o�r��B�_�사-�>#=�W&��x+�U9��ݧȨ��"w��L6���
���|*�p�����嘩#���m`�9N�����F���V��B��W��k-x�jt��ZR�B���w����Ѱ(`����� ��r%#ޒx�2Җ)\�V��}ﳦ��_֫���D~��L�;] ��4�<7ʛ�dsO�1�EFz/��f�?�26�ҷ��K}R��I}k����zh�g�>�g0<�0���r����u}�Ŋ��Q"Y|�=�CWX8�;����W��L�WkA�*���B ����"�9tވ�8n�b��ޕq,�z�I|QL��#�x�}��i�Je&99��x}oJX'X�`I�%���vC�=�S/��d�U]���,��uI"���[���/"]+���)^E~�Lp�^�4D�u9K��f#D�B�G�^(WD�e��M�A��%0N<�@����%��;��ۃ�{�)g3ue5�)���OU��k�9�.���u쉏Q����T�ݠgO��0��&Z�)~���u�f\pġ�z�b�h�C�f�+9��!��	k����΁'�M�=��o��7�p��9�Q0Z�����_�M[g��K�4��k<7K�䒠>f�(�1������H&?��֕�=� �,+Y�5�rFW3�n�I�����o��ġn"~�[��R��������$��Rp��:���t~/����0vr��irRi\���|�X;�h�n�ߗ�{������8�i�,Y�N+s��u>��	P��m^�sG�a�s�/�3hz������IS(��z�`n��F�ź�� �J�
��F�4]���p9ddޜ� a<+��P�`3�9:v���,����V6c'AG��FU]�9>d��1���b���5�5�����'��]U��G�?^8d6{�-���c� ���4����Ε�0�r��Sh�L�V]�ͺ�#4zn�+liS��ä\�s�U,�#�K�4̶b�&x����Y 3���K�t����;��]UdPF������1Q��40��;`g�������Z5!�oQH����cE<����e0�Isڮ�Ѳs��m���@"Nϟ�R�m_����xHg�8h*n>b6Z�>ڼ+�9)�����E]�� ��tS�tQ����!��K{��B�񮔤5�Dҁ`��EN�)��NH�+�����~�\����nywC��A��IK�#���c�T��,��������4��3e��V�LiUT�0C�qz秔<�c3���$:��DL��
�h��}5����!�<X$�-Ȍw��.~�֏1��J���j�TeY�x6��o"+�%3'�;4����.�r��k���@bBB�B�� ݦ�{��5�NR߂���0�^��ザ{�Zm�ɊNx8!�?�^�L(jsi�J��E`����MM� d�����.����豔2T��N��~�E��� Д������Z�?��\�-y>o�p���)�h���B���+��v�Jݤ����O�\�����g2��w���*���S2�O1,�tGo%�͚ i��>L��N����Lm�T���ߪ�u���Ut�s.���q�>�������`���4�NP�ص`ڲ����W��A��!�@��Ĉc"�� `^K�w���E,���~��O�.�:%�D�(Q-�����p����<-J8w4�����j~�︺�Ŋ��b*��# �X��Kϸ��X4�|�y8T����,�'��3�}�iC��b!�^�gL��͂?z�c2�/\@N+�";E,B��,B�>T��t�E1���/,�H)�F�h�m4X��X�-��qe2&�4����'���t��5)䉵峒[ʹtFD���{�?μj��qȥ�PRݾ�aH�u��0���1�[0
�;����-W��e�l����jc%Jy��H��	#�[|���W>��0�HT2B�q8p�1�;��V�R�RtSk�G7�[��
�/C0e$�����A�AO�M�[�a�����Bt�kh"c�7jD~���Jbqx?�%ߌ�Hе�ٯAl���A�6� �ͮ�}>t���J��'I�Y�C\�X�x��"(S�Ȱ5��EA貧,ph��Kq�j��H������7��{�����F�T��4*jlD����E�;ȯ���qc�R���	�{��g:Tӗ����,K�Թo����Q��ɛ8���Max}`3���Z;V��RVX��_{���	�s�N�F�Ĩ(�q� ���w`�C�n���c�e>% ��ĕ��l���q�_��*鷸���5W4c���vG�$�|; ��LGy�ٞ�r��z�c��|���C�w��� ��m�_Je�����Re�����Q݌`)!�!PU'J�lL<�8 +(����/r�U�^�[F��վ�A�f������6�O�+���c�(�ɼQ���Œ���f={V��?[�R���-��V$@} �ނ?,&�F�9�I���?+ʥ����]ϏYep��S��Tc+��콞[^GՒ>�3�qW#a̺(�ê{V8t9��G�_���� -�΍��Y~$���v@R��r�\t�NA����C}��g�a6�[�e�k��j54��ccp}Ot��aD�ѩG�U�ꑥn!N�k�g�o��g��B�J��(��:Xb�GF�ByzL��q�:��ϋ���Z�Ŧ]�\W�*Տ;��g���Q����L{*���;:[�
s'�RY�\��I6�p|[���(kh����"��o_`N��<+�z������̬�l;��c������e��:��/V�<Dg3��X�ma��h=jQpe�j\�_���)Z=��������d��hl���,5h��}�b�H�v���ݶ���S۠���cL05�:P�p���5@'㌘�Z��:<��a�9�Y2@��l����G>�?��N+���>=R��ˊp�j)��W�-���\FK������K �|}цe!����T���}7\m_�	���{q����_�k"Ծ�/�Z*��ȃݾe���� ����h�V�����X.\[@#�*<�,SI���n�U���ut���S6+�m�b.E#T5��b��V��;��Ǯ�`�;���`�g(cQv}�h	�63�?s��1Zg��-͹��g�۰�z/��N��y�n���X+��Z��q�_*��\%�����)��*�\������Wba4�ƭM���|���	-�����z�1��P�:c�­����e��S�ų�+�PR1-y��H*��7/v��r�E��g�*X)m(A����-<��Hy,|Qa}FnsrO�/?hhR����}����#~Im�n'�@6)�m.�����HF������*u�@��6�ݟߐ�7�
��I��[�w:���Ϣ�l�����pz)F�,L�I��̘˲J��Z�>dV�ܚ$��x��5�1�tFD�����V�-��˅E�YM�� �����K�J��V|���C�h���Wh�<��[�n!2&�>?S�PǨ�Dn���%b�Grv>u17�#FE� "��k�S)0,�6X%�#�A��x)e8 4����2O���{Կ�!�{ɰ	�����'K�{�@���[���|�CcHC��V��W���Q���Y|	`o��`h�5)��[�KD�=�H4�|k�����6�CSd^�f���H��p�؛Y6�To�;4,�����B�����4��QP��'��F� 4_ť�Kv��>>�-�������EU�Qڌb�� ���[ӿa5�h
Rpw��±��+d^Z �`��t�zi�(�֠N�Zyߋ�F�kcћ�T����� A�9+��i#�@�@��h�-wㅅ�qh?O��a��a�1�C@���.4W�&.���H*=����>N �+��i�V�s��&�\�Q�Br�l�M~zG�"��4�o�d��[�c�t�}i�A��K#b]}�c�jIucn��T�cq0��5����UEG�z��wy8)�:k���%�4z݊�o��dq�vz��Î�6�����W#	�c�Vv���ا�@���ƣ����ƫ���?e����VU���+5=�9�B@2����HN�?'��n�]��f~�/B3+���- :�Q�����Q��Q����/��3?R{Kb�Q�i��r}z�;�n�lw%O)em<�=�Z=�f%u�h9�`!�+&x����,��8����\e�����'n?����8���J�=E���Z�rO�U�_0!������T�ՕV�ĠC����4Ye*@��WjnV�;���CP��J*2�������&�s�+���j����HC�X���@ĥ�� \1S�1���GMK�{��|����F��k�y�Q㳵@o��cn�� {	�����A"z�u�Λ���/�6�T�D�Q�SӔC��|`ΰWŬ2@�a�0����ˑ�X��e�8������ȳ2s���hv��p'	w��0M沌���� �E�hLs5�n�]<���g�h���9�]'%ە�T��F�`k��dJ��0G�Gg� E���6lPУ��4N���,�����DyiGͧ1�gs;��9� �4��K�<���W�+��?pO%��Q��k�q8X��2�[G�t �����V7���[�����7�PI޺�=��n辀�����}gw�)u	���#�gCDX	�K��m;,sC"0x.P�ҠL�����g��͖�6u�Q%���}��ʒi��Y���H5%���B��K�s�-�:}/H��[]ܦT�>ETh�T=�Q�?9���to���*k=���W{�������M>JS�̰gK�'m>gɰ��^;O$!��4+��~���c�.t��Q;�f��\9��.OՆ��A"��E������0��.�~R���.���aV
x)��:_��uB�kKǪ&��M�6
^���OL��3�fw����/�Y�
��^~o��8!�E����0��`>�)���%X�	w���]aM�o<�*�a�G�u�ڄYMt��g��=��͹3���&�9�B}n���+���.�������F���t�y�<������ƪ�p�[ر#m��v�GJ��{l���
���b���OR���A�tz���<��/Y�kF���M��s(|�?�������VW����-�B9�k��hlDń�Z){���޶�5!#%�q@SG���Cl��� L�� ��;�m-��w�8ҴAxO�p� f���}���ز9�j�ed��a���!���J]�Z��f�	������Ų���m҂'�m+�ׯ�ׁ��w�כ[^��(�ֿPH�6���a�!r�p�!zX��rdc󧩽�Ҏ���=��~���P����eR#�m���M�RGF�P��y$�4��S�6:`�B35b�W�2�?lG�*������Z��></v�HA�VʊW#�}P�K��k�$�8�Q�����˘7���鿡���:��Pnm<!uU�cO	i��Q�f�n�H,�#e��H"*���\�g^�P@�=h[��dx6/���	�Kv��`]�.��s�3Q=R]��Gp� ��B㍹��wkѿ8Ơ�PɾX5X�ب�c`3@�e?<�`K�Ct2��P� ���I&��\ڒ���P� �ӻxpO��C�}�jL|!b���Ҋ��r+���Uh� ���9�J�"����˱�gّ��i�F�uoC� LfTjb�!;��>�) !�gu��Iҏ�w ⻣�AA�bQ2`��yW�W��[,��}J!&Dd]��A4���ҷ��l}i�������^��+t�w�~4�򱫪���夘��{ �n�7����a,rxD|�?хT�-�`aԿ���1���$C$E͘M���N�u/�1��"g;VS��*��N�B�e�#Ta�u��j�U���Ƭ!��%{��&R/Y�� �8��O^#�AS�l��G��:"��"&֚�v?�	��jGb�6�<���6����S��i�L�V���ګ���sO�a&�k�pj���Df��'�/��7���&;�qV�����V;�l���&n�_�A/��*M��RR4��:Xv��I1�� �R4�2�VԮN�NQ'�>�ikv��ަ~MGt��	�d��-IO��d�F�y���ϭ���]s��ǀP�Z��L��P"s�ݞ������v[槦=&9 Ӧ�����M�z��Ni�x�%-��򄁢�y�0�����h^�+u��]p��h᥂���6	�ƫVzS+i�HUqbl�w5�#��*h��J�I���l�=����R޶䥣�s�x����x0�/���0����8ӗ��t�i3k�H��*e&��l|�S�$҈-oQЈ~�zY�P�I�J_5��LZ �z�;82S���,�!/��R���q������Ϧ���a�a��R���G��k��{�*��x�X�b#2i%8�"њ�����C"ʌw`N���	�j��^.m�'"�J���%n���(!j9��Į�o��)�S'�\"÷`���9���㭦,k.���[���ʨ����\�2�Y����S��h��@+
^$ەG����:H�����$1y����(���]`�]�P��H(���}[�W������[���IW\z
?����h.k�LC81���WU�al�>G�,�q���6�WZ�	����Զ�'�}El��R`G��B����}��b���KLfk���-$�
�b��ǂ%�)M��T'd�a��h�R
������}j��=,-Z�B�ԧ�ʞ^��F%��^�p}kX�r����;�T���n0^i�oR�Pw�fF��7��K/阖�]cZG����=<������"&��<���+<r�����A��p�;g+ ������i���������ny=}�ɠ��I�����	�d�^��N�AkA�;�b�
N�
k�y����k���!��Њ��ʽo��,�!)j�^>Q!~�Vw�܌}��**?�fY+��8�b<+��|H�mS��d�k��!��b>��&%ဟv��R��X���G"�����6���k��PK�����]	���x�y�d^��O�G�d���uVv�If����,��E�}��?���9Nfl�>ǡj>\ܞ8%Hyϐ��Q���辯�8��C\�S�j`��������+(���{��=1.�{��ܘ�"V�ck�H�6�S3��ms����ċ9Io�Ҙ�[��e=����|�	I�Ob<���y�\�B��z2������f+�մk���Cэ�nz����n&l^x�xp��T�*0Sl쾷n{w�5	i�l���`Ə2BOy�Т�3��暉�~x��Q�������hWP;D (Be���RS�E�gi����D�>&U'[�%@�?:6�\a���{C&�B�H���A����]n�۾r�tC�Q����17���#���ى)�PY��W��_��ȼh�-�,c����j.�����Е}@����K��8V���O�� �|��E�º�ʗ��(��\�������qؓ�3I��Ȼ��~��q�H/����I�#Tz'��=��P&��V�[7c�QբC�N���x5r�9{�)���f�L�9�b��B㧬I�d�!�����GA��'GAO���r�	mZ�%x�ePo��;1J�&���O_����ƄF4GS�����c;�C�7�lO,�����V�7�k�S�Q��IɃ��CD!���֘��y1�z��c����^ѧO�S���B4t�D����?vB��F7�~�����Y�t��-���o{�ev�����$��p~�����~�4��1��_��$S��аS-,j���{�7�T�1ԔU
S��j8&��s�'KF�/C��_��L��H�%mq�b�j�"l!�X����	�m1�a�ddɑ5M�=����}7�,�w��EV�F��*�Lt�v�m[׊rɏ>�a�ͷUo�K?|pb׳��+��6���[' �˂I���@a�0��B_��4@	~}�ڻ���`+ˣ��K	x+��M���'}\��~?t�N�wR��£����N��n+ԝCcq��n�BP�*GqF��cp��#���m��\эJ�+1"�Y����Z����j�`���!8r��6�Q���U� ��9=����`O�-����#mJU�m"����;�$��$�]�ʉ��� �*�c��Ճ8��T�R�˚��u��ˊzArD�&Ϊ>pD�� �-��	����|�i�tR�n�����ʴ�BzZ��	�o1�w�#�Hz�;�Lш���a#�*��?P�ݥp�St����ϟ��?�#\���8�U�|��%��F$�Ta��DD[x�UB�%�,	�=>��5A?�ZOc%��h�N�7�il���D�4F�4��8цo����a����rH�ƊJ�ʜ�R�=�f�lf8A��w��z�o��=���M��I']'��6��T��y��QlJ.�.�s\��֚�)yHg*��}IXƱ*������x�o&�,��Z��:�@��\�V����������^�r�MzǝJ�&`�����rgma�L9M��?3��5�f2�gm�>���@�HH��i�G�5v���C�R027,�X��!�,�+���w憽oR���5��S�=h_8�^ۈ
\�$�l����O�����K��%��77*Y�����ٴp�9�%8�1^�Xx��u�1���c[ձ7��@(Ҙ�Ǝք4������B9��׽/l .�1��D`�zr�e#�d_ఆ>UI(��.^D�N���7��Jk�����B��s�X�Dӯ�;#-�XS�n���v���dP�`�V=@H���2���1ㅞD��ё��9����P���5m�$H��-��ܐ��dϖ��B�0��STɟ���X�F��få��\��t���B3�3%A�� �ѿO��<Z){JD�햳��Ұ�~�%�X���P�qK>[�(͔g��[�
�4��u4�]��ax�Azl?�Q3��U����g����5ה�
5���Y�|>�x�$�y^���?m���'p,w.����*	1��a����o���Ti�]E�ix�GO+0��q��馧��/\���L��]�н�c����A�����;>�p:2s��3��+[��6�gZ�5�[-��8p6���")��CLDN�)��O��S�	�����FF�4�){�_��-�l�\��;/<�[����Fb��V�d��C�J�U�k��4�W��2�H`U�����,|��Ai4���Q0%���s�Yه�F@��m6�#�S��S�m��rPg9
��v�|VL�U��ꢘ,p��x�5��ni�vbT��圢8z�X�'�}۾)�fU��42���^P�v�4��>�k5l7N���YNtԣ�EL�SB5�9��|�PV~@���i��t�-j���w�Y!� �4=����䪨��ז>�U&k��k`M�0�M-�d��`}��K��CJ�I�N���B���|�j��Z�FIm8�~J����"�ဴy��Ջo�:�tg�:��p�a��>q�0_��.�����FP�ŋD�X��}��k?bV&�ek=\5�߱����5� j���>�[<�сu6q�[��N�H������ �����ƪ��z��W>E��8�/Ў����R�+�_�)y8��P��l3~c�qw�B/���q������_Qϥ�A�,�F�>���g��]q8�38�+��<��� ��d���%$!�/ɂy$�������H����[�� �Ɋ���oI ^��
�;�zV��&�e�tr���0	Kk�8(�/U�;�� �ϒ"
z%g[e,Uz�#�R�8�A2w��˜��/RF��!%M-�^M+�"�Fr���n�)�zQ��JNN?ubV��z.8-�=F6-~{%���$�,X��%yyt�Z���Xq�հ�*I~���,6�;�����'�"�i^�-��&G����zP/O�^W=�%M�aq/�����<�, �.�$cB��o�zk�J#�7.�?o-�E������p
��x�0q���&���7�\�؉+���dR�ӻ��vI�M�H/R/�BY��x8a�y3�>?����g8�lP����P2�"�=�D��Uy��0�T�7����9�kn�\򽑽�g��bU ���J����ؗk�&�L�4"�4�~�s�N��x8�'��E�$�����)��GC��ɺ>�2�Σ���t3��n���k}��.��z��0���@I�*���8�5mj%\��U,S
���;�������P�P���6��'����e���s�2l>�G��rE��F�@^�#��^�*`���R�a'�������s��NxM�ƻG�5���3������y�D�Rd=�S"����,���7顒���g�(���l9�fc,�r�v�J����cvha{-��ivҏ�����+£��|��6;��47�^0G��Ym����@�p�rp��A�w!�"@,�N&���j���Wo��;.c[s�P�MOP	�=���5\t��ڦ"`+94x�	0{�n,@<�.:���y����K�`ŜQ�� ���������8<کj���\uK�2����P�{�\��_�!ߌ��rZ���+��;h�f���뉀VLB�T�A���R�jn�1�QџQ����{ *�^���`5c�;Gp��/H	��`M�0^}"�wV�2z��D����&>Q�g�fMٗLEo��x�Vej�	6.�x1�]����~�Ȇ��C x�(rAk8"J��	:䳗�B�`Z���/A7�a:Z�I��R�xh+\N�,3�:�e���.,v�I���R�bP�c��W$vYAf*�	<y��@�&�q�@&x���x��:Ep)�Ŝ=*��xu��%'��xj�.O=)���iW��+/�.m�����3'���*�f��>�N�p�Węų�����U:����e�x�d�O��7No G�!ܘB�]���9M~&�?��)0Z��\��$��G��Z����q�Qb@�7�Ex�Z�Ho�p07�G�j D����N>��Cz�a|5|�R��)�aղ$�k����p�UIK�h��$+FF���t�ȕ�Z�^��F���6V��8�lV%b�<.�9ז�/7��C豴J�2B�4a+(�H�[�У�Y��T�h�w��ED"�]:�_���X�� �g�л����}z�7���]]8�Ե^���H���&o4������/�	Wm�^��K=�dڞ&+%�}�T�⋟���)���^�b��F�\̢$�'���)����y��6^���%���M��޸��f;#ա�m��� ��Y:�-�=�g�s������bs*\_>e��ԝh�ИZb�wbܰ�+��XƆU4�G��Ac��l���$9���Q��RhЎ��S���7ea�K޲��F��$'be��!�ť%��_�����i	��[�4���Y>���L"�.�n]�5�<Hh�j�XOW�LΥ�*,���mh��{9��lMz��z�
m�[Vn!<�&��R�U��×P<��a�����L�}���z@�4��K�I�0"�gF�U0�Ӫ�4ݶ�kWh��|d��� ��"p���c����0���Jb�Ia�C�g����c(�W_"��7X�S/�+ʜ�Zr�RZ�r ��" ���J3{?��#�Z
s�1�� ��c��X���� ���%h��tI�A�j���,�s8x8#E�\L'�,A��iv!٨;X��7]:1haN�c� ڀ��-~��sD��Y��� ��ۮp��x�Į��EQbΖ(2���_��ݤ[[�;�QFa+I�̏Y��A�<�����H5A��bΔZ��Qs �Hd�0	f�.��m���4j���$Ofr�#�'#�b���h'���Z�b�E<.{�Xj��j䃇%)���U��=�G��~;�t�
��� ������ŜAaQ@��!�>.=x����b��b>� �ɍ�2�׌��d�o���_�5S�lQ�%�[���M��ɓ�YR�@��ĵ���S��	���!�6)�y�}�mt7'#���<uWY����f>J��&�?�Ky�����]]��H��� ��.!��y�E��Qۅǘ���c���XM�O�s����:�R2$���l��z'p}�Q[������9��e>|����Wˠ�P��P��M��/n�)�ʅ���c'R�	+h4uF��c�w�\dR^l���0 -��܁ujY-�%��uUrjh�q�SKPvnq$`��Ix]���5p�єf.Z�b^ 0��`ov��H�����Ed�dhD�B"RN	���?�#��I���@�w�� `�\�/�,�e��/�r�&��S�[�>�m�j��-�+��7{���@���:��� �4�K2���p:|�xB�Pb�����ĊFfqȃ�Ox@W3ȴ�D��N�0�5��T�'�6.�sşߙ"�/��Nǯ+��N.WR*\�7.�bb�G�$I����L�6�:�cV�8�X�����ǽ��?��Ty#�>�A�60|�X���Mň,Z��@�����`���P���V��D�sJ�@eB@$q���HJ	݁���y�?y͂g���n� �l���j�yk��
�~W���\�)nYr�G�B�Wg���$�1��u���m|;^,�� �,��"���#�n0T��A4G�<j���	������7eF��$�^��I��RI%���^��F�r�N��6��Z�l#���j+��s�"�u�B�E��I����2�D�Gnc�G>ε����v,b�Vb����&�\,�CZdP�I2��;�P��y�Z�ǹ <o���v��I2�n@ ��	�	s�H���`���{%�Bi������d�+��ݏ���-� 7����$��q����翤!P��a����A_��h�W�j3�z6T�е��{����p��=�/XQ# zp�5�����f��=a���`��rap>�X�F�QU��D%�-�D�W�9ʈ<�׶�ȩ�n
S�����&��[.��`6V��EV�a�:}q�Y�;E��ܠ�X �O�N�%l{<�j&>K8hC��0�P�E�>e��Z��PrGM�g̚�v�)miW81L�h�K�ǚ�G����Q6q����
s�0�
�;�3j~=sd�z��ڠz�k^!<�m���_�+��1����6�s#��	�
Bl��[5߷����0�?=�1J�HÛd��};��u���]����V`�Դgy��Wd�ߦn{��M6��]y4z7�IT?���@<`�7P�985M1������y�C�	� ��}�A|:J�b�J4��D䭯�֎)�u������ ���*i���U���LJ (H��b0*nUPe%��+�\��