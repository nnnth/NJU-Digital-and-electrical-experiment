��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�E3�hoA�zFҿT���8BD���!O��<�n�eg~��gI$.X:Z�ԉ�Wr����}�� 9`��K�f>�!:�9�!Pe#fpc�������v���҃maO���bm 3��c�b�H).|/�6�N,΁��f�[ x����c|_��Op]�c��B�G��-�M��u��B�ŭ?��w2O��W�0�N���p�°�t4.��X*ŭ�)�RH�D�{2��ՠfl8��x�x[siKݹ����WQ5�I��NK�p@�'6�Ϳ�uͷh�o�CL�� ��<>�e/�#it�$�F�(������
<..��I*�  �-k��O�wfqP@Lc��<B��JU��d���o�V�i+��Ʒ��v��o|��{����j8��9(�j"�ʐ�OB�s���7u[BN�MgQ�@Z�����W?�!��ګ���o���{Z-�8$f�H���y܂�b���2�b��L��v\�+�5�Š��c�D��Gda��]Հ�a�]k�p��E�7���pd�R��{��t�P^�sسd0�2,���п���w�^��` �¤��7���Z<�Θv��{8���Rb��"�M[�G��vy�)�g2dH��+V���Q@��ٿ��_js����L�k;P<�_:V(�H��_�p%Z��r�]�э���:�$/Mt���Iq6dG[�v2�+S��E���F`�	�@5��<DZ�R�ݼ�9T[��������D.M��$:����Fc,�c�b\=�㴁[�e�Fo�|[v�	��D����l�)�2F�F�9�X� ]=�0��A�55�v���ҟ[�D�� J�����g�	Q)�Z��>�ꧾ���6�2�L��<Jy�H"�vJ~p�b�>�W��0�f�l�p6�"�����^�U^_����fW��=B�`��#2�ex�R���^B��TdH�O�!O��	��zv�0l�Ҋ����8a� �_/��ur8�M��X��N���Ll�x��FP�8�ʨ�ʸB!�M1���b�h����]	����	l*�{���I\r�/�&T��}����c�����C�y���(ϸ�ed`Մ��-D��͹7+�/�
(�L`��7N7N�uܸ��+ۚj\��ߡ�B�%ϥe��Pm�����s�T�R%6Ę�|��M���_PX��\[���M���L�=��+���[')���zm�b}ɢm7���|�1�,�^Ip�Ι��TX%/���+�s����#�f6��f��ڎ�^�O��oEWa	Ae�tL�/���?5wޘ���0�ZD<F��e@���N����Lø�	�6,��1���?x�h)�����:��t��H�O�� ��Z�$)X ��)��.���/�h'A����};� 3��&�]vN���#�n��E�
g���aj����PH@p�1�r�z<~y�[�&��D~�j'˥ƷU��=�:@�ܨe	kM��@'4�뻛�(?!l(�%WgwriQ2:�8ʬ���!�8�FI7�¶�ѭ�*��zOGHhik*߼��/�/԰zx0�2�������x��Ťz�u�>.��$Tq�Ѽ+�*v��v��IN�dK� T���޽�H�>������)�"�w�<��Y���^�=2��Q�NxPd�䑾�&��Oh��"�į,�&-	Egp_�މ/Z��*����T8�
B�I̜юv����y�\���`��{q������P�7�s�G;�]���[�����![̬n	�{W0#���N K{Ǉ75Q�����N�CΎ�0��S�4���&�����w6�'v�j��Z�j��=����f���	��Vi��ip��.����mK��}ĝ���=?N8n�w�wda�@ƶ~YN�8��g�����a2B��2��w��f]sO4Z��8 �k�q�/ ��i32�G5���Iñb�d�||�U �l�u�)ٞ�)0MZ�/�eKl��̱u�c�$0.nC'~�crdI��8���ٞ�/��b^�L�GxXF�ѻD��*��C���ĘmBS.���J孆���ч�wn��7Թ������X_��͹Jd�k��TG�DZO��v�d�6�������Cl+Yw�ǃ�K[�T�!)��9�ܝ��c�n��a�ɥ�������Iq)�[�)��$&�۷Z},�*=!���At3��n��x���b��V�~�\�͡�x�]��N�o?˔�%ʞ%�|&� �A�ۥ���˸��d��ޣvZ��*5��G4�a���l 4�h�L[����ˬ�`�%��y0��u�9�1�[i}|{�MLP�ζ�U��M����=���R)�X���[��D�ۅX�j��|-o��'8�۫g��rZ5|�����i�>���)�,�D` ��(\-bs�ۣ�� 4R�i^'��p�Sg�6A[����*%�~8�,��'�}nJ�
s���:׋�l���&��Ly�	���s�m�Id���I��/����x�7E���<l���'�2/�nR�/u|�2�*Y+������x�ܥ�f�w"s���Pj1�⠆��؁�B��YJ�x9��=H�x nH�4"o\��r��0�ޭd�r�un"_`��A�u~����S�UDb��^I?e���w�����{���ٓ�4������P,V�^���x��J��L\F��C�n�����;�����^����!�}Q�ed����i��N�n����'X�{�ҋ��2^��B���^xU#��2�' '��{*���|׬+E����,�l܉�R�C�ݷ	8Dۇ� 	=p���e�֍�[T��k�Oʰ�:�Ih�Kw*U��~?b���П&r?J�R(������-	���*�	R�i���$ߎ�~�'�v�V�'rq������}F	n�zB��nF�4��DktqΥj�������̾D4����|�a�~,�W��#~�$�R>���{̌+ﺆ����7��ߋ�L�ʑ���2�����JV� ���i8�04 ;i�5?�ޯOXr~�ɹ@7ы�y���"2��'U��\GhG��{b�ɰ2��0�;Z�@PB��G���6c�bF�إ��^2��o@��F�����1�'l�<��L��*y�.e��"�"Ey�#���9�
�<��t�+.H(x������3��UJ�Uh �)�� :�����J�[�%#R������}'5�'�H9�t�죍y�'l
�xټ��ܚ}�hI��۹��;'o�4L�r*b1����*��m��9����E�4SaP�� �}�����SkX(�_Z<�d���u�kx�ve4���
F$o��.��n[6▿�1v`3U��W����Jp��1��i2B����. `I�\~�4Z���A�3�M�u�Q��5o���1oR]��7&=���<n�C�� a���X�A���8��]�k�?>�p����2�/�������ʚ�-�J^���O�yN(Vrp�\�>	3A�jY�_3��n�cOm*NAa[�H�g��f_�2RCk�!Rp����Wu�Z�!�|�!�L�yM���p�mƚ�[�~;;!c���LV��J&0Z~���
 �=��o~�����_j!��+�L����?�DD�,<�Mk�g�ӻg�ܩ��o�}�/ &��9�Z.E0���ca�r*QHh
�L$(��)i.���Co�l��t闋]�le����˿�i������}2��}�\��O�s�f�}�!������m��c�=f!|E�j�n1��,�K���|wFM��XL��bYY����~L��wǎQ�ʌ��h�R��w���^��ʝOH%P̬�CJ���P�AO2���y�ɿbGK�I`����n=WS:D��0��8=��R�%�6�=��SGx��B��Z\!�O�J�+P2�����̀+�ڦG��@x��ܶ��~��FǵE{)Df��P��/�_.�)ȋD��<Hk��\���n`���{ކ�nQ�$T:66�a'�О��u�"ՇB��;z��� $��k�tJ$9\���vV��E���\�?��^=@"�'�q�WFH1l@���B{g��P����b>��ڏ�tѱ<nO��A��� G=f�oB
��6�U8��JD��{,�$J�0Zѯ�7��Ksa�|���ٹ�Q@\t�BokR ��G+����W�Sru_��N���ݪ/�K��>�?�00k�x���م��l1?��ʊQz�E��ť�����Po���V*LX1��=��ͱ�ճ���Y��ש0`��&K:-"�z�.��Wl��q"�5h�0�(p�O���f-SS,��c�����bܖ���62�~'�QM�:�W�g}�����3!�j٬㞭���D	Q�=�H�vDVCFPnW��oZ�4��A�G2vi{�B���	rg�r0�Q��6؏5�n�%"�'<�)��>l1���>�<%�Y��7�Yd-��5��{H���L�G�m� ��y�vX� �a�B��W5ĭ��K%0���QJ'8�Sz��D�շ���%�@�@Ў��A�ڐ<���u�j������:��K��U3�>Ѭ��;�b=~r,�������4���6�?����ؐta9`!�!Uʎ�pJ��bp�/w]����?�y�'4�N1 ��bMֱ�v?�z��M��a7��2���Aܳ��b����r�3?�3�ǅY�A�b����Io��YMٵ$�\��t��tR���*�,h�a���=G�+jo��@�����g���א�J��WؑD������1����/`/rd��57�{�9�a��p�5�����p�ԙ��E\Z�{����~H�#����0�ѧ�h��5_@�ɝԞ�˟��`XrTB�@e���[�sZ
q����eZX�X�t�WkI�4����v�2��փ��>�4@�r��,��ó�%Iլ�9��8<K�������(�.t$�����$��������Y��yQ�=�i�%5�5����.��
��]���C��;/"�"�e2~�{��R���`�y[�\$�h")���m�m�9#^���@�D|��Sk؁�*c3�P��"�;)�+N���#�>�s(�Y!�EN6�w��.5��We�� ��϶c������ǼE�E��H-y��V	O�s��/���MG�*�>q���XN���ܖ ��dn�/��N�����l��#j
`�g��-���X<@>v9�/g@~��/ө�J���>�YV>�� '�r��dk��I�V;�X�>��s��D��1��+�ֻ�&L69�ط4�(���=�,{ɭ���%�<; ���Q�X�Ԟ�1J���!n�v_�;��� hl�b��䭾yxM����VZL#�W�Ÿ�s��<�x���	�MrW��f`#m���Hs��]px���WE,�M2�0���̱C��Ҝ��(?����LC!�d������7Q,A:@��o.T&	��c}W���D7w��Q:Wv$��E&���$aG��$�Q�q��I2�l���s�&q��L��ܦ4��w�K���px���㿒���] xva��t�KU#(�,e�+'�S.@q8XKP��~@��$f85�E �F��Kb&wH;���<�a�z�����
�g�mn�cؼ�['�B����x�k@����H�\�\���kf���c+�I˜Hvf��hvbB�.#�d�9�}\"�M����k��dM`iz�'vJ����@���(�l�D|ݮ����l]�0���'���J���F(h�j(�o�* $Aɓ�i>g�}���WГԕ�_�ko���b��Fn�VU��9Y/���#� ��7�"b��)��4UC����� �����]70L�Ҷ3�Q���b�>��C{4ᄴ����e��7Ȩ�G5)�ܠ����ŕ%`�/
�B7�kt؆�lj{���qҟ���w�G�?�*�$V�����y��!�/a�p�h͐l�>;���}�l��j��ML�u������M�|(�*%����B���@�~1߶��A&d�	JL��l��ҞUg���b���lU�mz~�R�S�T_������/��nDڥ����*y��5�0�A�qN�NV5+
��l?�8�?ӿ��A���[����d��2�w�!���kL�|���܆q��v/�wUez�w��ɏTE��6��L�MG�PΩ�D}�]�ӟ}�S���gwx�{ᆔB�1x�[Y&�T�tG�;�AX�*�N����	L8}p�����&-W��%4Pm�'����~�����&O�pf���R[�P��n�oWښ�阭c܅�0�6ti\�UB' 1�[��N��������x�����Z@���iȋ0���(��`z���@�-Ǌ��2��Vˌ��Բzy��pM��|��>��ʈ�M"��g�|�L+��J�F竿i�?�n	��k���D�:��*F�o�1=;���1��ڶqE�Y���|���zJ!A'O�[vꏣ�" �W�E5�N͝L�|�]��90����T���3Нgطu������	��x�X������Xlp�� �z��n�!�6\�-\5�ڶEN�E)cg����mt1v �Ù��%��_�`�gy&���1cQ[5�b�>���k���L���^`Q����m �*�K�tt7�	�,��US�[7|�s5Y�}M����$�����1ت��G�����e�((�/CƴwQ��EW�	����j���hy\B�bg�Q�T��c��e��-��st�TD5aK�a�����4y=����R i�����T�=�Ұ�=7P6t\���6����q�Os53��v��ȶ���|���=��r��
�����Bg��*[�n��ȵ��F�4��_9�G_tW����	O�1#�B�Aw����0yz`��� W�X}�I�	�����p��ђ�u��#�lA��p����7�h^�d��Lj���˃@���8d�L�p��">�7�bYT{./@ײ������钙����F�4����t�(G�xh�]���fVM!Ayz�_�s;�����5�A���#��p��Ñ{�e�n�_�td��83����1�~�����o7���N�w�����0q1��	�x|��,v�]�J��K܍%:5�g��+&!�� F?�#�It��m�=���B'a�*�>��"�&�қ0��HjB���������\�n��dzFv��i��ɨe,��!T���	d���v��n�>4Z�l�gJ���Tj����<VVκ��%	�zb�[E:��4ĂD��w�g�������egExyc�*;�	�d!ˍG@���:�hK�q��f�筻�M�ŧ�%\}��b)�ư�T)�C�D»ǌ����ة6p��J���È
?�FA5.��P���F�B������3B�{���\H����;�:+7x2a��sG-�_�vk��������W��i/������ k��������:�_&�6��!���<�%ˏ%A��'��tO������[�����3����T�)�|�鮆F�U�rp��\=J�ڏtn�)P���
W�����n�fҫ����!�&[R��~�Ss�@x4B�VCŔM�`��z��ZQ�Wl	�G<4�R�8��s��h(#!�o��o��=�?��s�����+y�L>����<@I�al�?������YgP:�i�F�q��X��.���}0�%�_�-�?�E�-����
Zam�L�NC+×'~�;���۳f�DyƂ~,���7Ө�$�s�1m 
��n߫m�m��qo�5�	p&8)��CK�vp��jg�s~��G�������R��9�������[�rʿ����'u��0&�{�q͡��"���� ��[��$ʲ��E�	Zn�Zȁ|F4�E�F6�$�_�9{!ޕ�z����}�P���Ίai"��_꯫:�Q^���̬�Y����c��we����hK���b���n���Ioŀ~�cJe��6n��?��&���̷���\D8xg�W�djB�H�x�����=������#�]�������y���wˢ��eJY���:3��%4ڑ<��6`�k���|_a�.夎��	�p�����]ᯍ����Iu�m��q�7'�H(6(EC���L��_t�-A�Һ'�[8ʆG�8�T�v�s��Ч
ݫP��+f\@&%�T�5[g��9 dgiT��=$	<�
�G���T�R��U�B��}�P�$��3
���Q��J[Gۥ)��o�ꅶ�ž�	T��W�#/���rd�)����]v���89����ىkE�w���՗B<P>
�
�б�U��um�7�F͎���H�*7Jٹٖ�>��1���4r�Mݴ�U6�c�"��5���t'h��P-^�a+4'1Ss�5>�o�����9��y�jG�y�N7�X4',xF2F��n�	��}|�������SK�;-\N$C!a��I]��8F+P���LOt`�r�]��3��)8����i��t��0�Cnĳ����!fD%	|E�R��:J�|��UOT:��TI�� B��U��4��Wm������4|!��\�|�o��#���ɦ/*BR��h�Nc>#���;Z����2�]��&&m�*3���_V���ZO��B2�v�����h�d���?T��0����4�?j)z���|����	����}�P�� -� �J��������8�(���I�;	�
+��:РD!��}�ʱW�2ۄq��P7
�.��Y��c�Dp�B�g|����g���f�Xz�j��iZ4�"�ok�L��e�r�;�77N���8��pi�o����$cɩش"b!M�t>�S�$�Ԁ[r�>� �L8���qRR2�����~M0�ܪ5V�Y٥'FA�7}�3~V�ڵY0��/Vo�s��
ϩ��Gw�T�bi0���Xy�f�97�Q:H�p2�ܝ���,����٤�y~|��� w.�#�D�{�D�0�M~�=Xg�mu��mщ���4E'+$H����JMw�c_,����V~�|�=Q3|��k�ܭ�H4['�ohN��Fq��â�	�s����-^s�⵲���頮�H��o��|;?�����B�ܬFc��90�"�Rͮ����)z��󔜧��*^��O�Q�����'NE��}��,)����3������iH6��~h�c^L���[���lz]�,:�s��n�H��2�����W/����{����&ohk����5���n��V�c~�&ɽ?z�4v��2~���e/���!�_��n���p`���)D�)t͏��;��Q�>0c��gg��'��������\�>P۾� q&�q�H�>@���8/f���$���@���2�Ђ���FȍD�/��{��;�Ͼ\�k4��Yvc��>@�\a������Ȼ�8���:X�5[�+_Q�\��QG}�"a~� �<+a�	eZ�)��i?��m�a,��6h� ����2�R�/�Ɏ���H�#��	������^kȂ���Y���3��ؤ�� ��cڧo౷x�wƚH����H��s4�����~?�
Mn�S�5d�TeW:�6����x�B��U�1:!�P��DE����~��+�Y�t�ҋ]����<f�����ƎgI��#�%!���P`�h#4]��kt�s�N\�������G:K�������X��m[�%�-���^�v�j8'fj0�'�B�b`:q��4�7�a�ԍh�����`qe��N�W��	ɭE�SVeaW�#�Ò?0EӖ#Il	��(� ��e�Q�(�{B����I���K�,���X<z�W��[�I�*���o����\<�آ. ���A��gܧ��L��j(ݛX���N�~��~����~ȝ��o��Q���Sp0\ɓ%I��'&0�X���T�?r�U��S�2Z��B�s�' ���&t��D�!���<f���>��M���qЏ|֮���(��;�OF>�W��e���^�GE�D7�������	ʡnk�7�_�Aa:����EK�	3y���9,sUǬR9������#֕S���w�ؒIp+џ�VB���eB�M�����Ȕ��G%�F�J�n���8�I�	�5�rEb����]U��ژ�Ӷ-�$x�hVv�$�Dj�b� ۵;nu#J�-��yq�%͠\�s��bQ�NE����JC�+L^ʣ̶����8���12B9��U�ɖ޼gz3�kv
˸����Z�\����v�k��(Ւ93J�L�l���e�|���W?�ɺP7Й�T����*0��\�b��m�X��Y���c�N����KSw����#
yYvlS�E�$��CP�m�6���<+�[���Ƃ}�7u�l@ ��:�}�'��hXD�z7z��=XC��UO�SX�����'�TrG�i�a��c^�n���߁Мҹ<�j�H�Җo9��$��"Wol��[�}��\�f�Pyo���/����m��cm�H��D��[�D�o
x6�0&eD�c�V����|�� ߒ���"���߳n�]�bJ r!����ܫS�G��$�8_�@ٓf��Z?:[2(w���Ø��m������tn�s�H>>T!`3�&��T4�s�
\>x;ş��fV�Ŝ�~ӳ�$d�zQ�Aq��=�!�e:=r���(sqJ�i����+FbQ�l�Ρ�����h:ua��jH����f�#� ����d�M`h�Xʅ���TUҭpUf���t�T�(�|`F������v��/��A��9^nh���-��X�>��>�{����/LB�����U��L��X�O��&��/��_v�(*p$_ �~g��}�49<�V���w8�������/�9X:� 0�q^���U��VOf���<���3��������
5�%Υ䳾�ȴȗm�aj����_�����8E1`�
���nR����V8�\˒y*��ROޕ�+W4l�����KB�(W�����q��I�p� �M��-�c��&\}^�Q�>!%m<@��:LB5Z�~,�U�?,_�{��<,��on�햇�{���,����(�ď�b�æ�)�X��M`z-�'����$��� =����x��^s�'
Fjm��O�����~��'�`ɔ��P)_3V�c�a����6ڢ�!}��h�+v�}�-��wr�h8�ӆ<H��R�Aǽz���\@����2*��d��eG T}�����?w�p�ҏhg�R|*��`�R3$����'~�g3ao�U�I��&��'��N%=�����Z��m�F��e�G��4���9�*D@.C)`�t�(�sg���z�N���p��<�ye�7.���Z
�q�8ӡݚ+{�"�j疕��ǕQ���C�S���Ӳ͒sf�,�>�YvV�Soȵ��x�~|:�r���pQ���!R��@���.$���@�Xng���=w`����N����1Ov/����}�o��(])�C`�8W!�:����&��X�O�T�@霅�B�6]WW�U���(23�6q"+~�K�
�g�+��14w�ha�ܘw-��]o׮R~�f~%8>X$�,��q���Mx(��HTS���X����w�J�Z"0T}$�`�L��qR=4*�� A�D�**j�3�Yض�~?K"�u�����t�o�Y�����^�8>��t�K�
�[�Z7����E�S����c�l��[�;�w���C:b��H >_�_t��:=��|�],�PJn�Tf�q��O�����x&����-A��������+޽F{0��VC�R�T�7ߎn�YL�/%]K�����Cm�LG�C����ۺ�p��"j��t B�&H���s���=�{�>�9L�"hW�m9�BF��?
*@K��J?O����r�.�tS�,�tX�"����������7ų�&͋���,Y�S؃"���Oj���I�C��YK�n{]r�rw�����|F�Br/��A]3�jBxJG���?��Q����%���Wy�`?~�%Qu�ނ��m� B����n@��h�-�S�3vMT˔Q� �P����G�۪�G;��,y�6����u�J�p��XsF�M���H3Fy�����/&`D�H�\��f�@F����/�PW�hX�MC+Q%���Z�_�?Rb�Av��
b;I�Oގ���Ϝ�2�:� �l����>�G���PCv�������&[�U������:�O����L� K}̬K��H��O�x���h���Y]�]�2z�v@:���RO�U��P顐������؝&�)ީ��B���0�{��vi�y���,o��g�GTh�����N�oj+{��U���m߲G������&Kd�\4��L��7�F�4�KK�t�.��0�{��V�1��������������u��G���(:�R��e�I���(2�+ z4Z�3���JAoR����()
���M����z4o��>��!	 PՈeͪ��J�h�>_˸��f9M'��u�3"s8d���W ir~c�'H�>�L�Y%�; a�U��n���@[~���g�m��B=��<H ��&9�R���W��2�B����p_=L�G��6����Y�xrv�@��Z?�?�3�Е���j��r{==�s�m4	)�:z����X��Wzf�A:�oO� 4һʷ�Pg���P<��ΑѲ2��� �V5����e�쿼&����#��`n>�Gɦ]�G#�:dA��D8�EL���
WԞ�nC_�4K���"QA枫�A����qD�u��n]�A��j�d�X���9xu�������yS�ZW;0�sf:���V��ff-�\���1D޿
s�<�`㕼\|�s��p!��Ԗ����z[0[����@��A��L�$�|�4lY�W�f�@֋�~�H?���k�C��� ��r������ҧ"+][.Ԭ:����o��IIO�}��)��������b~�6$	�WV̀~U>���?F%�p��n���)������H� ��I:�=��=Ofla�D�e%�.�攢�2��-k������RƠ>��)�sj�<Iw}F����#fb�~&L}��d�-WP���G�ĳK�F�ˋ�j�Q�sB��wS����M2�<,�-��N�4Kv�W,d��ˎ�n����(r���]j�게�+��\�Xu<�J����I�] o'�qo�P����'6f�<�'+<8:q��S�Ⱥ�q��',vd��%�-G�ha?����@���Eo��u�`��w����z����i�7-X�q!���z�,�T_1���ø��\��������9m�^)��l��:L�\�kZ��$IQc����kDwp�F���6ӉVFn�Ȝ�����OP����������ȑǹ~���ʽ�1*0=��VP�ӝ�U�G�P��ȟyw�B.s�8�#�kub5�)�(J�"]��E@�U�0�������T��9��r`�5�|�$=N��x7y�}�O}�h/����.�ʅ�=��g�<g��U��wFc�p\�
]���C�V�N�~�U�����a�c�:w��9�:N�i��x�4R�|�N86�E��ox�����RQ��&m�V���e�����ś�d��ʫ]�V���PT�t)���s�R.t�k��@C��c�B���#w	�aÆ��|���ga��<�7b�'V�"������Ԑ�}�	zzκN.7�CoKy���HY��}0�[�?���P]�vE\;�K9�FQ1��i�M֏s8�Y�h�ѡ] Ej��H`����4�3�*�@nQ�p�4�R�z^�x@�4��F�fAq[���\�`�s4�	^7���2�	��� .�9���pA��_KJ侔����Ā1æ�}���m�@~U������i3�P�KL��4}[]��Г��%�o�#C)�d����d�Id拼�-Y�|0�?k��'��X���Q���j��.�&�w�Ů������w���4�^����C�]��B���	�$'�
!�g_|4}��+��.�Mċ���+�!��1ɍ6�,[�ɐ=^�˼r�5/�|�ӽ�Ca�fa(ͦ,淆�sV�[�X^l�Y�W�1ZJ���̮�xh�Q������a�3�6�x���/���Z]��݇����ƛciw�&��]Gg����AA�\I�q���a�����"���1�L��Р��@Я�.�n�7���Y�Z�Rz�7�����%7���:�-)�G��y/Z����b�ͼeL��M,v��]�5��uV�o�j�����:lb�);P_����5͌�҈���û�ͺ��t��z�IL�6}/'�h�xq��T����"�Z�}��MB���9Ge��D6�ل��!0�ּ�%��{�xG2X�d����wi����ڝ��h�����*k�ؿ��́�E6�?ߟ%�y���hz�ֆ�M���~�_�y��������_���נb"�/� ��rI�7A��y�E���b�5;0W���<��I��V �j��X=%����6Xf��~߬>�h�2L����Ge���j8{OЭG�O�BY�����y���� ��b���(��������O��⹪=ױJGtkv��S�I�b����Ó�ٙ�2qK�z����K�t��� � �`�"q���m'O*��Et<��3b-�[Ί�f0a��l�k�/���$͊���V�-�0�������&���2�I�5�mI�^U9��|�i9������V�{t;����zN�����|e4�����ھ��+y��4,t
�Ę�*���{�����c��������}���|�f�����������8�)�b�!�A�/$�Tz��*f�xܿs5����������C��Lg�\D𮱑�}�y|3�uߥ�1~�����b�1�� [/�~��b�T��������)�=��l+�j�kl}���%�ӵ�K��Š�y)�pb�:%�Y�E٢�!_B�l�H���Ia���Ww4�*J𾁃�Ö~�nV5k�&��=H*/
e�`��_'��N�5�Y�RQse�cS�U�MV�F�$L2Ws��4N��-���ߛ�+Ȝ}lw�ĝ���7GJ���?���{l7G�#��jw�"���9A���"A~*i�g.��F��Cy'2��[��u����
�|;��  ���{1���"�;�}V���e�G�G+�tn`}��Ι�{^�>Β��M�x��di��D�X�i�d�S�F����o+/�!�o
�-����,°$�
�<�������]����(˹u�T���q-(l4�J���pdפ��0c*b��Ύ,#��ee���=��~t�MR�]�'�e�:�r�}nm�|�~Ďq���I��o/�7'=i��ӌ�բ���lz�P�4�=K������o�'Bkd��0�R��㬠�qi_�'�>����T+ښg�T�~�D&��Yl2s��s�O*�N�͇)R}}��c���8M��BY*I�/�EE�Xg��Z��im��(�y�ˇ^K��	�f٭�"f��V�g���m�O��qf��iO��������_���#|V��q�PZ���j.���(I��S5Z��Y��X��6�H�޼�ɩ�+ �`6�X�	=�!??[���(p�=����-�2Q=��8DH��Ȋ9�\��;��%d�7&h�6����h�^�p�_�������>��B3�8z��u���V���q���CD��$7��#J��;��!�8�!F�D
4 �e���:`�mt�[K�#"j���gR�^
W@�X���	��m��
Т&hLEZϸ��6E���,0�������1�"��z��N�Ŕ4������dѭ��e�yy�@�r�4���Y�L���o��d��A�:�B0�3������_ �-,���>@��Ւ���Z���J1�g�[0�z�f�hl��E���G�a�s;b�Jƻ\�����,���˃���+Ia�Q��[9�,?��V���	͍Y�;��6���k�m)��Z��P�o�%��ۢ�7hkmĖ�AM�,��؜�c�>��]O4q|�v�P}��e��@��n�)��-vl�Q�)����w����i<f^ ��6q)T?�T�B��ܵaL�&V��%/�n�d9��a��˭;�z7��حR�kk좴�}(���4��̻��F���Ÿ�.���b 齢;�I���ݡ��'� �� 2�q��N������%����ҠXI��L۳Kaa�ȦN�`f�����,>��L�#J)���%�� ٖ��D��I�"Ex�A`�%�3��������\2X-L~)Nme��sdE���@��W�L�մo#����X>���?��m�p��ipX�N�*㕎b��&��I��Vm�ݫb�b�A.n�q�أ@�q]JW�L	��Ŭ"����o�������ŇV�h*򿔾�샛�{�L�_���ׁ�PD �=R�Q�q0�^7S���>!�����u�5 u6b��|�KG�"��>�!�:�����f��pO�:Ҍ��r!�qlX>��9?|i�=��2ɤ�����:l�9HTO���;���f��]�kz�|�d&F�x�@]A���E�f{M�\0҂Eq��v���\,�3@�����Y���8���y��1�p�/ɺ�]��o��mJ_�p�(E��s2���DܡT�E�!�3$(.&Y�K�v{&�A��+MU�����.`k<����G�~UM�qpL4�]u��fxLL������c��'p�WV�
U��/�uk�ڜm�P��\6�m��?���hj�Lԣ0�p��C�e���v�"��ϼ�].\.�?Jߔ�Q�KbTl�c��d�f�2<�W埘\G����fj=���Sbו�W��X*�b��AM�-r-"o 
�B����F��?���܆Ƕ���O�Ex=����lI3�r�����1������vG�,�s�������	����ѣ�rxQ�z�H�NV�PI%�c��e g��9�j>��9��\�Ϫ���7�	�8����](�?����ϥ�����`-�Ϗ�y��#Cv�K5I�e�s��
���1͊+[������;p�����
��2�;Fk�P^p|S&�������˃�i;"�e��iu�{\�5��%F�+Y��4�/2o�������d�U�F�k�=
�;}��+u�O<�z^�P��1���Jt�z�!�8|�$�Xf�(|ɹ,Ó��[!��d�Z#0��W�����:M��^�H���*���A��h�v���#`+a����>�s_e��@ö�:	[AP�ƀ��� ����446�f�c��aSB� %s�W��k!>�8�KD�Flm�5z:�?����`5��/��0x��*.Avot������ҺR�k��-��f�)�>C��PX�"���{��
��Y�ʈ
�^�!7�t���e#��3�X��k�a����Y/K��`T��{��T89���܈���|me�;�.�𣃮��'wtۀ��Zp?��K7j�]S'iEg�λ�$T��~ ��g;e���4&kMkG���I��@�X����G�6�iI���D2���g�Ȋ��w�m@�M�'�'�)�O�AE�u�����H�N��Zη�DC�����P��!��C�̼7�˦M\a^�8|�p�8��#�kzg�k�n�~�ޯ��`��8��*?�!���"��a��Na�.����,$����n�}n��|bCÿL�h,_K����>�#��: U>��_�U�8;��:��Al@ʿ����X��&h�����pw,��N�P*�.������xU�d�	���K�?Yk~p����|(��y�ӳ�p�=M�q��\}1R�x# P��
��u�Y��#�}�Z;�ת��/�K���:�d*�~,ѓ��,��K s�&
��=��� u�j��IC�n�'�~o3w���5�y��[XK؍����_2�]
�əb	O���<����h��䨑�ihr8�t���O'��抠��g�Dȳ:ĵ�[a���U�5) �:*������u2L
�3�COd� 3�j��&���4���v&^6��""��4X�S�$69,�|?��C�(�\$z9&^��RF۫Aѯ/]:=:��	U(@a���Y�|���� ��s�jB�h���2����p&��JR���#E��-"��U/K�ˎA`����Wc����h��(@�y�����p�ӆt ��PPF��\����-�R�Q���� ��׌&�l�[�,��X�c&X��.���)���5�N��Q���a������
�z]�$���-��!��]K�r�l�=;e$�
ԴGf�Ĥ�vk_V�,��rz٬�d^�&�����B�Eh��3�O�z���)L��}��cD���~4�yD��r����~\Y�L�I�J�_�[�M���|s#��܏���6�f1Bp�KX�Gv�z��:�����5��_M3�9�	�R���?��]9z��nbK*�׼.�1Y'&�j*h��5Mx~~���p�B��vLàՖ��O^��a����;���K=�Q��D�w�_�h&�! k�;OS��KsQ�l<��œ����������;uܭ�jF)����� �{oM��J�P2�S:��l�a	�Ej>E����7c#T��,ɽ7�W�?�n���$xF	d��>�k'�U��J�a�M��1԰r�_��"�t����nu:c1}v���#��^�uo��~*�;��F6�gr{RH���R�y���,g$��)��h��{ ��~ɨ"A��c祛���N�+c4s]�t*<u��l���[��`AA͑ߞ��Y=��K�a�ݮ���ta��+�a��a���Ė�q�hJ)с��tx�fZ�����@=i��fyFȟ�w{�f�*i��#Pjc�w7"<�֘�v@�<��ըA��\V�@�C<=a��K�J-G��n�dV�l,�3R#CY��x*��'ԹN����ŞϨ����!h(����_�)�|7f,Zh��s5A�6u�+dؖ����p��l6�]�}_~��u�v��[p����, 0�Z�?��pIS�=1�V�A޵��]f�.�x#��2��.��%/�:��L���J/�c��1�a~�����ù���I�:i2q*G���	�o#��ي� �$�8k]=*:�3�vYʁ@��2��{-v0�S)��.A��)��V4\�W��q]�r��ǉ�|�ynz\:R���#��o����&E�ݲ�O�	����=�$�	�!N�4 �~e{�O�� N��_�G��2|Y1��)2~�DI~�<^����.�U��Ҹ�[�Ź8%�n.�1[�->�4���Z�Ĩ��S�!O�P������8X m�����g8��O�a���B,�Cz���Ü���'4�X�s��(�bT��"}����e�x*�����K=��.�S�s�5h�@���=�=�Z�Y���Rql�a�	3(w£��n��E����x�;~��lz5����4�/�̲36����o�]�7�D�>|��<}r�J�!�� �)w��Z�9��s-2C���#���}���(�"Չ��bQǈ6�+k��)�����m^B={zb� ���@�����<m,*s	$=.����6��%+�\���-2e~[�5�;Mx�s��S�vU/�V����Γ:�A`�����������_�\������6W*��? �:B���4p�}u#���u�*�.�)�:E3V�,������S�D�G��Z:�Jգ������$2�j4�<Z8&�Vd�=��
ܱ��	N{�⋓R
#Os�/7��/YЈ�\<ht�"HPqcC��EE�o��d�ά����3���!�<��$�����T��M��7q��j�%�A����U�_4�юaB��ZNU޻ء��e1J�=�@��Z�BΉR$[n���KN9mK���J�"d����C�܊_+mr�����v%��c0�[U�6H�N*����u3��0z�2!�A.��V�B�H\VSuz(�T�*�����lX+C����E�Y�B�9��b8E��������t8E�q��t(��=p�O�UQ�U~{�F��yǜe0N�i��@�/c�T#������vN���eld�ю��+g����ʣ���HGϼ��<��=U�@j���f<�?E��+��/��׋��;7�9��S�QD��ZЌ|��l1g���Չ�}� �")��R�+�=����߬��r��|��h��c���%�b��|��ٔ�Tm�!&�ކ����fhҰ� �%+'k��È<���e!f��w�4a\#���.�
J���0v-IO�s��]�w��Wǘq�_�+��Ј�%�}�c�#4�]L�Ƴ��#y��ڮ�3ӳ����}�j*�b���ȁ w=�d�v.d(A�UL�=�O.PM��ſ@�2N*E��8�m�]��E:Q�B8� :��p�/�D]JI}m7o�W=C�� +���K����yh����i�)!���8���gաR�z�Ɉˬz"��*�5$lA8S���D�AX�G3|�8��{N�+��	�SIa��4�gπ?v؎���3Hz�Bs��J��g3�m� :櫻��(ڝ&��2q�Q�$�Ǘ�Yu����R��:��`��W�B�X�*���a�4��e2b��>�3�Q�#����CꌭH�2�;5���.2nq��J|p>��q2�C�����af"g7z;�x�K��u�4�⢶K��^�?0ruA��DoX�%4Xt���b&�T�ͺ�Y{���"@��W����Dmu]5^~�cy�cv��ۨ�!:KE
�=}y�.\w`��t	�l�ݝr�G�D��Q�0ԛ�bp�P�0��	_A�	���,p�#b��K���כQ-�\!��%Pd�<f��aƥp�Fu��Ф_vęT�QƁ~3��fJ&����.�S��ţ��� �H�&D9D,;�/��V���%n/k�L�8�:_���2$�,(�V�{�9�:�����Y�j�Bc������]�	�G���F#����a%�F��Kfk�W�W�q��5s�u���[ԁ,j-���R;0���X��k�Z��g#+���=`�l�f�ؽ7M=�1w(Ǳ�=��ߪ@3Z�m�N�6uM--��'��>���v�+�	���]�]�>d�]�9�� �C�T���:�������x`�A\���]Vue�ƭ�3*`�J�
�~bC<a��Q�>���r��?���y٭T��d5D;Q@���j%6�j�Յ>]B��1����'	4RE��!Y�=�!�ܹ8↎���S*ir��M��*�'����"�8ɪmg����������*�a�E�t���U���E�����ÅKi��yt�J�9$�捍㢤���7��p�=RG���:��,��K@�����XB��6�4|i�"y�^��Xl��� Sj�qK��?ˏd_�S� �"��(��>�V�5��~��d2'O��X׷�&Ϊ�"t+�_P�4P9���g�ԗ������!�ᬑVH_&J���č�W�}���=��p&ʥ�Z�*yv�n� ��*(F(Ŭ��&)��@{f���Q�w�1�Y�敌�!�ԪБw�k&�`{��"!��'5�)���e�]R6�ܩ��dc�k:#.�u!�+ٰ��)}�B�F������c�`:��u�Z���L_._�5��&���C\)�%��d�;*cQb�'��b�bCK�PЧ�����JF�)ꦎ. 3�ݠ�om��}/�"�V
��1"�(�u�y=�����^"�!�Qە���8Hm=���c{X쐗�m���\���
>�1��t.���9V���$k��-ڳ�`B�-l���A�}%��K��v>
���U��9f����F2���N�y����I M���]q��E��K��Zم�K�>�mɉ��;��|��OZ(Ec�3�ؕ�b��r8�6"ڑ���a�&��F�Y��`���w�Bg�$3�ܤ��r�]r�jՓD�f����K�C�����E�w�[��fH�e*q	BƗ44E���� $������J-�Eފ����/\r�#�k8���;@fOp��L~���W��Ѫ̖�������t�؎~mfN��ǽ���Y�e��� њ�7�H6�s�f��h��u�����ַK�Ͳ�~������JHJ�画�2����\���B4�':Ž/Z{L�6NJ��dW��h�Q*ç��wa���²��b��Z=��؆$�"���3�ώj��=�e`7 ���5�ǒx�Y�B8o���TW	'
�f�H�/�"0��I{V���.H��활�5���!|�@�?�d�¶f���9V�j�@�lz�;8|�A�CN�V��L*���9RAur�����P.U�>j��f���'�MV��B�K�zm�#2U=���[<�;�߷��~��:�v��N�%�����v���Ӊ~}nZ�'c���F?L�c5�s��)�p��2�BN�(aѽB� {^�GE�ut���h�!eՊ� Z��\�)b�:�]���};&���6���Mm�␄q-c&�@�N�(|�}*O+���<?����ڬj��
� .0�mƇ�?���j��S��l���B���U�y�����d-���?�~�}��9�C7	�C��כP�'J��*DY���%�rlȚp�m����t49��+u���W���X�^�=��<��c���jq�	�-{�1�f1&�:���d�����x��=�
j<?�_���3"��v�ՙg����R�WIq����xiH�U�h"�S����['��#�l̠�wt�ĉ$�X�K�J����[pKr$,�Jbj�L�l�[vT+蟏D�QCC�W3��ڝ���47���皩#c����[X������MA���L($�C���srL�����&��V�I��F9�$�6Lڧ����,��V��ü��i!.��M��l��$�o^�/P�6��J���'�(T��G����V�4��^�M���^�_�+=�Bc�3�̵I-�T;4�~/��g��9�]b	���B�ف��8e�o������LJ�� ���J�\�͟�̀'7A���U4.�<���v 9:�i�`i�S�SF{�������U��2n<�,�Ε��
����s~]ߛA�a���#i�]=
$i|*y-SA.�
#)�d�NwwG�,]����[.Z�����9�X?̌��L� ���LX�ѩkG�]���W<f02%'��z�Gz'ΗO`�3�8�����K۱�'Z�%c��T�fW9Z�X���s!�7bI+]N+�R5�����m�5׹OC�d�h�3���ȎdSIg���i:�=a�Uc�4�:�l�$�S4Q�>n�2|]���������~��4{�2�2`�zȇ�'3C�onk�q�.�k���aNy�F6�����B�g�O2�u�6'U�5�P�_�'���6"4Yl����x�>Z7�hX��
� ��|�����%�	�9
9y��&�t��Q��@�$��V�I�o���(ſ+_��I��#G�!|�JIS>�p?֣H�
�J��SM�G�r���:��Wg��BR��?^$&o� �ن���=u�ޛS�kh1���gz$�w�:�j�vt���Y�r원W�Ȁ��YEq�����z��Y��C�XkQ����ۀ�j-Yۼ���f��|Μ�������xk�y��υ~�f� ��!��9��
�U�$����3��NU�!��� x3��F�T)�y|%@���d�W0⬀w�x�<a����qJmU���V�W���kN���L�S��#�Q�a�Gp&O���9���2Z�׍���Nk��,8�L��f���븣��$uÔ�����I�2�&�<g�9K�T]��#@��U�)��`���Wa)�/�m��(e{~��C:�@��w�8��@Qn�y-!W%�Q�����:����{e��ݬOe@��0d���񔹾(Z��������KD��� wH֙�J�g�|S��	��d쭈�������E�C[L�F-͢w�ͼ6t[��}I䳉�at��P\��}��&!�hي�ԼďBMj��A9T�yY%^�W���;<�=#2�R�L4��j��*�76�St\�Ԣ������ Yh���*�x�[���8?*�D�����t[,}��Sߗ��~Z	�J����娷�*Cfc����B�{�A��d�jc�p�s�w]�KY���7](RU�#X��fH����.����w!����	����|Gnd�7�����.����t�Zk�;�
>����v�Z��P����
�,���"���=����l�J�G��ssE�W��j�Ca�a J�/����!�����I�?^����X��/r�������#��H~�uj��Ț�"��h-y��X���EA8U˹�s�O��#��߬ܡ��g�#�điۛ�2�C���� ]�+c�^O�/L�l�MbT���T<�,Z3U��>���E���.���&xU���ŤHP�T	��X��î�wk1���|�C^,	z>�ʥ��0�io8����h�p�{'�<�[n!�H!���~�Ć�l�"��W�E&��A�J_�(�b��j܍Ј�7��/��)j��o��o�Z'�=�h���O�(V�d��;I�˦�w©��/��t#���q�����,PM�w|�m�#'5D�׈Z5Z��`t@�t����'^Ny+�꘏��	J�&�p�"op�Z�W�Rwzw[R��V5����9FVk(`EQ�#��~�o�o�N�����Sƿw,���,7	� >c�K3~)@R��\��n,�]���������ŵ �l�\���6~�e)pR���Ӥ�cM�2����Xf������V��.��هK����cr5�II���W��7�A��0�yK�^W(�C)��(=��`��&�2���$\p�����*��Ť�{��?;�s��z�[`�j���Bf�1����Y.K[��Q��J3��UqU�0���Y���w�p��Y9=�즉�+�Sb2J�W��0٨��i���)�n�e_�wd�h�����ɓ)���GL�Tl��k��M=���B�æ7ɧn��D�v���F�p}(6HzP�T�é!8��߂Qu���Y��0�[(0�|�ȼRn�+�qM�hc7�o�Y�}�z�K�k��5�u�M�ޘ��w�XQ2K�0�I�ŗ&/�����ޜs�|�ߎ��V�O@�T^c=/�����A.��ʯZ �KC&=�\����AnKg����޵���eR�x��^�T)O���=����R>�o��M�t�;�6|1Y�wB�_��jY�~��p�<3Y\~^BSzA�^��%E �Cۉ��=P0T��U�*��\Y�y�tÏԬЯk��bôJ��CÜ�wKi	K�:<�4U$in��x�η���0l��*����e��פ�_̊����J�C�?�M��:��&{�&���ab���%ΟqHD�x��>���c�S��ʰ�j�� ���K?mBJG����Mミ�τO���M��S�`�����掍���|[�m��Az�B���d�uq8705��Vw�@u���!����>�U��	41�R�i��Q���r��/9�|.��y��(��? ��Q��M��"�s=ot�=���C��l�=�	��#��؇4^��+����^͸�t��M������qL�tZ��W&e�\z񋻍<���*ܯ�d��[X_hO�>�?�Ed`U��;ێ|�nZ=�\��8G0@�Q�aS���E�)-����Y]���z��z,}������G4��^�M��/e-ԟ^a����%P��",,��ќ@�9e�N�f���6=��|gC�MQV��B�����d��1�
��7~��2>\	�J�Bw̷ ��������KS�8�L��+S(�XC�V�3]�թ׮�N
�����H4i�51o��M�����+f���� ��jP|��9�*���^t����&]��̈�67�H$$�&/�|\��:��1�����#�j�,�#��ck_��\��J��Ğ��,u�C��������!��<���e��k.7<��N<��r&��v�-^y�V��h���a��v��.�Gە��t�'�pBe(���)\}�S�B�v]n�R�������D��ؠ½N�e�Գ��3�h V�J���L��h��{����Ymw� nI�s��0�p���@��Cgg�t$b����uK t�( ��Y�#?��Z��{e ��g��:�!��Adq�Y�!'�|���%ߊ;a���O�|C݅��Ŏz�'ײ��8�퇿��Sj��Y���X��a���x��h�$�P�f�I�?�8[�����X��	�����J!8�Bx�zls����E��l����ݮ�{���3C��ۏX�Se"J�kD�����T�6�1�MO)�y6n�pnW}t�}ݹ��,�Î��� ���"IF`o�����ct�%8>㡥�l{fk�JEӧ,�	ۼbCn�b�F�I�����6�M��$i��ʥ5�e������s]� ��{՞*2�5K�WֻZ�j��$,W�5��x�o�i���e�	�	be�����G�։���Z*}Mg��+�^5�J�tԔEe쳙L�n�����������Q�1e����>��e!����r�EP�REX�fs[i����1� =X�F���RԔ0�YH=����
��`��l����Kq@�f-�԰"4�U,��9W1L#����[]������BNL�B�>��B��^����⛘�_H�Q�S�+?��6�"��e�4ys�Y?��Ⅶ���p����XhKtKw�����/��&�~�0#��vh��[R�ݏo�s�H��ʄ}vY��wS�\� �4b�+�-�����/��Iy���SXn)�-�6 (W_ 1��X����Y�h��3$Ә,�.�Z5�(%�%���o����	�]
�߽��*�ү\��u�0�'!s5�n=��_DB�������o��͇I���$�h0w]�y�|��2�10��#�D�QlݡS�7$�$m�����F����i���UYv~��FM���'iiO�%��)g�����_��QU��bU�O�½Ċ��R �/�[5̬�u���a��2���]�f�
R���nEmO[;�.{�^�*nB���-g�l�`�U�W���5�hc6
������P���%=AR+�����AX��Q�l�T٤�����
5)��)�?��c��f��ga�@V�o��yY�ң��?%]��G�=��l�g��!z�7t���XW7��Ԑ���_u
rz���(I͘GuA4�9�饃�5ۊ�"��L!8N/sD7�$�ݾ��yFn�M|vi��fͰ�h�c%�J�.��G�����ϗF�0֡��${��ul�,}K9�T&Mk�)��<��*%P�vxP
�,yqS(��1�R��P��*��݄��V�~N�*�W"C�G'�^js�M<�`��<UI����_ w"!�O�u��rhr�em�pv��n��̝��$�!�u�+Ou���x#���ޙ
�P,he¶Q�$�"���:GA(Iӹ�s@vF�@���pJ��µ�b�*@��{o����RC���.D�s#�?T����~��WSu�4\��O z�4�d�G��؏G}�V�_Z����䟣�έ�q�#W$>�<*���h�rO5�kSHi�+�ME���(_���*��l_U��ht!2�����@����ʄ7�Q%�2QK�O�G��.Ō����x%,*G,o,N�r����e3ۜM�5`�S��B��lW�"n���p=/����Yd���gU��IX�I���WJ�� �g�0��#�;��OI��p��_ۺu�`�^�D[LE�L��#O���a���:�+-#(qZ�)ӕ�tv�w�:�M�Jw��hf�cKAv�yx_�[F�D8�T�R'�Hi�Qq��@O��R�3`��Ț�]�0Q`�»�;���>��S/�#��V�k��-�~jtu�-�FZ�{�Z.��4�O���,�|j2g�)n��z���b�~q��O}�F��qm-�T�Z�G�r�H���ԯo��Lfn ���.Ԉ>	0�i��8�S�S�0CۆgP~��d沏���WEX(��(�W6�E�(}��6.