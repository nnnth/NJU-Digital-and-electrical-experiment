��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�Z��K�9���4���t����~D��ϔ�Lm9G0�� Meȯ_� �ny�5�����P��Z2c������:���4�-�H�@S�O�]|�m�w�>�\dq�ayoҳ�Xw#lm���8a2�E��V�V���+���0��Uq�8�����K�u�c���B�:�A�א��ɅB�����{�:6����$�i��Y�TkU͂�iy^�^�{�(��/� ���vS���������/me��YJ%k��M��jm�$�-��xTn�9��D�/���Q߷_Y�ڜʰ��C�g��?B�FY���apu�R~�d����{1��Y7x�J���G�R�!�>��,���h_D�ĩ������FoW�~��)=�3�������	���R��}7�Ը5?�'�do/>�+�}�"<a���Ӻ��Ķ�ϳ�g�4��lI���'��"/�WV�Ջz��4?̏��{',[�Of�ON�X���Np|���9w����%b6*�������Fs*gg/�.�� ۪
Ҩ�R(�'�*��]�+�Y
�$��>cu���>K��k��z�M�i��ZjHL�&N�\��%`�� �E�t;{���νl2���Y*i�)��4���5ٖ��j`Vd�5�^���I�q �t}o­�+�j��+.��\�X��g���!,�c?��B�����A�):�n�Z"������-?�<�a\�W})W˃�L�DK6�7�6��ܡ�Ԍ�	Z5�E�	�}v�����f���9	%&Uk��#2 �%�2̎a�P{��E����EN��?��[~0�e�����.\��f�h���v�B�uک%�> �\Tv��J�N��Ks��q��������V����t�w��ʚ("6�æ�����LA~=e�?����z٣B��\�����$?���u�ۡ�T)�Z�}U�n�͞~/�ӫ@�)���,�+s2�r:�����s�8��&8b�*��;�_�H�=.��(G��Z�+���
՚��N�w���	.�N��ٚ���)�9�U�qb����-Ye�S��Ѹ��/y�Ǝ���Յ=�6�|�_�[)�FZ����Q�AB�&�t������w��ټ!1�H5�*�*��d}��K1�&Atj":i@v�!������I����BP-��MP�x8��+}�!p���6�8V������QV�/p�
92Y2fȦ��m�݀��C�>/�A��'W�I�cmy� =�A��Fl��1ITO�Xn��=�B��Rb�BuSާ�-���)X*�>b]����W]���� ω���wo���N5
M�s�ːD����[�u�}=���,��0�};����=%�A�מ9l.�i�e��?_U!ķ"m���U����RWm�6W'�ǺV����b����sD"��D�5N�.����N�j��0�z��2W�>�B*�HP�>�ᓾ�%W{Dq2���4���z�qL��=#�ys����F�BWw���CҶ<�w�#���̜"�Az���<;Z��8V�Փ��<��gc�Olf9���W�`������W�;O�l�'���=8ڮ+�#�H_1�����hm�UN/�f��&b5�͋�Ȕ��ȞM�D��3�S�|{���>�F�-��cp�ٽ6OW��^��>���M�e�]ܓA�3*�o"g�����<c�و�e�u�mrN�!r���J�zt��p!�dr��N������$�>H�0Ҿ�;�����_a��Q�J�JC�
�V�<��9ɖ�Djl���}#ev���$ъ�����S����gCڟ�(�M�"���w�v�'�%��)��2r랎EEɃ%�����v�ϔÄԨgDh���ZG,��k��P���䄂4At1@��I�
��b�3f��"t�m�=;�����gW�z�F�L$�y��T%=�A�W����	����S�����:���<�p���(-�Cz��_�Mc�yۤ�B���	Tm �^ml8f��i�	��NkA�z�W��F4����e^y�M*���K{���"�s�@W��MP��Ґ�2�i��$�O�u>��������϶(<�{|�x+��.�`�X??������R�Å�hMLn��:���.K�h���\p���w�n	y�6����7*v�jexzȧ$ɞ_̚V��v��F����ʔ�\ģ\^�Ě@%�� ��٦�(�Ă�e��ԁ?0ꋐ'��U{�ߋ�;�}]�%[��:y��\�#_����.'�������2�>���n�PC�[3K}���&��U�Zy}���	)��ש�P��UR(#�Rƾ&ռԣ9���^,{�h42 �RA]�b�G�IV��=B���1}FmkRy���Y�t�X��R:%?Ar�[zUI5�Z����;�ʌ(gM|0I&;��Y���X�k;���C�,���}+��ͺ�9y�ko(j(w6�jGѩ��s۹UI��M�������=,���:l2"*Bcd��ש2q���L�2�H��Z���˩M�z�U\pq}`��S�\!Fk�2�?��A����{g}�_�F�x���ɜ��X3��V^�l���⻂�wEXqmmCЀtL~�s��JB`��B�K	��9G.��d7^s���ɪ���=]l#��JTvq�`ǀ9���rm�Z��LZ��G�$�.��I3o�*EW6l�rG8��r���t�'H�������$�<��� ݿ��bV�2qH���g�V�������Y�r�L����a����L?/�\��a�'�}w�#�uD�[B#]F#��g��N�>s�op}Ae+bܶ�2ן��m��aR0�0Z6X{#oH��J.m��us��D^��C�Ѽ-^Ē���RlÙ���3�:NɩS��2E�3���9JΑ�LS��(���6N�nHW=QU=Q��z�%ӽ`��g�`��x"�xc�>g�����mi	�i�>� 5����h�Pdm��'���	[G����n���0;���[��蜰�0C�O~3�ä&ķab��-�܉�(��2��E'<$|zOU�@��{���樵�``]�ChQ��oY!p�p�!����R�O���Q�F��Ӳ�Rݺ�R��T4�{��`3$u����ֻw9�N͍?�D�Z�S���A�V9cZ-�$�B�;���~� E�+}!j����ß7�'WS��mL�m�T�;5YG����j�N�n-�z<{�1/x�ۢp���h�7�I��e�fa��\%7sC��j�|�J�m�
�rN�����(��.�nK�2��x
$�<��׮YS'�f�-L�?'�������*@x1�FO��hH���5|2ʏ���a�Lf������"�{j,�9���q���`!���j�$����Sl���[���"oa��w��2��IS�GӘޥ�7#�38p�m�zK���ϲk�\�iV�*�bd cB9��+����r�*�KX����f�����=��5V&"�Wnƍ�dl��Z�t�m�2��2�ґfv�&"�6ɯ۶x���}�֗Kj#׉�j�NL�Tv�)>X�������nYW����hj��m�O�&�cW��y*-�!���;2%�N5�cL;�Z��-�!�Z"�z�Z���^�[䭕�hs���薋FZ޶��	-�&V���pe:'x�e�^kg�_Pl7��A�uw����YvU�����ZI�N���%l5�6vG1܋��͊��6eػ�@�~�bG����g��o����(�I	�5G �*P Ei�#T�c�DSX��� m"�V���X��|�����dP��� W ��Ag����SO�Ta@0��zB*C�pfi�  �lc"�!�X�Ɣ�e���q�ͱ���ڨ;d�=-wf�ȮVù���M�o�q�t���[n�k�b?�.�D/�L���ġ�7�gГ/�JY�V��z��2sd~��e��`5���@�Z�`�J���.���8	#�0� ����4@�M�/�Q3�ck���'�s���̍����&"�����2�-{��0�\0��n�:�8�^�M��-�FpƨF��ʙ�k���Ӻh�B�� C�b���J���;�=:%J�tc ��<e捓�T������WY�Vã�yd>��h���c���犆N���S�q	���[��O�7��,�m��]s���#��( e�x�M�2�i��d��|;�; ��ᇯ܀!P7r�+/A�<yEv_cKR��:�E��jnaA��v�_�s%��ܶ�r����4���x~z7c���x�m��b0��_�F�&��F�e�n���S��5�W��6�P���,X!����㺯��ˎkH~������A�3��\ �G�!�J{dc
��;-�B%
N�\U,\��exQ�%e+~`��@������nɲ��V��v���$f��8'���X��(�X'v�����?�f��}�TӧU���fz�¥�X+�r��'�/�û:hՖ�oLE�rt�/%:n�$�������Ьڂ����CV_�&F�29�g��nsaS�PS~�����_ǃ
�
�Y+��}aV���?�đ����i|����ԟ�A}���j��=�D>�c9�o�
@1
�	/T��6СY�k�H�� eu��=�:��,ʬ�t��rc�]�E�x��Pvwr�(��G�Q�a����[q�~J�۳�hm������\6����?q�AW���6�,r�Ԏ���;��Am,ɴ�c��y��n���7xn�A^��/��=�k�	�)+x
���w���Ĩ�R�Kj��é�+��g�ġ�����:�s= T���rA��	��=B#M�<Uy9�bֵ��m�cs�����0�qs(�b���\�CwP���c�vj�y�JC��o"�Q��|8�yǲ��g� J�Kx��u�aJ�s����7�oZ2m��N#-�%���_�Q��}m=,�����;i��j�)F9Y�u�4��w�)�$`����*���s;�=��a�F�ͮ4N�\���_�X�>�C�o؈���[�0W�4�|�RU���8��u��8)�~���E܇<2��@u2���p�M��$�&�T�k{yh(����E�(���f䒟u)�g:��.6�'A]zX�WMv��� �+�ExwD��"i!�K��(��R�I0c�!�@�����l=�wE0�Y`���/وb��K��<��j';,��yp�g�A�WU����)�"C���{գ���-����ӱt��[&�08��i&��A2�77��&;���0�g� �k󷭢Zi�V������R[���h#Uq��/	O�A�?�r��k�����3۟�~u��,����n�%$�B��*5p)%8�����=̋g�N(Y$����\l�2)O��Fn�G)�����|n�'Z�V�h8!������G6u@���q��>�R|piU���*��`�NC��Q�]�>U�?px��xo��2���w��Li�U�	�:.:�L�߈��a�\rh36��k�z��t���*\��w2{F���#`2�x#K�}gʜz�M�������5a���s���:�,]��N��ǃ����O����z��=2�{�{#�mڠ�0
�@�$�K^��Z�� ��c݌s�>i�~�
�TH�v�]B�luS��r Қ��{�����+��C����m�z̼�M�d�WI�&���@�D���	��:�g��l[��ϒ6V�����q��ɵ�w�`|+7��^��9���+`�V? m)G��ibT�-�%����'��f���[�̌�}�����Ɛ����v>���BD�F�6�^�o���gh��A��0E䗄B>��n*���pi|�o�k� qazR��Lη�-��qS*LH��z�s���� ��<AZ��E������2��Zcl�.'g�G$�l���m�XE��s�آ�D�<�y2\�O�ƣ�I�Ԩ���O}�A�97���!#HZ6	�5!����ƒ�����Y�6��1ꤳ�z&�L�6Gm �fF��$p�p7v�4��%��pc����f��6 T	�ũn,�?��_���5�D�~�?��o;�P��e�
$�-K.�����5�#��νH�T�k��x �XgY��h&���D2S��X��H`�7�c�m$�0r�-�=U:u����^��!�H��覽`p�.�8?�D�K��o�n=n&�W��	���#!fA�d�:������l��`*@��W��=�@��2:d�R8�qw�*�y�|<Z�UK[�5X��5��#��s�'�A�B�f�k��[*DoGkI�Ku�[V-��>��-�eU��'Z�V[bja�.9���NCU�H]	�Y	 ޏǬN+�S���U��\���ֿ@ߖ�b�����Z�*��p	٥ks��.Դy�!q^D�n@�%8Sx�jQ4�Q{�ɉ�W�NwH�KIt�l�\.�D�z�1��"� b5�xXd0�GP$�/��R��L��z�4���\�m5A���N�u��5Vz����*-�ӝQ�Vx�=fB�m�0`�#Аp箢��\�>�GA�T�m�W�Z�&9���ug/%{Ud�o��D*��/�A�Bf�[F�>9�a��W��Zf�}�n�2��r�M`h'p���Y� A�#�$TO:-e_xc��!�}?�tNBIka�h�̶�A���0ĥ�`��	��yi&�q+c$y��}����/� 	w��fɬ�rM������'S���~��}C#
"�M�3��.�c�?�PQ��Q�1M��/F�u����T�&ӭI�	[���?fA��~���F��=�
�m� �6�jʵ�����f��mAOM��~��G�P 1�^tp�Q��$�z7/���x#��:\nn�p�����'���A���I��l��/UIZcء����q�cE;e9*�K$��s�e}L�L�� *^G뇞���2ǆ�DQ�*��ǝ���@�?aL{L�7�8��d��#���eN&;	� W
�E�T�EN�/$.w{�̂��`D0����+gknGw3uN(�$∊!$/�In�n^e��IB%h!��㾇�e��S��e��_�����ʱ�QJe��}��U`�rOq5N�%����uv��}�ڽ� �8����x_�p ��+I�'�gtu �S�P?����UI��ω�/�ƚ���>��7^�����X�v���<�F	������֩;$�Gf� �acoJ�2�ӎ�i�3���{��Q!^��%�8K�����}^S`�
����&��{r���_en�<J)	En�$>��?���m�U�U�0s,��z��t�ayݣ�n}�B-���9�����L6���(D<�k斷�x�i�(���%�>U���m�������7�O����y�-:��h�SL-���`
(��Z3��Gl�Ea7@���-.*C�l��54A�@>%H���D!*k��������U�V���#��Nճ�����\�TG�B��� G@ό=�㉞�9DȍE[�n7r�O�,�o"+J��Z=����Ao߿91��'��zɓG�5i�1b�g��D%�b�^f�ṦIS!��1��/b5EJ�b��nOp��Q���-��,'�6}^!a7���Y����A�M���/�Zm:}�E���<��r��('݈&�h�L[��T�u�,��hP�ײ�,ia �QU}6�R�Y�"��`�md}����Ze��!ȗ��i}GY 2�����������#�0�{aYT���`˼ ��ΙQ +'��,��+dLn��[�T�3}�ښ��m�����0��Q߽�Wq�UZ|��M�B!���`\W��=�W֙�+�) �k���ŏ����D�`NFuLa�����%��%��5�ʗ��k&Ō�㡨/���
��x��|��M���r�a2
ucBsꏷ�� ���L=����|or��Du��9��l-Ԝ'�������r�F���=Yށ���3��z�wM��DQb]���t��~�	��-a����πj&q&�Do�k*.
��5�T�� ��Ge �y�AVM���2��@Gg%%<%�`f�m�gmT���i���9
��ހ�7� �ԓy��X�-P4�\��T&IoE�L,�fŕw馧����mr/��Yu
��to��l��.���_�z���!ۂax�mE����1�"�l��ͳAi��7y5��%�ˎA�M�JK��]����eQ��8?6��z;�m0�y�:&@�v����)��҇d��T�{hB�æ�\��{����!��.�й9&���tEP�7<K�	���L�*��[� .*�k,<�7hf(QHÞ*����?�,�P<V��,�_4XJB��C��W�A��Q��F�
�����L�r)
X��7i���Q�/����H��c��Mb�%K�'z�������Z� 5��Lbl�4�o=� �l��P�ƹTS�G�hC��I��\�Y���UN����C#�;�t�$&����Be��3J�وtޛ�7VB�Ck��tt����D"?���L�N�>��E�0ٹ��Boj�rt�f��R>�=@#	��	��⫚�[Z�<,7)$Rr>ST��N�u�M�'�]bS�>x˃'�51i���yz`��D䎣cAVy=��rG+��cߒ��H����{��|���0�} �-�Ն���1n�i� W�m���Ď�)���2��x��ޤ6�o�O�*�!�эt�F�<�fm��[S��(����S}�am�������C���bs�a�^Ux���QA�e�˯�T���1��q�-b두��u�  ?����Qn)�)�xͥ�vF���a��ݑ�D�� ��>_#|����t�^�%4�e�>kC|o3����#�`���.���03�>�����V���� ��4��mĻB$��=|�8�7R��byJ�C���ì��|�L���0�f�lT6(:�s���Ye����G}V�-wL(�GG�	��P������F)����I�C)�D1�5�E�ۂ�9�$�kv�2�ȳ�)� /������+.�)� 7�ZRm0�mU��
��fe�U�bSS�i,��D�h����@�O����n��jA����X�Rk��aC��,���ce��EMS.~�ʑ����&<�|�:Aך|ݧ� f.Cx'�F�qT5��� 5	#c� ��i��!-8nʃ}.b)�.&�Fm%U��S�"GbE��!?�l;92�JB�D�]�,M�?��/�dl˸R�I)�s�۵��P��-Dk��:&3�cc���
��ȵ�+Br�����E�0�'fT:v�L��[~����y 2$$߆P��H����ۍ��n�&	.�9x�Fuk�Q~�O�2�����(�	C-󛐠�>s���=mI1���V��.�O:�v+Ӭ��Fc�M�JC�c8� `K�ŘK��Y��0|�4�|�
킂]��ch
��^`6�Ї�0.�k��K}�q�����3��m2&G+"��h��Et��/�� �N����A�9�a32������N��Ƞ�i��S�9�2j��EHR�r�F?�C=FیЧ��0ҭ�T/d�N-`(�׆����L�T���%-U���{�����S�Re�m�b�+c��!m�?�N�׏�x�� ���LԁI"�8~�X+ ���>���Ԍ�j6D��d�x'B�
z�c���l"�	\��O�$вQ�A'���no��O*�;�\i�06�p{�#67G[��_#�!��{�O�Ь����=��<7��6c-�ɻ�V��|9�0�n�D�����7�s�B-��� 5�P�#��������k���˱mF��r�|,�ԍ�[�Q/B�$k��&js��5�{�AſX���}Y�d�F���m|�5����d��=�F�9��3_��NJ�ϬK�[�����`�q�u�y�Ln�H���~ڿ�Y1z�$#�]��c��o�q���<eNBa�}�F�39��M��m���h�I�6$�g��Kt��7t�4������)�.���r�iy������0	dg�h�jr+&`����Sn��ٹ�e�,��%V�Z�0
�9���Ǟ�}!�3r���N��1��S���ڋ���:{1')9�y�Q0B��E͆8���OM |�DI�(�.mʟҭ%'!��E5�����d���z���ۡs�����C~��p����������t���zA4'�h��G��B
([@!V.9�Qbx���.�3�Y	0%�|.7��x[��cK�-%�.�0!�b
"h�m��^�������[v��D{�F97 �NU���+�f9vk�:�߻�wǲ�p-����{��
�+^��Q<��v8x�_O9�2�׹y�M��K��G�f-�@��	�����Nh80��v��С�}Xh[$Ɵp�����Ƭ��ǶTY�7��R/�@^�x�epq��l�:��]�?�^W6���/Ƶoy)�+�̰��t�*:�}���)�uս��)K�����2��bW![�oy����zum��x�J����$tis,���ו��Z���v��Ů+���,YKSNg�)��\��ȫ�	b����j㿜ٍڈ,�:ũ�_OS�$?�)7T��X�b��)ɔzS�
>J>��kL�Z�;�����P�+�P���I
m"!o� �A��-l#��I�ሾ4H+�t�F��`��kG���{#�[3k�8�!�G]d6���O�(�-�ɠs]�<ȵ��#��~Z�ڨ�����~��2����S�rl��6l?K�\�F�1��뒐���8���E���������͋+�Dۚ�:�<���;H���c�Ű����rxgm;5�C0���Zp$OSA�;M���e('��]��B���>F�6�4<�UW>O3NS%^��ܥ�����*�_z�{V[�*��W�Tβ�wtPhX��I�6�Կc�e Ц#E?�<���ߜk��h��
Y�@%��F�!��ER ����udWľ��� �B������]`�(T�֭`c�(������
H���;��b[���F%�����'u����sT3$�?���ˡ�/�"��JH9��G���mPc<~�Ԩɱ�Z@�#(�X�K��h�Co5ׇ�� H~4������"h{�V�ŧu�%.J>�)��=0���������Ǻ0�������V�z�V6�<����F���B��Ƥ"�0�c�j7�h�֭jl�z���6�*S4@
8�3�n�3�'�Z�R����KR���!�o�\U��R�����fPXͶ��{m��*�YF�=���q�WB�#ܸf���D��*ͯND2OH���úm0B�CQ��'��m��d5U��|E
�	o�t���i�LpPZ@���M�ku�&�2��#;0��^}#�����6�@����U�6YW�I'�J 4��1��oNW��+��� ��T�0.Ro�'�<�� �4����li�h���U���ȹ�w�����
�t����Z/�VL�7M�@���5�,��>&����p%޷xKூ�|�cc�WB�)�����v����u)0$��#(�v��~������)�D�u�BE����_�gFqu��1M��Ͻ<l?u��a�"L/��Ǎ^u�0�r�,�,�㫩��8�+,�yT�����^��7fi<%-�`vr�P\�زR��./P���H@#����\w�6�2���q+�)̍���Qd.�S.K%�<(�}&�s�ӂulG�@��ѻ��1�% �X�}��״���u���;��1b��-j&�����-0�E��;��YS�嬛�)����'���RP8����4�B�ab*it*��CY��=6�3#��o�����fOFK�C�ݡ��ee���/��6ҘD^~v�A�Xb����0�6^@�t�Jݗp�t_�:	@�5k�H�[�~����$/)��'�`�)!t�Z<w���{��*�A֟�2��<�2�W}�O_y_&�w�M�s/���5N#R���M$^���F������R��3��:+�X���M�U/ž����@��!�(7�(�RI�l�W�i���@��M��˲*�x���A1�X�B��a�����@��
��nL��ْ�ogL�ɟ"�t	}M��'A")��gO�Vn���@�0�.�E9N�U:xr@��}������qmga.�7�(��81���:�D�L���d�r�d��wF�5 eueȿ8�Vp'A+�&4^l�����J���1hK&�����7�:*�8��U$��uNq����E����l�u���ʖ�1Ay!�\PWPm�� ���
M�x8�w�sU&Z��(�����$�f۫�R.�UG�&�'#�9%A6 %>���Ό@œ�Iր$������ef-P,'Ut���x���`�S�K@@�E)�q��g�Xdow��9�I�Fur9�a/D9 i�P��S�� �XG�I�$�=/K	�H]�J���0RM�ba�c.5�"�"�nz���������@�B󴡱��)�:�봱y�V^��C~[���?H|����0����k��M���"��a��b�_��zOhF��=c�2�2��^��\��AU���0�ʶ��S�V:�+��9#���¿�B��b�Δ�ѳdn�@M�*�]�((n0���x୭��'�9-7��j^�������{�!�N� 2������[B��,��5���9,����E���R�I�<��P�AQ�0�W�m���������p&!���/ĕ��Tq��o�tס�;�^h�%]�AR�"r�/��^Fr_I�M�#l�Q��f�g	׿�={Lm�?S�H����(
 ]�]�U�雚��l���%�`�{�Ip���I��J��9��ށ#-���g���o�dE�Mt/�zImx6x����vO�?�ңG�k�G���jCz��ו�;��W"�X��+��6 Mg5u��o7��GOßh N`o�<?%��!9�G�G�QH��v�%�!�O�󗽡�6����w8�>�A4J�n� ���B�~��$�L˚�� *^S�g�5L����G�oy8Q!Y��dC�'/o��W��H�G��ȃ���\�=x^�u��% [u�@,4����w����4���_ �e�N_��I��l�9j]��	�o�G�HE%�x�=�j�lF�p�S�ST�q|i��`D̶(wm��|Lu �3�7f����'M��`�����,�]���X�>�i�)d{�ȐH�		�}�igzVaN�z�L�++���U?i�3��H�D�Ѩ�ښ���Iwp�r��q��b��Do�l����^%�s͑|	X��IMd���>��4�k�`�/�g[�s�=�/��T���ם���rj)2�Q�7)�?�T�h�	b�n�	�[���	�-ɬ��IRT�$z��do��'�����Sx䰴\&���t(���>�<�r��kh!h����pܞny��+fx=���7Fr+�Ck�=�XC�U��=.Dl�fe-p�Kߤᤪ��Mq4�
傽,\8q%���ĐT�!��dI�/���S���
o�ƚ(\�i2Y����a�4_����Z�ux������~t+�&��ݏ��Щ���}�K���4obC�<l�����C ���SF�����l��o�y��°�4����W}j���H?ȿQ>���QT+*��w�!�(�L�n��~Dey!Ōn�,��`�!�M�/M;�]Q�Cy�R~����y�l�Z��|i��.5�Ƣ�Ъv���
�<u����"�X�'�y��R�c���j��6�ytm-a�H�4�O�w��eG���Y���vM��v^�3=�A	�7�~L��
�즣C���<�֔(�����N��ïk$*x�q��a����l���|U�J���"��8!H�e�$��R��y�rP�����:3��5�2�C����q�V=��nպэVc��L�rS�1���Ă��]�9>k��H����_��u#�NQ�O��C�b�y�y�h\�Yy ����x<�����P����h�G�s[5�ż_� ��z����.a|S�*�d��f�����&/�e��	[(�ad9��I+k��"�rs��^�KJ�z�+�3<��4�G]w���
\�$	���yCx1�#�ɏ9�Wn�B]߬h����3Ը���}�h�0144Oض9�}e�]ɞ.Pܔ��s�AC�l��]�j�}ن���is�c*�­��>�%����h98XӕM<;��~deК�Z�����<��{P��� }��5�ͭ��#I��}��=}�O�e(�^[3~A��j�4�coO�W�K��_�#}Z5�H1aH�4ZT]EN�<h�;ks��� �P�EY.��m^{;���_�S�S���W�!�o�&�WeĝA�L�-m����"�������p�:���ج�,s����,��4WD��?��J��^Pl�z���w"_�5�^F�W+P��L��m�L��;����z�CRHQTF+�������Kv8�B��/�\��������wtj[.�0`]Ӣ5�=Z,k��PP�z��j!Z
�&K�!�K�A�G��a�7ͲӁ�!~3�.�'�i@!V"���@Pd'~�t7^ �7��?�ycg��|�d�W��)��=u��B��
,Hv'W�s:o�nW�D��zWW�?:��-�ґ�!����Y�2�U����z�¡�㼭�,hXǳ	$'��T�P�I�R���/C喍�U�I��o֐�	�j�o��9Ύ�(+�������Gc�Ӹ]`����MzڤtWM?�'�}.�l}.�f/����,�
&��/W~%���~�k�q��Dش`�2��L��E}B�l��\�#���m�7Y���Ey׶<t�����"�	�5�!�G�A5y"u�U��
;����Q��VV�$Dؠ�I	��{ޙ�H��Jm�D�0o�UT#w�	�z� M^/�1.r�Gz�[ ������ ����{�.��w�$>'Pf^)��&�3	ަ}S jwn�Ʒ��vV���/ɥ�N�ԣU+���8P�x�or}>۩rvn�:�'����K�h�A�a�  A>���u�����V��u��{���|Jţj�]���������^�T$ο���$&��o +o�.w7J�+�<����n�j�B��'F��6�)�P�"ð�^��5��gZ��꟨�S*�S���*�둛�P�Ӵ86|���e-]P&�sl9��))�SI�Nu���ng��b�\�������� ��C��j����c�o����m�Ճ��>>�OH ЍDO�n�Cy�G�QLȨ��
Z��=���G�Z��M~T5��a����;zQ�s$ 롖9-״$��+T���I�[U
گ4���?�*��'�L��ʝH�!}-÷g%�).F,و�Ӊ�
}��W���Az3��^a�̝l�m�`�!��Y��?��e��f^�� ��|����!�^�����uߺ�]�I�D�jTK�m�'���R������\a���v���?x�����n!�9 D�Z��)�2���:P���D��*Î�[����Q)i�pl�lGN�p2�
y(נ��`G�EΊf��
,
f9&óf�ğ�f�Y�������������Ң�yp��/}=��fa�7mS�i��x:�S��EL�zq�a���!E<�x~��%���r���w4�8�l�c�̠>�J��5?��9@N?Qy�7��>��j��O}Z^�M�>�.=�y��(���n�Bn_=pKZ��\�
ams^���	:��y�H?�����owq�JP��Av�5�5�p2$���4#4As�;��[��~]m�"���u~��R8�!��� V$�&�j]g��I� ��c�DJ�Q�1��ɦmJZ����M��#QVg��FOW��{�̯\��쾀��>�d��ð�ё�[t/'2=cQ�K������9-+����	=����o�ސ1�G��_��-lU�W2����ң�&��J(Ѡ���֝�8.?z���w%��Ax�ѻO���W�d��^�~�p�>�jΓ�wD@^m�	��_��rq)���=�9e�v�zbƸ$��S��_�@��^h,1B� �Gy--���>���~����U���ڶA�V^���U��޹]V�X�^����d"����z���c�z�}�#��ٿqd�x�ab{�=�\�UR=�Ep�k���)V��V�u��A=�`�����h��d�ދ�]�V�|�Ky`��,à��� �`��t�� ��S�}mY�߾'P3��.�C�.��p�|�|ȶ��|���U@���O�;��sm��ү}� ��]��E��BDv�(����Г��,��;)����D��ʾ���'@��#a�����vDV���*�n�T���ʂ���H��h����G����w�de qx^-�� 3�%���]��m�4^��И/}b��1blW�/�Q߾k]�C�Z7��8\8'_�a��|R�-+Ǫy��H`Ⳏ!i�(�^�,Y�_��OB[��SS 1z�%�R�7���@պ�,Ҭh�KJ�/�'%'�
ݬ�X�5��SAS)ɭ�:@m��]����Û��G�>3~5�Ի$��8Zt���|�X�E���[JK��� �!@��9�L�5;���ﹺ��mHP���8��Z����p�ȾVM�5��dxL�ˤH���u�Q�M�6*J{)���H$�<��L)<���Ŷ��lk?�mUܵ�b����\�Y$j������J�Xn�P@R�j�q.�=xԣ��+�$�Lx���rR���`��r>;#�gz�qlaP0��:�	_Ln��6��t��@���߷�r�򽝘��@C��@� ��ǥQ;Yu5��7N����
i�'�I�[�]��(���8/����0lXNs�[ꇏ0���ܗ�V̳}���� ��(��W{��נ*˹��ۅr�7�|����:s�	�(���"ar��N��+�tPjWLD	�)9.A�1���/��O�SKm�e��"��w�.�5R�y��O%�2$�ǵR.Ã��l��-�5��B|jejL'&\��L�]�e��W�������N��h�̣��A��%�j�ؑ��}T�ݙ_��2+��{��˲t[ �����@8��'ZH?K�����G:�>�,}����+����%�SA2�Q%��k��
Z�A¥V��c ��O�"��H����Ŕ��@���	�!�l�&�<��@���fE�\�gf�Ť����z��F��aKGИk���yul���}���A=����_��|Xb�U�� ����:�5���ؓ�������;!�!�"�v}�g-̯ł�ړT���7_ɮ&Gѱ�8`�B�&:~˿�C�G1e'��>�����Yv
]xVf�P���&sh��PZj�1�{z�A(�>�~���ˁ��^�8;����xi�[�T��pg~��m�;�z~�K=CCSJ��y�$?�nI���Ή��k`�P%�+2q�.�Ъ��d�с�q�[�R3�%��N&��.{�Ӷ.|L�Ӷ��oG ;�$K^i\��,ޟ�kmXa��Iu������yP���K��
{x��̽�\�� �P���ꏱS<�6�0��"�PhX_ާ�8�UԾ�x��Қվ��Jj�դ�+3�	�ޭp�m�yÂ�淞ۻ�T4�v�+��0y�pO��[f����Tmx.�ƲR�sN��n�����>0QCo��u�?n���k�7��33���I��&�݉�e�nWBZ�=�Q�^cr�f�h�����T�L���G��>�͒�C�=�C������ZCB���i���t�ҷ/�x,�D኉x�� ���SF��d']�d�guTd��bYHrg�t��n�=��`�
��i�Z�*�'%�����ڒA�WI��~�Jw��9 T�Ņ	Z'H��y�ء�1�5�j�.� o��s���&�:Q�.m�e8/��o��9L�`H�Jp�D)�1����^w��O��9%���y��h�$�����PtMՖ��N͵&�.^���`�b@8�d1ʨ�ѭP�n�n�_���M5�������w5f��?�� ��Sɤ|^l���
���y�p�� ���ʟ�%������c!���-��+"�L��5Q]�a� �h�B�c�Z�4,�������
9V/	(�!�X�QC'��k℥��,�﫛�3q�h�F6�o�A*��w�'�޽�~��:�����WK���E���D��t�����5�
����6�4d\E����z�w�dt��Sy|+13�1>c�f��ϛ�t]�z{�%�NV}�i�sMHz��؂
�];��(p�j�H'��ո�iO�|�.��^-�O�w�#�R�7e�BJx�g,��e&0Ji�/�z\7p	U+��te��w�ʙ�	�)C2��"���=KC��L#��Bך�'��t�X�TL��#�������H���$�^�߮�4)����%��zT`K!�fz3��n�g�!�r���T��$�Gd$ͪ��/c����t[<� �or�E7�՟=�8]�|C�R܅	��%�(�[��󦓾�Rh
�e���G��{�;5��j�ɴ����rs�Q|ʟo%��H�(��ǝE�RB��;(reW��HK�q [��p����+� x��x��e�������+FS�1���ہ#�b^|5~�����5��:K#V������m�Dz��I/`oh���a�r�l�����	0��oܠ�b��r5��(<ۺ��5;�"l[na�l�����ivǿhUc*�ץ�m�ܞ�$��X!c�jN	��R"D�6
4�e�"0O���)L�҉��l�j"j`�J���_&�Vx�QhɗUb 0�oW-�PaF����iW�V>#���Λ���'L�/W��@���u����o��Ǌ�18�NKW(_I>̳т��N&j+�`�K�m&��`KS2"2�geY�֭~2�����Q^rX��&��]�䔤n1L�¥u��� _�EMs`6���j�:�#�۫{4���Q��~˝��Y\;Z\�Ű%��64�He�4�R��U�a'���A��s���3��� ��iC<��D�=lD���Djh�����t�L�S6Y��u
��@�R$�/՗���L��t�ݶ+�!Yq��o�(�$2*��P�8��I��$T��.��<e���띛���E���3���{��ֳ��z���S��*��g���S����x��H4
d+t��y�\9���t�A?����gh#�U�eA�w:D������yq�g�C����0�?{��#v�W���ٯC���'�����cDшX%��������V��ݘ�hT��$�Z��%�ݗL�x�a��a��F����簥t:�sW�Q�`4d)֦��тjr4�$DY?0?BX6��	L���ÈMKU2��bf�]�Y�XJ{9{�M��y��atlH�	�W����V[�+ܒE#@�z$��þ0	���Z���k��V5��[�k[�$\Zܪ�"��ϰ���,c8q�q��.����4�=2�R;��kwM�͆;Q�t�f\��V�Vt���n4��t�z��D'���skEa*�`ɐd��_O��A���+� �q�#�o5
�I�g}�Y�x��}�=�� ��#�ɥ.��|RgWK'�.�t%�O8��[E�:R�x�Ȩ�뽯.S�.��4�=Zm���6O¬%�Tt%�a��ƙ��R.�K1��}�(x5	O�'�Rf�ŧ]-W��C�9����g(�������Ky�m��y�,�q\o�[�Y���&�6��P�R@Y�:}Dg)�?�C�SG��Eg��fLqs `Z�Wn���A�ܑᲯ�qíGG$B����f���`40	����t�CI���� c�G?g"�\���<�Snm�:9�8�CMT+d�s��

�� 3��Qݗ�G6=��AW�)��XG�#�L�r��p ���An���Yz!�hv������'�R[1�5�_7#jRac(�1�Pζ[����R���t� =@�X(���K+�dJ۱���隧���LO	�JK�N:e<�(��6=7+� �S���*!��\ܷ���wK������S,��2�n!�O���C�s�mm3�G�"���%�H5�����'�=PB�,�lF������@�f�^�O
[d##`*<.Z�p`��x�r���xC(���2f���R�`X�~�������k������z��L�������ڈ�u�L��@��>�a�ʖ��1z����5�:�i�� �E�l(d�)���i�D9ͻ��H	�H�)�R�zS&e;VC1�,s��71`��q���@�k�&09�_���OD�
1 $=�\=��=C����� }���Y�<[��E���ˑ���t\�_�xc�g�a2�V�y�jvSxW�|]��̚�M,���_���M��wp�5�YRl��ԃ��w��Ϯ���8���>8Z3��я��L���s#�5�$��š�z!���=Z����#��oZ�\P�V�V��<x�@&/p�Dv����,��z�H[�K�!�)t㳈�V��s���Li2��"}��P����)"XqcK�o�z��Z�+�h������l~��=|�*��xǲZ.�U�ϱQ��P�+����t��t,�d|7;8�5KP���-]�}N�Ȗ���O��ܯ���':���	C{S�?��:ه`غ���9���`����>�Ț��C��a �l	�vG�ɀ�p��ڮj�ǃq׊��u'��hu'������1�C]�����	/��ɻ��5�9�	2��[Z*|D�A�9+}�����ځ˿ξ�D�C��sr�3���s��l�A=F��j$6E!r��q)1'-0'�+�3[�Ξ�k
�މ��a���"!��v����@�[�I�79

"4[5َ����M.���(�d�X�&`Y��:���C�O�_*���3�U~��Xci���}�<fV�M�Pq~��p�������T/p�,���^�	��[����1�%���3j���O굎������Q8[Q���L@�� `
�4Ng�5�y��������N=渉TCĘ��n��t=5��%��kOfQ�(l��?1�������K;�'T��h8
|������O@q�^+�5b2�|Ň5"c�x����~���W���8|���d���ýGo���T� �۪�l�w��\��#1L�J!�2�O��冦?�ϓ ꭼp�.��� /���B�%M-��*;��wmmL�3���P��e�����ڮ����o-<�:D[07��Gj�=�UV�%Oo�_�V9mb�[�=D�jC��*�N	�2E3�>X�!�_�Ĳ`M=�) A��b��
~�b�.ٍ�K������ш���@A���]o��~1�",���y2T��N�Ғ}1�_�!@�`���=%�\
c�Z�$r���*��A䧯f�3d��'dX���C;)!
��5Y�ڍ�#o��b�d�7�TM�RM+��Z�QF�r�_љ�k�g���~N|b� �6��$j.�
����=�����8�*�E�:�0uH�N���!�-C(�o$aX���K��JU	�sф���e_r�yI�"$�R�}��PW�����:�lĝS���A���l���"���W�p� q
�@����F\ȴ9-�huR�oLj)��ݭI*�ߜ:�VUtSnJ�x�Q{���w������Q;�
wS�҂ǵ�����j�ǭ�'bZ�L<�{�4���^��x�����Q9D������s���-���b8�z]cj������sXzT;�_̑�*�8�,�]�a����ka%
�VX"c�4�߳��U$>/�ӡ��}�����4U�)֯��d'gB���C=nh�����olN"Q��^8g2)��7�5}����xd�͑�e����%[�v�!s�%��u�B����@,�j�Z�����K����zYnMw��q=G�։ �_&��ϰ��+V��G��D�p0{!�[��ꖤS��qr*���I�$e(��s���5���&^>�4��r��{�I43C�v���U���Q��ߓ���}D���Q!'�\�\.�<���]H~���[��ވZ����X��|EW5��nX�)����f�,��ɗ�Rj�)9w����'���������-r!llK�"Qo�uq��1�Z��&��̧�s�ۏz!!���8Z�x�z�J����A���]���^K�]5EڻGqI�bZ�|����8m���̺K֎ZM�ax��&�X�iY��>���
p�:����wu���%iH�u�r�!sZ;h#D<m*~�=Y6�h����$�f$�3�oUt��-��#	��w
Z�O>��U���p�0m�Z�@&v����q�ƛ��d�j��,�=��hP�I"���ְY��p�S���c�ʣ�ŷ�6%���0B�N�FY�7#4w��wu	�C�➙[��M,,�}�ӷ%���R;��*����ɯr��=Ƨ�q����·,4�Oo������I�Lސ,m|r��(U�O�oyP}�����C�g1�����vMβFS����Z�d������+�yx��K2�+�Sڻ�\ޓn���y*�ej*zݾ�6z������j�pL�����t��"J˄�N,�[P�`u�0�:�)!}�MC�&!3�
+j�<��>��h�(H������*6�0_����-c�ʷ+ľB�dTza{��7+�:��l�u��i�:�8J����% >v�4s�Xb%�yd@� ���]o�~T�����H��ӷ��P�h�t}����u9���,6�Y(�M>�{u�~ncɘA�l�>V~�y_F�$,�>gtU�]��w�\yp�V���o#��*-}�?��3IY�(}|�bY��u�����kY�5n� ��?��V�
�K��c���P�߬[H4�S;�M�]��/8*��U"qtj���`��-X@阑Q�u�d��xѓ�����6c�	����*L�,���Vqx����E�,\��*F�5«�n�C�F��TC�wM��	\�&$3
:T��ei��TZ3Ũ����I��_{Wvӈ�p�5"�%B�l+�M߄baO�����D|6S��.� bC����̫D��Z��n��]�`�cD���)q�N@4]�K�w\���}#��ϼ��/�l@̾��z��fGӣ0�KcW}Z��XEGD�vF���W�P���*�pR�U�'��"cE`�#0��R<���˪��H횲�\ ��Ua��l��r�*]�i	��+V�oy�;����Kl�= ׮~MA�Ҿ�yzL%��M�	�������^uZ
vi7�JV�K��E�Q��G}5G2�����ǐ�GOX�J(N
 �Fէ��^���۞���!��� ��{�y�	\Q����M������5\̝X�P4 	��/ kӥp����-�P����S��+���է�������5�bw�@2��*��{�C�!`���8�����V�hl2�`�U��(��>����;Ӡ��>|�9�HدeC�VG��G��:X`A-) _�Ҿ�S ^d�&oY�e��)���*;Y��z�e�Y����?T�Kf̿4a{�x�Ȗ��%�zO#R���,�*���/�}O@�갛o2	>���dU=�6�qG���F��%>�������
]viJ�0:p$v��{�{����4pK����L�Yܲںሺfnl�!�Լ�l�+�6�/��<ˉ�{���H�	��_JF1(�{m(�\��i/zA1x6���NאEOiqg@�����3��KY���tK.`��Qb7�Uh��<��m��*��4&j�~�I�~s����Lϵ����\@ <��@�i�l�2�hS>f��9�3Eݺ�hw��<�7�ʅcGǺ
!�����ѡ��]�O7N�i$*�gҙx?O��)�7V�;�`G���V.����iƓ?۷���<'^��9�<�N�ȟ���Rr��~z���$�}аx��^A�L"����c{5;˩R���ʿ	
����c}�4���h?��]�HS?�gĄ&��s���-1�����և	��H!~�]����	jXC�c�=�����wg��9ʄ3 6JG�R�0sPk�So�I�y8nT�j���v�Ŷ��{%�m�#8W㺡P2��34�*}�Kc[nO�\Y�l���c���J���4�e2r�<B�ؒ��yf�t�+�+ٚ�O�|�ki`y1�X��ں�}-�v��YQ��g��|�K���Nsa�A�rW��
�H�4���ͼ�KDfΑ�1*�����Ԅ�LǪ�QG�!s�9d��I��JLj,9ǣ�m³��gw2� 0�"2QP�/��g�߿*	r�v������H´r"��1}u��,��b�f�0YߧU��h�̛����[�����Q��� �*0n!;�	�
�rE���_Е��y���<�.�9�����*�Pq�m&{l��βz3���T$.R�(�{�����6���5 ��s���@��D�d��	���t�k�l�.�[���㟨���9�;Y��EyE�O�b���r�mg�����O�5�p�+�q�K�KH����q�y'@�B�^m�ޮ�o�-���e4b��Va;���m]Ȱ�4Q��VV�pm��g'ѻg�8�`)}̆6��0���!k#�6�N�̂����5��s�ݕ�.=��A4�)_ #G��{hc�}�@�8�~�vf� �sF�x���J�oپe���$����LM�c�(1	1�ag��2��C����L�DJ�A��+@s҄p�tcz�����et�e�[�϶�oK��>l{�2�(W:cq2�׼��aĠS�?� M?O�SגҞ�$dK�8;�;�V�|a�7EP?���5�~��<[
;I[w�j�\]%!wy��"�`�߽i7u�4��F|w��)�3�Z6l\�D��t/��5���l��O��gzJ�D\���Ty��l<�7���´���
�Ǵ�'��ARM���ȫx�i���8!���c�˚���#��yꝾ��V����g��t�����"�p�s������L����ϵ*b��ȕ��J �QL�y��t�J�3\�e+�l��VZ��]P��7���/�5���T1��*p�c%oD.�����UO��Z��9����S�t`������sqA�7�[Ubd�Y�Ar䆂���@Kg�ML���A�&��!D*����e�bݓ'J4nw����::8h�	I���0�q=e�����; ��O��ut7ah��z�ػ+���f`�D�b�f�S+���p�!��6�Z6�i�
?��ѣ�w�g����E���ܲ��e۾l<�{��3Zj��en���<>X�2Q@���_2�NꥉY���u�#Y�1���J�a��V�s�GГ�B��h���jkݿl������XK>�m��a\��yBJ�������s�iA�Ñ]�F�_P,N������t"( s�N����ѤWka3-27|�N?i̩��xzc����ĺ��/K��݇XZI���.I�_�7�4v������
���� ���mU�t�ϳ|�����<cT�j��pB�ʭ�>������X�8�_`2�?
��KQ̼ `d	{OA�}
��&�oAϔǼ3�v���l����F-�;&0��$��=����C�~�:���B�߳���s���S���dh��f�Aح/���aO���o�O��nL����-�<{�eVƶ�J��N���i�{&�x�'�Ł������cŭW�?��n��O�?��1ÑH6�}�#�=�S��=���ΨS{Їܿ���6�{YN!�Y���=�eV�C/\P��V����y?�m�Kݘ��w~)�����z��Uܨ�b7�v�6�[@\K�L���J�,d*XJ�?=��\pި|I�(5�Ssco�A��H[�9�^c(��:=��7�3x_��������l,�������sDg��P�)X���˥p�;���1N�z�H�>���bw�(������A˨���@�D�^OVLԩ������J�͟w�3�|��)�zf��`iD��N�-�7������P�#��U��>IØ(I�
o���Y�(ğl$=��y�;�8�l��Wjj� 	�f4����$��>I`t��A
/�LRH��fY�[#�m�MP��� >>�泄�*9<y$v����_��w���
@: tS�Z��@=��	k
�8v�>�~� �C���Y�*_L-2?^�ܪl���y�${Z��I����h�ؐ��N0z{c����l��ʵ��Z+s+6r������(��&5�oG������t���қ�QD�8i��]j˛֜�|�~�@�J�e[��ɥ�	o�E��f�?��ȡ,9̽�	�6��Ӳ�tnvQ�d��Ѫw����Fa�������Q��C���OH���Y�J���+�*�:�h)C�K~����R_�n@3�$�Y�<M*�q7:���g��$h%���H=�W�*�e�e���+�v�t���@�6�!J"{��2�U�rGL3�G╿F����V�m��&J�#��GhQ,mBg1�T�H�̳ھ8�H�L�x��i�>V�������Ek�K����i���8���&�S�kMa#.r7��$ ����i/�����!H`ٟ�Y�$�A������z7�Z�Qǧ�+�#VH� ��ݕ��w����=}	b����#�!u���UXl�q3
��/�*�'��$���Z�� �+,uf�?�i��:�EA�z*6��^�Nʠ��zX���j����'(YI��վ�%>�<�?.���0gTz�?�]�g_�7�����Kݒ$Հ�������.����f��Zی8��H�5�,*�>u-�+�
/%��f��
��U��Lo�\����ܗ��@��S������$^T��Zx-����n����s+��f���K�֮ʢ�HSO>�^h��g�\�~	��difV������P�@���?%�2�r*�/� `>��"yF�{�#2��3�ռ�|�LY��|�!�To��a/��,�$��h~M�	=W�t�2:X�*_9�u2�Ο��h��ߓ��ux��nM���#�F�ʄ'l�Иb��4���3�P�V;�N?y��qX T�4���%1th�/6X��K����@Lj��#�x�.���yD4�#&���J[�����(�Na�����i��[�lbZ~�e;NaCj��=VS7��͟����e�5�#n�������\n��|s{7�J��3�E��C4�}`I�?�\_DZ���N��[G�ˎ����A�U�"È)���o	|��y��J��-���ȗT�#\6E{�׈I�Uì�{��2')k��CMdW$�٩��Em�ڦȤ��oH����z�T�i���o˚�Y҉��^�p���b���7t��t1�qU�f_e�2�w�)�,��b��%"]c�O�xܣ}8T�̲ԃQFʬ A��"��-�f|l�ƍa��7����gr�p�`�l3j��Q3x*-0"����/1#*ب�M�$}7����O���)�Ҽ�Ӓ�c����C�m�O���M��2�<i�K������g#��9e�@����λT�q�>*+mj1<��fS_�3��|rNW��>������SQ�r��/��UR>ڸ~��qoE?�1���u�)���8n�h���[���C�&�:Nc_y�9H4�C.OM��$���#5h���%��E��vp���`��]�7&�n�mp�v�U[�;�������m��e��l=Kg�"Ϸ���'k��읉��ڄ8����?�΋R�O�ff�v���}�_,�<�|�?�n���|��U����R��ŗM�LUv�;�6����)�|z:��W�����ꣴ8u�ʇa��^�yI�[��6g��B�j�Kǁ�6�C+[ĺME*wR�I3ү{���6�)6;��P�[�s��9tsO4��i(vv7̙��GX�� _�Q�S���)���x������:���e���v]<�s�hwt���Cw0�	�_�v"6���.��57S�uK�N�EݧI�l�`(}gE�������O�U䩽L��@�`ʤL\�� о%T^�������u>�V1-Iڥ�!;V����#����w��z��j��/��yV��أ�k�{�#�B��L��e�	�G��V:w/��O�iA]��L�Ri�,[;���i\޼ʐC��vJ�7}��#��N`Q�{0]C��$��� �� �3���y����s&����R�@��œZ�<�)-�nX�}�Fė�;A<#r��+�WʋŚ����o4Ґ^�����+�b �e��Q�N�������|��I"��X7�-.957d�6ʞI�hX�y�5�HBʙ�d(�(�;zY�� ���]��y���OѼL6n  1i��͎�ַ�#"��v��ǹ�?�o̿�M��m��*�͙���h$�[
'�jx��"�d��x�ֻ\�''FNKQ�*��y�<E�A�!=3������2�",#q˾Ϯ}�,�X�h)�If�z0GW�����k�Kӽb���SaB�)�p�}Hao>���h�[�cґ��Od�7yܑ���:���1����G/��� �Z�f�))�C��I5�;|��,��W5�ݧ��tL!����,���K����+�	�}��!���e�\g����h,�ۻ e�}���̓��h)��EK1�-�#�ͨ^fH\�!����Ӷz��CFA���H�lj����K�%fd(T[Om�,n��.���%��e��c���z�Ͱ�P)�ى����Fп���^~ی�ָ�G,ĝ9��]0��t�[j�/qS�,TT�|�`'���
d�����O�O'�G���R�hL!l�Y��&m�*�����<eX�ww����ޝ9�޴�7��pS-,�y�Gv)�\N�����-
֋1,,q��.� �!ƃ�߶���_�"���;tp�NP�iQ� PP��TY�6�	�)�l]�P�4�	e�̢C�H��<�NT��'B>���wI)}
?��Ťf�%���般Q�&�֋����酊��~Ah���c�"ި���x�ru!4���Z�R���O�Hv���U6�{<v���W/;����	�`����������)���y/��
�2�h&3�)2O�gR�[��#zO;au�3X�'j�Cܭv�7�x�g*�Tm~.������UΠ�=������tJ�B�{�ל�#�j�U��h>��6(QڙQY������:�T��I�/_�ꃋL����a�=��q������y�r���0Fz���G�)�
�D2]�;�ʐ�1�k����̛!+cs�,c����G��(ݱ�S27��L���v�YA9H�c�wWp��H}vo=tE#l��.55-񇓋��U�<������{�@����� �G�E舿�A��`�t�]���[��h�	sΫa���S���e�h�x�I�=���B�W���f�!ylK�oR��p>����*M��(B��^�"ĕW�ީ�sw��/�+�ʮ��L7˦+k	m
�0��).�5��i<x1��K�F�v�!��DF\�.�-hT��f���ȒAF����g'3��֚ۊ�*�j�5��ٗ�*���1�m�c�JBb�-�Ƶ���D)��NK@�;�>�[Oq{kO�	�_�('�
���Jtʤv�~���ٓ��}i�zI���}w�K�f�
��a�2�曑4Δ��_��=�&�C��($o�����Y�FT�2�&�{dnaN�ت��VW�\� ҋ����()^$���Z�%���M��i4>���`[l*�R�]�r�����ɮ�$����OTc���=;9BM�]>��(Aܯb�{v���$��)'�0�rh$�E$d��b#E�H�{�p&��~8K΍kX�7���ЈF�#��c�X�}���P=!A�xKnE�<��_����e� ��=����B�y���ZA}��J�jPF����,
��U/�f,���J�ܦ'+0��W�Q<�G� �]��н8��cճ�i����k���G����~K��-G��h�iv���}F_�	ׅ���G�y�њs��rX�v��l��H�NV����z�D�t0�����H8��T13옯��6��c$r�(��ڨ*!'eMPx[M/��6�wV�LA�_��E�콽5_bH~i��y�݊��ܩ��=�n��ׅ�Y L��^p�U��q�K{M��í׊7y�Nuq��äI�@�go�)��J�^t.qF�R����S���'R6�"���5�\���ΑS���x0�/�L� )�zu?�B�*$?� \Tڙ71�^7#��D�2��SC�:v
aD&���5�s�#<_5�!��p��L�|���F+��C˦D);�r��ܖ�\�Ψ*��7�z�3�t�&\0j�?�����r$��������_5m���K����xP"ٴ����8�v��W`& "̦��,cC���r�:�JDy�P�K��A8}E��h	0:�?���o�0�!�!��/%k�@j�h���%Ҷ�7(�J���}��М$�!R��b���;&6;|�-q��'F�&@!�*#5�����ͣAv�p���)4�P�@���djE
IJ�k�?є|�M���[�w��/�p��҆���n���s����N�?M��\@�]N0FB9�i��pC;��P�_V�*��,�^y��;��p̸����0��D�8�uJ]�����{�/ӹ	�$�4�Y�ȃ��m��'n����{U�o9(؟nS#ޝ�NU��ڊa{o6ʋ~��ۥ>��m��o��o�t�A� !�V�ap�48dl��8.U��ŕ��ta���/f�s���Nw��B�`Д��;�y�rBh�w�I.�;�]�V�&w��D�̺gq�	�D`�G���M�����:@���0n�Lc���xkXɜ`�p}R�Oqg�H�9"a�_���Uɇ��݀M��o/߳NP�����,E��
F�1h���	ͳ�d/���3$�0��f��)X�I
��Ms}���8C��JѺ��o����du�r͏��ϑ=��˙��Q�7<N�'H�z2���oV�K\�^X�W������X�4�Qm��y���h����\,<��0{1�i�E��+�xTdS�]e�FE"��-��QrМ��ƃS���L�}O�ۼ�w�bA��Ɯ/��E��<�F������up��=�|e&�@(�X�k͘�MP���<�z���|B��0�N��?��q!h &��Jolm�(��Y2��55�D�9��T/H�e H��A�F'��p�	��n�|I&z��I��..�}b���ߙ�\�u#
et`L�NÿR�Dx�"D�B>��K�%ހ���(�"�c��M2�c6kff̗�bφ�X���fdj^���X�C���i���:��Hǭ`@*�!�9p����25G5��<L����+�^�g���{�	�%_�\G~�6*����7>��G�l�1���Yn/)��3e��߇Z��V3:#��R�q��S���-��ؓ)�0�����y��Et��1���Ƴ�شz-"�*��r&W� QMi��x���ú�� 2�U���?�#��cӕ8u�HgR�R���!g4��7·����h1|�(��j
�;�S 	�J���VTA�lQ�5d<3�.���0���,�醕ë����n��\!�����j
CG�/����]r���4o�f���O��{5��i��=�|�k��7��'�R��
H�FW�x����l�]o1XL���m5�kc�ӽfa�C���hż�}�wɿ�[EK�.��kA��v�9Ы丑Z��� ο�V�����Y`�Q[�/��O��R�1�e��3SB�/]hA�ǊΘ�Ą:|���g+ҋf�#zb�ƚ�wƺjTڵ�#E2J�y�b�;} �i��W�S0֫�qOS���=R-C# /�@���E�';�ו����N(X�kU��\A~��^S�ߙ�8_0;0U� �~���{;���Ÿٿ9��ɣ�y�>3���2�$h���oF֒���h�v?��&��n}�p��S�#�>Y\mp\��վJߴ}�Jgj�_N~�YX��P}REZ%7��Ѩ�_��V#��pi�4��9?@Z�k�مll��4�'��	�7j`.o��_X�[ل���#���a6���#�����6 �Nj���k�Ihwط	#�?���9��t#r��O� �ﳫ�N�����d��L�>
� ������;H��#��3�Fp����~��]��MrEc�A?�$�� �j�(j��t�� Q��(.��<vI�hD����Qc���$�m�T�q�(��|�{$\�X���ƺ��,���j�+^��	4x�f�!o���[E\�:B�\2�������D��	E�j�#�O�%�M�)˹�j\<|���7d�FWŘ��[�c��?�ߐ�O��4Xh"\f�7�.K��L�!M������gۨ���Lܧ�����Ed	eM�^z����'(�+7ϼ��51�q��M�_���I�4��#��О�⃸�+�z��
>JL�e��q���o尺KdxN)�^�?����8���W�=�e'A})&('�Xw#��l37a�����--뺛�!�X�f���3�pTX���<)�Ij;{w}��)�K��� T�_=�a�Q��<?���r�u��έ԰���Vv�H��s�K�'
��������RL1+�S������4ٷbQl
6x�p�@1}θ���''��X
d6l}Iuk��� ���n:��Xë"Z�_<����+r�O\���vmRư٥KKgyTu�l����'���ܦ��� ������*Ԝ6E�\̚��&=�T��rH�+ޛ SBߍ�0�FW�j��z����
)�9�2�JWY %

��H/jn���=EW���#d���h�yպ����n�cK�,7]�#� ��%Y*=�I\�x���,�[�I!֘kv��9m$�� ����ɧ�w(��E��U��#8Vm'fn��n���,P�׻+Un�T��a��}��-.�~���-�
8J� �[�n�ސ2a��<X`��7�G�Pi>(��𲔦F����8v�����R��V�q.���-	��۔�Z���I=(N�#K���_k0��_�o��Ҧ��?�m��%���o$���%i�k�sk�����%�02�8t@�*W[)�|0�� 0�q*G�r���2�g�:�`m�^�qYܴ���˃�#��߆*��tE}��������C��#n�R����sE3X��mѺ	�H�b=���R��k��)�5R�ӭ�1hМo�*���_�>l�I?�ѼCl/��U�f���~O����W7�M�doԦԥB�đ0��},f�c�O�&�!��M��c��1r��<�y�Im�S^�^�ۼ�;�����|��Ɍ�~����Bۥآ�+�_��a��LL�]R�Ewx=����`����_PU�Z�3�pJ�,'�G(̏���D.]���N����y+lo��C��ZC�˱ %E�:���O
Џ^�!�o*͔#;����(cT���CI�R2�o���=
ǣ���ly����M*��%���Fo4Xgt��{��'!F��&�'�k	���˅k*�<R��I��&�cc�>wq{5����V!/;w۵joie����9����Y����A�R���[S����ho]a7������r��m�6Kv&X7Qϥ��D��qi�m��:Ү~$�V�M�&��U�1��
&b���~�MR���P��:�8�����bӤ�:������Qj�\f%O����@��VK��t3�����:my��[��u�t���q�$�k�z��i������	i��� ��Ia��*���C���z��{c��I����v4�1���<O�z-��!�Őm7U�X��)��Q�&��L������ng�͖�d�g�%�T�bΒ�cO��5��)ҵ%��SP�r�q"UY���QT8L�#��kdQv;�KC/��uw�ғ!9���Ti�j��g��"���A����w�bY��:��`6� �l;r*9�ێ����b�SN���g^b��c��`>G�7]���" �&�	R��}%�d�f�s���x��o������7��'KP� �����rFB����v�%[��2*L�5	B;��,�o���*U~�����vQ���P��Q�59���3,B�}@�������f��q7r�$�Re���Ĵ^��{���@
ٿ+1-k�;"�ĸB���4�3��S�[*����ךI�5�V��r:Ԟ��Sh�֚BtE>��;����C��8x-ǩ�ܭ�6��vN+r�"�E�P�T߿�Az\ϕƫ�fJ�)-��R��FOG�e�h�.la<��agJ��}6a1;��1��i&kD�sE��(���M���|٪ci��񗡽耏�}��,];@�B~U�H����$�p%�g?n����t�-�M��<I<sk�®NC`U�/n1l͐]���B�b�q�%d� Ȩc����MFVAM��3W_<�lZ��R4:Lx��"�P݂Ɠ��B^�5����,�dW���A��3Km5v5�~Y4vE3��G|��1�$1�������e23�x;�f>��&R��@'���f���f���>�XHh���bs�Q��e����/sCy{�N�u�Rk8 |��W�*\fCP�(�:hk7�N�E�u�R�+; �ՌP,bޝ��l ��2�O��QE@ec�@#�?��ſ�F,�0��R��_c� ��:d/�^��K��c�4�񻕬֕󐑿s�]4�VSU��D��3hǥ�:jİ�sť9��4�����:��x����W��J�("�ݿ���6��E��[�����Ua��R�;[%A�9���L�q�.9K���Z5s�����ugɃ�@{����'��-τ�Ć���f0�fe}�,�ȧ���E�Y5(�I��WV��exK�����.fq[�2ү3��[�G��?��:w�U���vm4���qb�a+�Wɢ����M3�]��v�6�4�^(E6i?Y[�u��]�;��"_�*�������00e>�jń6B@nv~�0m"�h�O�<>�@�=d��8/�������nMXk��|�
_�YҴ� X�5��\�Ι��O��0x�$Jh��ө咶d �FH��%����~7���h��ƕ.ؓ'dR���>�bCV2~-"��@M!IQ�	�o�r�yG9Ս<�E�eLKs�N�h�hHW|���Ct�F��@�_J
��$O@3���I�.��z���#$��4W��KWz�:�	i���y�o�W��ec��]�!Ig�N)��"��Bt�88����,�nC<���`3���	�4���b�X���Zj�����I邏�/M�n�|��K)�����Y�챉	bM8[FїFL�Fċ!i��k�,�������nq���;p��7��c���E$+)��3�<^ȕ�\��s�)�Џ�/5\��46��u޶
i�]���yN[��2""��]��n߼����r�\Fx!�i���:��&l�]�u8S)��+jv�Z){ZKyQ�O��:��4)�==�����T�����[�aMN;%s�F�;��r���B�_�k}}��թiBb�m��V��!q�j���
lj�٬�眔L;dBi�p#m��-�&8� �
�ǩGb�n?�+���c�sD�'0ÊeO�|��)!p%�����ǚ�<k��hŭ�n��``-?Au���1�0_H��Iz^����޺��y���:=�/��ݨ!��	��٩_hV�1�W�i�L{���,��*�?*��FKCW�������Q�;A+�F�qȖ�)t�l�=D!K��j50����R���4��nf�H^̘�&��g�U�f
���:�����Z-A��F����ܨ�
�a�vT@r���e�������!_��DԱ�S,�ژv�����h��#[�O����(�Glz������ç��.I����	�GD��3�M*\=��u�;��n0�R�SP2���UP�x�/NS뎣F��(��a��f��0 ������N���9�N;�?:��V6<�W����}�6~I\b�T�ȪU����I*8�7v�B��%z�qܦ���6h,4�Zuf����ɷ���-�aL���w��u�Zlz��E���C <��ęG+�`J��~�q{^�#-+�E�P\�3ʾ�S��'ˣ��F�5��Z&9�,!�Ҹ�O��n�7������6����:&�Ha�9(�Wn'���B���U�ԅ*/�L.�/���o}�L+�yQ�;3O�����[��f����)KAnD''������m6�&6�ۦ��\���·~��g=q���<l�LF�-�a'�Zl��t����H�P�~��"��%����%��L�ɽ���k|\�,��x�}�Kg��6]|o��)Q�l�t5�8X��~@�(�)�MY�s讎w�=M�����}G��x�G(�2���έ��Dг��Iaw@��טH��������N���F����*�G�t��y�=�y�>T;{�y���An>���4�Z���B�b�lJ~�s�.z���>�E4	��\�R.9Er鮳;^ca�g�'��5Za<��S	�x�.�w��k�N{��z7Wh�ܧjD��6R9�"�!�N��1ty��y,��1�	��q{o��ĊO:�ޭ֛�ڌ\�#\Ot:Z�|��6�8�J�����9����Y]|��<��eh�4�^�-����`/�'��1D�_���B��\��9���]�_�"�y�t�����@VxP;s�X�3[ԣ���Ƴ�?]�SZx�e��p^�6�s��� ��~����~z����G�0�ls��f��38W�(�s�
ޤ�����`��H��eo9�S�.�8�=�\�wČ��P՟*�~�v=�L�F���-�W83�C\�$��0�,b��\���&��E����n�{�l�+��Z�~ވ�y��a�դ~YWz����K'��䦍$����G�A����_�˺�C�X���6$Ëh�0�P˩���^/���`��*�d18�	�i	��u��Oks���~t[��]���h}Dz�0�[�"�_Px/�{���B9�65 g��"z�-�ҟ�w�0�0����ͯ"�����a�Xw��gA����w6ox'�*f	=�[��s������*r���w�r��c�����I^J������1Cn���\��yK){0�S�H�Qs�.�d����[<�Z/�&A�7�l�w��֥�l ZM�~ �Wb*�ö�R0Na��O���6L���!u�f���w ��\s�l
�0he*�NC��=gWGg��%>��r獅g'��A�	p�����O(�V'#6��wɩ��.�����r�fɋk��Z���-�v�WG��u���N�d1Y4׌q��s��6--�n%jc���x?��Ͱ�9�!��0"Bn��ܗm{��J���e�qg+сL��<�;��Sx�S��43o�r�ݎ4b��]5��̖�o7�f�6}6��9�omACAz6h�D��̀%=5�-���x�X�.?�6��O��9 ZwD�k����Hq[�O��Q?��KN�T�n�Nx��W�lF�EG(���zPy:�	�f�E�1>��1����l�3j�R,q�_
�)�6�9 � �N��oo�l�n�9`+���
�ٷ����B`{ɺvu��w��܌I� �x#��X��ܟ<u4���c���B�喅�u�&p�����{)��n�b��@�t3)#��)�z����r�:���M�F9�����"x���Gi����5$��{��b�\	/ V�.��/&%����.7��w!�F�u��K���d(}.m�FqHHץ�|�����3x��x;��f:�u�fV��=��Ӆ�9�v�E�9(�٘F�H�:t�@!&�ZBlKF�(#�+���˅�b�OOτ�m�Ay�s�!�d�