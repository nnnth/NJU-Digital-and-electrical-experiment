��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��ϱE�e���0�
1��@�Գ�)�E"m����ް3	��[ms`���.�E�x��K�x��H@6�0���ܵ�n�a��rI�N�+0wѓ�U�BH�pd������u���� �L{�rwMOㄜ�K鮕짙4L�����Xǥϖ�QC�Ĥ��(Tϯ����V._泭�<����Y�C­����[��7�ܦe�'g(�#*	��q�N�0t/[���4f?9�)��`�hN�����2�(1���/N/1�9���Ts��K�I�⧮�K2�ࡹ�6$A����J@��m�v�w�e�m�yѦ\b��w��t��f��-�[�ݵ
�� Q�1��^㴔� �瓷��
���IѴ����#�I�L<�"����*�X�X�-a����@��r�M��F`�I��.^��ؓ�E!$������������ �c"��衤����%G�	ü�� V��WQ��Ria��3����Ç�Jud�8���s� u���
���3u��"�~o��U���M�$T;�.�[N����>̺ԕVڙ�.ˬ��Yy#��˗�C�@�ɨ����3�a�NZ�/�ZA��-FC��}5�����ܓJ��+5<�5��R׋C����jX�W ��/e�A4�z5	�Љ_�C���9�����A�ݺ) O�c]�\'Z����y`'!��C:��K|j��bk (ʖE�&�7��[di���R�b[���;��?�4U���[&�0�dԮKU�!6�7¸���A�g`���`�l.���H�����?��E���5���m�+nfGI�"h1����Z�]�<�@��"H�B/,yT�b�����J�P��-!����p������E�V�?�^0�Y�oB�
q-y}��}���ߨq���y�X�d[>ŗ *Ps��fC5.�j��[�9鍑��J>�ިzGqYk�����N�B��#��& }M��k��8h��ɉR�N�&?���} �$:�)qECy��X����M����5��cR;/h��H���dp�\�^�f���q����g����+�vߚ�{�y��N��7�IS]t!�H=C{��<2�t��*~T
�
3��XM��')e)��JS�Q�@�6gJn/�F/:��DS�l���;�ޓ�����Q�.�y=աj׈й������j�^ �#;c*[)'f￱�̾��G�+I5� U�T���70�㆏^�=���Z`���&0��E��~��銢}��~F�K���L�RZ$�ΧD�.�9ya��Z��S��䣬���SC҄B��4�@X��*��\��5���$�m��F�i���>'W]
j�Ma\, m���������	���U�ol�2⽂�텏L�33e�+�AF���c(�C��N ���/��ZS1�!��p��-����L&�s��֮�c
V��ه�
+}��݉�:�������i�Sȴ�����^F�
vAZ������,��n+{�7� �7�0��^!��F���4l���CZ�ŧ��ӝ
�,�"73��i=��t��)�C_��<����<�6����O���0h�O��k=|K�!/ށBJ��R1���.��*^Iگ�]�ؙu<�� ���՘�N��9PH�h�'ջM��-7p���l����w�W"�S	�*��0ՠy/�p��f��^�]� �N��)�'�[������kaJ>x5_�[���gQ:��|�ڥ����<�R�ݲ�Jf�+�)�9Џ�6z����v���C%�aY��g9��hQ0}g˛/e&��G�1稚T���xf�)
�MǑ g8Po��.�T�I�q�w0�L�ٮ\'(�@���B���Q��P+*W��8���"�W�ב����= �ǃ��V#��c�wP��ԋ���j�U LH�؛�׬�����_��(7�H���xR}.Q��!����OYS���i��Ն�**��oj��$ߏw�m�� ��dӹ�!/#=��9	��`�}�e���!i��+��5fƂ�/�f7�VK�J����ȝJ׽��48$��������`ȹ�!�92�F�����$�0[")���JM����G���HJa�ovM���¶�������*����s�\�]0XB�����1��f�e�O(�G٭莻5��N\�p�Q%��lI�S����bw��-�6� �,�ā��7��ET�ف��Jw[;7�n�c`1sx�Ygu��n�W�4������V��S|I2��d[{hU���{q�2b�C���C����_��r������:z��>�����ao���T-e;GP���>�M��&����K�� Y������ǫtl��U!�Q��y1����X��5�z%�W���9�vap�+s��n~�4j0@�i���D���י�'�k��̌��)���N�tX�q��u$�P9\��H�������m7��9� �t�.*t�,�S0��闎��׶����Hs�*���1�2�q��_�3&�:!*���Ns aX��}5R�%#�Hp6O�q�q�`�hHɓ�<�g�m���G�JV��'�ِ6}u�t.RN���/�[I�wv{�����`��Z��z�J�;k�/c�zWҹ^�^G�(t�*��}l��s�1Ja~���Wmm���~(��
s��yyV�E�9#%�����$=W�f�.t�c�w$�i�a�۹��g4]�V�1|��Z��ߎ��:03����hP� �r�:G�7"?2��t��{-w[t����]DWt�ʭgF�o��Y�trl�N���2�*�|:��݅�]���G�A�86=R��z݀$�nQ*�'�y���X)A�7ȏ�y��npɸ[J�J��]�S�ش���9m���H�'6xt��,�?��-&���婧~7̜���*p} 5r�1��*��
%I������3K��wŇ�zj8�u�%�׉	%�z5��#'Q��5���SvV���d���-B��y�ɼ��ѱ"�i�|>��M�T�Z%��SM#�Ы���r;�mMOh��)�^Y��(�[	(����ݙF9X��]0dɕ��?ȿ�;��.�cv�}U�t�W�i���5���&^�\�O�L�h��	9��z����w�D8��+����+<��� �Z����!�2ǆ�����V�^�?Y]99G�������=W��wIo��g��-��b��%d)H�]�C�
��O��Q ��3����)!�i	FI�h7��5P�����?��|ro-����-5�ħ���f�=@�K�t)�]F�Ja��xy��n�Q�W��H�A-.����H�;W%0 ��_��dbIs��+�fq�S~ �ɰҘ�ƩnN0�B�~��˓e�^���݈�˛�3�"n,ٶ�9-���e�{:.��}�u4�X~�-��b}
��f�y�V��7?�Ĥyl�Zs�ʟ����q��mq<=�?����3iU ��?�Kj5fGK�De�w��q�
�gt9�${	�q1�S���)���a=�6�l�c�B��4<^�}ZP�U^�Ȫ~Пl���[Z��j#>�=�e{�#$VU�$����gȉ6��|�S��p�~@�/El6�hƗb�KbK�i�e=�6������>9�2��]_��7�։پ{�W;.�Q��0��OÄQ��W�5@�����S�*�������ؼKa]��8w�0�K�.��xNč�M }J��)��R�������X��H��(�j��4�%����r�4�e]M�B��N:I�����D��K4�/ذ7�x���g/6C�4�ԟ���Ё3���K�mp;��D��~�!��,�s��J�!͉���q*"�U|����A3WĿ�H� ���6x��#��$�a;3��yp�Q33E�Ł���lKq���3aw�":�^�ć]��\����zq;�a���+�N��#3�#q���ܯpJ�EF9ޱ�S�"Mpn��>��q��ƎAp�M�n�tY;%��:����e��*����Q*+(Efs�p�\�R��-�ƶ_E����+�C��r3DN�xX�����CG<"c�^�Ǵ����P����3�h�}����hf@�M����zL��2؎��c����Yj��rA^e�����:�ªH�4X��ݢ�9������.���K�����K�hI'��U~�\�"X�@Vf���?\#��c���k\>�̛K3�ҡ��E��gF�r�Wu�7�����@_7�C�'tc���=[NF!*�_t�<Z��N�k����d̚#͎'�~ȑml>ɸ�Z����KNDc�0������DG�Yp�J�@>:	�Q4�"Dsg�m����"0����TҐ�	C��f\��P9�\���r纋�ÅT;���|�4E)���rs}r�,�>���M �Y��m���N]�'ŮBX���XH����N3
��&�W���ȼ��r(z���]�-��C��>E�齉fy�`ݶ0��*D��`{����>Ӌ�4GkQ4W�Q�1�ӂ��MLou�d4+k�i��#��)Mb���Q�M�8�=|vQ�hy*/�Kjr�ջX������Câ��O5��X�7s�������i��rHĤJ����������t�0�K��8|V�u%N��Hzq=�i痃��G��G�H!�ڸ/��-��3m�t�� �Ud�������y�T��Ѻ���(������2_i�gsɓ�gR��	�kW5:�|&�*)AoČz����9M�����9�<�V�j!����}e�ZXX$:=]�9e����s.�^vvx:Q�
z���Oަ��W���c&�� ��"H�Q�	?�6��K�Z��77+�n	�a��K)A�$�O삨��L-��6kY�D(Q[4�����@\M�_���j��Mm��V%� ���ad	q��x21�QR/�X�q���J]+?�5ETFz���k.�kn#�M���٦>xn2��֫W��k���:u�i͙d)m0�~%�+Ln��� 9��iD���:9;��i�ͥA?i��Ӹ
��?�۬7�8� �h�E	cn�#l�JIf�D#�����*�`Ϡ�6(�]Qx��N &/�"�}�m^CL5b��z�����]<]�C}�/�#�Ps��e��E���F��f��T���	A"E/���A�|����/XBL4��#�P�Z�-W�k��Z����X��ЊW-�l�P�Շ��LU�x ��4�����*��T�A�H����~�X�.��ڲ��W,>x�q>2�i��d����f��Wm�f��P�<P����d��ç�����^6	"�Y_jS��K��R������q�=��*�
�x9��B�H4���{0g.�5�ړU i��Z�d@�7���i,�J���#�d<S�4eSH [�;��)�xh�g)���I�'����];LZ���E0���
s��B��6��:���,���*�Q�'�Z�c�F�bro�?��L���CBdv���:̿�u�ڲ$b�[p6Ps�G����N�X����%W,$%��JVwr���.�@��{@���W`�$�LEX�͞x��������e{�&X?1,G�n��� T���
�[˛FpXT[���7r�XM�������|��$�Q��}�E�Z�򳞧�H�yk�|K}L����?dO^���E޶$�b�4��D��.����������P�o���/�3V�0��,e�C�e�X�J�����H�p�#�p^	<�m>z$�����B��1��_��׏a�o0�m��ɖa���/���v���.n,�Ķnw�H��5�/j$K��,���I�����'ɠ��qF;	��Ϙ�1�.�M�bnVx�H���^'-�czw0G�0��N�]闂���D�GRW���4:��|�Ufތ˄���i=[N��F|��pԢ���-��JOY�ו����f�;�g�@�}%���R3�C�ᤄgr\��i�x������_�c�ƖAfs�Œ��y�'�\��E�#V�=cr�ak��B@���
5Z�QJ�b���8��GI�f:��g��c�i��5*����-� gX�];��j��mg�=�,*���Z����%%�&h�_X��B��-.�S�����u'�Y�BXA��kE��[|n�5R���z��H�;_ޠ�ߠ�VǶ��&_���OS��چ��d�Lq�?.'��?6�<1�Zۧ��ғ������m1�n���pㆹ�,��X�{,X}\�Ij�����/�dr	�X�Up������jY�;�NC��wgVl,ݔz�dgl��]g$Bi�w���^O͟�f�?pNO(���b4}bO� d��]:�����q8LF�hZvg�j�
�yq��vSv����!f�Y,S��l�M�W�H��Q���P�K�]�mL�!�=���՗~S��ls ������l�NP֕�j�!�_y�U��
��>�g����o^E���.�n|�:9@͉70��?"�s<u���K�v[����Ozf/*�S��B�]Q��ߞ%Nh���`KP���F2��>�(�jI��_I�
�x�I �������G���C4��&���{���^פ}sxD˭K�(�!�o؍<��4��M�-.$ ��'�ǪƧ�)QS�������mK��E�%4`�/6#�+r��̽��@*��X;����_�H�x�CC���W�@`�7�hԾ���2�1WC:��3!>9��Igjg�T�#w�MK�S|���X>�~Ԟ����^�c��I�+��f��q�Rsŉv��>���E2���ȵY�BA�Ȇ�'�e1i���!b6?W��T��cҹ ��z{���q$>Y=�P��EW���+��%&E&�fglO�.�IA�j����]ŏ<����QjH�W�A
�q
�R���R`Q��;�����ʰ���g�t��(I����yл��C��o��Ps }�}�Qp�� q�d�o�V�0�yU���8�c���~i�K=����oh�lt�L)�<��� 7�B�x�(=q!�����g�h�<���1��v��qpΛ$zJ��r�ɑ#��BE��Y� ~�I�lo���4�87��.�@a$J�pj��䛾����*F8G,ݸ㞢�����a����ϊ�ŀ���|�N� >y�,�/_����>B͜6�Ҍ׈U�a�xJ���U��<`� +s�w�t'�j�JZ��A��B>κA�G3���	�d�]��t����F]��}�e�y�U�� 7��������v�o��:���l��tf�AO�n�}�i��W\�E��2�~C���s�1���J�����E��̡�Y1c����K�A���lm�O!�:)H&~K>r-�t\Д���W\�T��l��f��;̓�<�_�z?e�Cw+���ܯ�I@dNe3�5*;��"�t���q����u��"�`[�%G_4��P^;�: ,�(I-s��.-�:<�%�|�}��[C�}�#0�v)�؟7:5��Xsٌdl�ŏPF�;���.��`��B�mC���k"d�3U�����9���hA��(����(Qa���UL��_�{eX'����e�n純j��0�M/"��|tE���A��UW��
+�ٽ?�\�a���4|�Ӝ�Yq��GlH�a3]�s��<!U9��Bd^�V�T%@����K����N!3�>%���I���r���%m�A�q�>��@b�nV���T`�3,���Ρ7�F�i���V<��<h$[���Ϡ�)E�H�@�j�N���}yϭ��̠k��-�⤇x۰
ͫ�C��:B�^��u�	�T��Ri`Q�����v���-.X���(� BG
?���]��7rqf�nKk��49�c��4wPa���a��E8w^z�<ޭo��A3�ݩ>���Ύ����KP*�mS�17C6���I��i����H!	_4�_p7a��*ψ��kd�zf��$�|�Ǭ��I��Nq��j�H�C�o��S!IC����䍛�x���j܌�>��O�S�!$Q���"f�4L�~s�����p�6�&�cާ�`���3��C�Y>ݷ�?s��6�j�ß�	�R��s�)eEV���	,�c��
� iMS�PL��8O&������Ig��<s�fvG�*5	)�P������fw��z����A���B6r�!�cA]f��Y���3�-b����0�(�Xa)���,\ ��TP$�D�9�yŏ>g:��Z�x�`���d��]�����;�'h�AL��-Hz�>�sЕ�����Ȍ���� �� ��q���,z�'��D�~�,��L�F$8�q��p՟2�8�'_��[q�Aܯ����jQ�(�Y� �ݱ;s�Z�K��!��{}1]�4���W/PQ�Amݒ_M�ި��s����_����Z��"�ߩ_���٪�fV�
��ru��V�<&6:�e�
G��WS'��Y�O�j����$��맓O层��yW:Y���8/�N��_�^�Ac�P�[0�7(�����Re��X}�BA���tr��/ɗ���� T	�s���!A	�mh��6|�d�آ{���g��
�I���9�f��������;��
`#Ӕ��tO�2�*�d*<��ƻ� ���'��l� W	ob�F�I�+*#�2��G�-�G�Qk�fN��Wk��8���4Jb)�+=��9N�f	��i�@Pi�/��t��{��NI�?�ri߆aC5�<��t��Gd�
�˽��q�;K!�=����ZHg`x�~��w/l:ՇyN����ebd5���L��s0�lE�6	��)��|�Z�1p�������pa�e���9%���C��.�~����j����ڐ�Iܤ�mv��	�TC �a)_ʻ�����|�H�Z�H��6���=�A��+�c���B�����n��v�g��$����J�"w�嶗s鍰d�%Ƹ�%�M���Ц�V�1��RNek�r��Wd��8���qc>?>�5t��O��5���&'�e�*8A±p.�7��K;�'��߭��>�ް�1ڶG�ƾ�l����|Ĵ��\�e�C6����`)������Hl7Q\K��-aK��J�����1�-8��Jk]
p:j�'D�M�3Р�GR��q�k�����G|��軛���#�E���G�m���;"΢D���6���b#��?&�/9�?�х�`M�i}Pcĵ|���u.�X�~n���*N�R}�P�A6l�<GO�̇���m1>������/3.���EU"&���v�)�k�Y�_ֽ�|O��㚏�U�#�dT#p����ƱN�d��G8��V�@$�w�Y��{;)hYWC��#6Zcd��Ƃ���p������!ED��Q�7��a�A"#͚߮X1���b�gp�ߑ��da�%��I�o�o.0�渽�e�Cv����t;��'�W4���ލ��^}*�jm�m�|�>��;�CiF��%m���?#Z6�]�.������t�����-���?(��h9"�M-%�t)��?|5��W�W3�(����+�c��>�.��N��u$�Q2���ZB).��,�#,������)��9J ��Z��{Wk����������. ��&��w���:D��s7����?Q�|�u��~���!���A�!�,BgwG���w�7wU��T�*m/����D\���`Suly�@��۸�]��l
�دv���@��T��9��8�����){�eMN��bD������7���bڊ�z�o��<k�ZEi.�T���@�Pڏ�{��J�7����n$ⱍ�]7M]�l\ϭm�S~b��^�6��ɔ�[�1�M�ȋ�E�����J���:\�J�r�j���X0V����������^N�	��eM��|�'Ӥ+*tO ��&�xU�Zm\�PKE�V����|�L�49Z�i�vd��R���j�3�M`�7u�YR�${e��:$a<�XB+��0�"���+L�[8�Hǒ��2��T��bs	���-��_����:f��a���Z2������DX�K�4��/������L�e&�� -l�>�l۬Z��N~z���3�6FIB`t��-G/��%��+.�\��%��M��&j�P�b�:�=+a�k�:�z<��Y���Ӆ��b���
��ǕR���:��Iё��`*���r3�.�G�����VT���?��W:r�zȽ)K#�_�k����+��l�3���J,�h_ �O�i����N(�
M�Q쎟�2៴���<����Զ�E��Z�2ו9�S N��ȏn��⯰(?)3��}��=#3!�)=�S�att*�P�Jm���?�鴓�f� {2��;�pq���X�e$b`h#��M�-z�)q�`=~�Z�c�<U��@�"}�W��P3 Tb6���._�9����>J�sY��u��- �͠��Y�%���m���A��]<%�'բ6zڹ��^).[-g�am5�';�F��in3)	�9m_���O���h��g���a༒�lO���Sҙ+�R`!�-�ԓ��a�)��ȃ� �O�������$�0J_苂��?��@��)�3)뀆�2	�F�BoŃ �r��x�CAA\ ^�$$K����&�6�U��>��
Y�F܍5�v�k��,���I_@��H�	+]vL����*E�c��l���HKx�,�����}(�M���v���,��_ו���!��ȗn�����$����,�)�!�HPk8�&�D;�rG�
���~(�߭aުS�Ԩ�yR��
��Nࢗzmo��#,8�7�W���mqxc�������=�X��@%�^Ш�A�=jShJ)!����t:iR�� �n�O�8j�ք�d�{��Ͽ�	���� �8Ca���h�.0�ɟ-i��i ��[�J}}F#] g��K�5]�@(�������A��+�����>2*����B`�m�*��|��g4�$ȩ=�
mxR��]i�F�*�/��
���	�&�N߶�h�X�;:X���|�u;Q�H�,T�`�ł����}�����D-�0�����K:Wi�ϯ��Q�{�~���e���������u؄6'W ���S7�iT�DQ�������.���'��b��X����ۅ�h1�����No�A#e��R�9^�U��%�o;��A|9c���VyԊf�-���7�W6i#�lH�|�}�����,3]k`h� �`��g��K�:dK��pC���ko��\��?A@p��E�2��hh��j�zU(��2\
YM� ���-�"�9�j�3x�����Qu�D��.t�=y���`��[��<TUr���T��JR�d�jb؎ ��UسQ ��˸�t�|
'��� ��"PDW�E���~��Uu�*���P�Ĉg��p��"oJZf1��tS1��Iϡ�ǀ7��R�`Ց~8#���t���y�F��V�Д�hwa��CK�M������E��n�5�V�,R���?�@y�4�ĕHΉ`X3��3(=yb�Ƹ��«ƃ�-!��?�Yv��iG�H]�ѣA��j�fӇ�\���k�!=���JSOY�*#d'H�~�y�4��Ź����<����9���{��@DqhYu�3gU��`�|c=�	2X�g��ݾ��Z����"Qˤ�[s ��`�ݲ�EipiU���t�gDy�3HDUD{�2G��ܷ�ͱA�&d�3�ݼ��:�9��Gr�AŚ!T&�9T��q}���"����2y�@NN±]%�c};���,�$.Nk@{����^,�Z��rS������\�`ӓ�S�*/9���/�RϾmy7VX4���2N氯%�'V�����$��q�����K��e�(>|��� ��4Ǡ<�Tv�~�8[��y~�&P�����<5ƿ�zW�yZ+*����ۜ������&���T�Lu0Wr�|��w��@�W��'��b�M�jB�>°[5�(;� �92^{�'���?2Bh�lc8�w�.�r?a75�E���9��4������$.�M���b�V��Ch�3%�:�eI�[wH[iQB�pP��P������ʱb�|V�򈬁.�m�n6���P�Pq�
<���#�x)Nc~[���@�{�@0�k�@D����.ˊ��_�+8�bb݇��w1dvm��b~��X������r�����{�Q_���齾�o�+.�az�U%�I����bZ�)@Ffѓe4Y�U0s�@�PU�5M4Z���P�+����q<
��b����� �(�����}<qho�4�'9ʦt���OJ����g��P�Syv���,�:;"y���L
�Ubp��נ��S�O��=���/�H��-��4�<:�C%�A��z�Y�ZyM rR��i�-��j��ǖ9�|`��r��5��+��`f7�R���3 sff�1{�@Kz�i'K��3s�؇���C P��V�M2G�z�1�����s�p�feCH���5���*��M^d�y�Z���m�.=�(�6Wb�`�B�9i���Բҟ���FV�r�|�U�,�OlA3�B���=1-cޯ3��j�&�%�Y����[�6�~[�}	ܯN� ��!�W]��6`VYD �*kD�.8jbjY@�� 5�O��d��8á��>έ�,�5sX��ڊJ��a�1�=�pT�3ժ��߭���<�_�"u�s�,+/t�OTs����3ڴ�%|�&�j�dU�/V�7�c�Њ�)���yS�m�<îv�bR�λ�|��6�M�R���b�4��,�\t1��a�Mc0Yh��f�ϩ�f��/�`��*8���W�N�=��"@{��2�c�<�����M�:�3@o��|�ҔE����^���@�3n{%n��nO.!�BS|�h9�f��l�����_��n[��筬:h's��,hp�l�d_�Le�NK>�]��l�ӚD)�*,4��@w#h� ���<���ވO\hT5?�g�]��i��y���b���(����F=���f�o�������#2�/�����)���+�K�;���贅�C6�V��N.#�J�j��X=(�㈄��Ff-7N�OK!+����._)������YI���+���r2�#�$@�^����;܎Ŏ~�8R�/�^y��AM��,�t�Y�R`L��
|�5�&�mrT�O��(q� 8`�#G���?2>GGH��D��9�ugP�l;3R�k�^�j��Ym$Ǽ��,�~1a��g���6^K�u�XJ��u������l��5�&�7i������]�(�C̔�q]޶�5ux��t���/x,^���/�<]�ik"Lf�HM�ꎋ���L2�%�	���BU�v`uqj�Pe�!J��愴^��0�`"/��w�?j��y�)յQ뢰���D����<	��4<��{�d�4��mG��@�Y�s�B͢o�����L���,
��\�`����He$OB��� ��l)����6~�.:�H�#��b�������A��.�c�0��R5_�ǰ�njx_	���W��8�c����~�<��,e�x|ޫ�7:�
쿗 R/�%'lΟ�q�
��8��d� 0�H��S�Pw`��ʐz�Vl	��N`:��ӓƽQ煊�M�Χt4>�Y�:��_���YV,^�ر��9�H1A�y�]�~���=+CM��;e=%�u�g �~����2�Ǧ��&R�3�fh��P�Buޓn%��2��k��Z�ظ�	F�pPN��4(���ѥ$�Ɔ� �b[�P�D�.J�"S��4xq��+Y���;)��F��I��� �ٺ� kP�[�.k	E�c9�>��!pv�-�Yf*��}�{t�A� o��a!Ho�n����S�+�Q�՛5.���V3ڕT����V��;ƥ-|t\��o�E�&jO�m���K�M�8t���AC3Ҝ9OLJ�p~kowv@�����ez~�nb�~�0�����!�ܝ������ܤn���<�A��2����[���C�
��k�U_&X~$����x�d6��|hp��
�&�����`Y�ń.w�m�#�EoH��/5bW�G��*!1�b��65����pˇ��zrSE�)"��k��讀�;/Z��c��[��SCɛW��p�3� 	���H(?H^��m��>罠��T����>�y�` ��ken`j&Z�r�6��:j��َ��^�aZXm|��>��qX������X��|i�E���!��E�h۳5,��g���% JGp�n�O,/=�U޸�q���|�Y��"͛^�{����S���Uf�ݢ/���#���tѥ�quy>k� &Հ�FS�Z�� S~�>A���e��ҀA�;I$��3G=���;���K���+q�A���l������i�pz �f���d堿3��^�K���ۻ�XNJ]�����o�fT(���sD(o��\�+�6�!v԰��ĝ,�D��~끃j0����pZ�O��
��^l^9�O�����6+����Ӷ$�KC[�Z��/.xIi�����u0}E�F��6
�ھ���J�0r�S�S���p�r=3,u���,L����bc�w��B�G�`�G�L$�-�R0���']}4�M��D�Y���UT�,�\7N�;�ҝR��V>�p�x.��#�=Q��趰�W�Aj&�N�a�q�c�2��A6�c*?|~8�7����q��F���Iyۑvo/OT�@VZ�8��tK��u��ʃ�S/���p�d�)B�+���;Dz�_Y�T������o�O|ޭZ�"0g+���H�%�$l%sM����>�B��r�x�{�G)c>��L�Z��X�ᮟº ���2�g�g<�la��"���_lb"���d��4|�7��J�s�wKg��"v l�QI�����g3~����i&ʮ�q�b�%��kxVq�;�OiV��1ڕS�N���36P��Ȫ����h ���`�`[� ]���G�F���o��:�/=����t*J�A2��n��w��D,׬�2;~P~�B�b�tW�s.�Z��1kC�ʀ1sZ�f_:2��2ҁp�o��{{M�B�wӄ&�����.8W��9A;XR݅��G^���W�:R0�������0kSXhqŹ]�u��X���h���Y���T��uْ)w���˃��'�H+ER��Z����F��N׏���'�b�X���tͯV��4c���7hK�)0GT�L=	��(�o>乷�B�����S ե�5Σ�+%r�T	�(��5�+��¤=��#�5{J5�+�z�	D~H��MK���a�ʤE��h���̟�ɆWkgX$}�����ػ�-T
�q��1��Mx_#��`����?�ٯ��h�_{M�@��~�I��Bvg�u���_�V��q������>�W���}H��	y1Q��|�6ӄT��C�8i5�"�]�S7��]�$��oq�0������O��G���Ў��i�*���l����S�)=�ϒ0;�bM�Q�%���{��1�[\�-���`��k!���)4G�;��[	 aC93*�a-xW���ɡzԭhp	Uf���]C�N+���t���஍@�D>��sz��~�:���%ǎ�·,
=���!�E$���;)�z<���f=��-���w	:����WЎ_��G]���}�g� ���ۺ��hO'Z^���"�H�[��i^�"y��
�Y������B�%r~m�����=j��z�IRAצ�l�un/����.�$"q�{��������\��P� ��߳Kŷ5B��2��m�'��<�Л��s�c��ロaѡ$��w�Qy������,7�=&9���^I���ӮV���g���w�@o���Eĺ��t|71��?���$2�J�٪"ܠw�� �`��zg�g�wLe�{��_
{���:��^�2fz�{qq���������f� t�z�5�:��o�&`F��,��2PvQaX����>s�Y���u�}ኅ�2lȢ�DB&�������.<3��\��˦�X*G�TH���b<�s�k}���(���bWP��B��i���������,u0�ꍰ�r�e&V�Z�^�:;�R+���]�m6>�$	�\�*����3�������S�W�Q�d�s,GLGy^�Dw/PM�hRE�b~�������s]��8��ZXO�^Z��n}�\)��W�k?�����7�
� |�x�����o�+\ÔJ�xZ�J���ƇOQf
->
����i�GΜ1�2%+D�-B�K��Q����]Bޛ�w����
�Z�ˤ�p��mI��r)>^���旋̺M�;Jc��Z
!:�l ��Om`p��|�đ/�ՊfdT�y��P2�^;����>7��4.VA�G��r�k+ckP���CQ���+��+�)�I�(#$�S�l��~�Tf��;t�ܼ=Y\�x�*wj��kC~Q��r���I��a�X����c]J7w�8��*��n�l-�����/!�$�a�ٸ��IO����x�B�kI+-�$�֚y�i���LG.+O�?)/�@��X�V�Kb��"N�r�p}�h��iu}kP����Q78/�'C��� �Cg�d� ���Q}cҕJ@ �D�˙Є��+/"�7� �1���ӿ�lh{G��%kTk-��l����n��������:n���l�c��?����?#P���*q7��/�x~e�kg.�17i9w<I �a�DO���T�l9�2Ã,L|SJ��e�7���!V'm�~+"�ݸ���-R�LJ�������Ѫdf�'�
��~5�V��5���/1��rg2
]��'���f�~2�c�ZX���,����;'�1�0�B��[�q6�����4�0c7�&��=��ڳ�1c�At���
s=H��rG��e^OfI�s�(�f�1ٛ*?��ޠ �;t\eujʎHC�:���:F���z6�9!�S��������Z^��;�^?$���!�7�M�r�i�r���x!p�cg�vbϿ�G�^�n~mD#v�9�%՞c���o)�Q���g ۞������~�#������S�ul��Z9�!,b��Q�WSO|�[mUҟ����ٻ�%XG:�]�3R��{�ɝ�
�VC 4@�,��#�D�{�l$��5��MƙӲ^	Kb��1Q�	�8p�1�_��GE��"a�k�%VtU0q��:ȧ��AvW������S�<�)��'��C����ߝ��0�ے�уR�o-�b�!�_��SH3��
�IG�<��j��M��14@���&�'.,��%�xF5w���T!� 	+jBʪX���r���M]�Yj|P1J�	��-�6y=Cf���_�@y�~@�Ǔ��L�� ,��cgj˽��s�ǐ����ƘW^x6�d:�4Q�71k��Vչ�\��F�3����e;W�6Y`�cs��ʼ7���S��F�����
�^�\�o�Z�a���?*�h��@?��|���j�,$ʿ��j�5����B/���&(VmF��K���o�2/�Md)ܦ�U ���Һ���y�x+��ka�_��ۓ�jpˁ���9AC���ײe��S�'ǌ��U�Mۣ�S[z��v@�v5;��x�����J�o�)�Yz�{���<A�`�Wh	#�NЬ��Q"�f
�ms��1M�<F��[���.Ԉ��(�� /�ơiv�n^fSQ��Via6o5rj:���]T��O���`@L�N"�	�K�1i�эv���C��݊案X�� ��8�oXWa�r�6;}r(d�b�m5Q�K��H�W�����WՈ2�P\�P6��� Ԯ5�2�a����S��8 t!	E'�G�g�M��H�d�P���.O��-�G��MSH%2)��n|g=~=�į��B1�)3W���Z ;o)��c���Y%��|:�����iD�����.+7����:�#?��5��4�/�N�h���&g���ի8����g R�h2�	����༄E�w;�(��\;���vr�I)v:�\���iU�S�]�ډ�<0'54�,_�����S����^�,F������Qya�rA��ww]��4����Dܙ)��Q�JYHK��]2�r�c�E	�Z��
�E�N�w���+�������m2��V7j�I���¨��CY؛�?d�U�ZC#8��&��@�˕��+)��_C�R� P'*�c�-S^}sV
���zW)��n��o��3Y����GE|�E���7��[�C�TG梠+��Z�l;{�޾c?!Uij�ڜ��B呼ysї�U@|D�vp袐��/(M��.�	�> ���U�jg:F�65;/��Q]jI!g��hLz�8]J����9�d=�H �X�4�5���5t�S��j:Z�7.�����څ`+M�`
�'��Q�S�P^��'��*�$)}a��&�>�p̹;)�I�c����8�����X�S("Ѕ�9�$y�u?3s������`g�g�!�����P��b��0)�[�ƌ��p��r����vC╯��x�C=� �S:�dp��~9�.�y>U.�����֎o�k��n}����w?ic����11L����wA|9|�`�e�q��Emb4�@C����+����Q �v\�0ҡD�k�ǐ��p׼h]32t=x�r�K��Z}�Hr�>�*[�5��z�����bV�h�g��K���a?�c��k���	S��ѐ6��������9e�&]혽;�@,1�h}�^��%�yL���K���9mv�rĠ)����4����/-)�$*�x
 �Y氢�t�h$�����mCC`g�瞈���pwP���l�b�cbe]G�I�%�s��/�O/��*�ڄ�p}v��am���[����/b�c���*�p�]���Ě�)���#u�������Pp#�r3��PO#k�*p�(�7���O�-��\b�����-1�x��/�R06� ,�Ƿ�e�����T{�[S��~��#��Y��?�~��H� %���텴�+,�AM�cn
��X�^εC>|_�6�dO�֕�[��Ū�L{�������&`�^�՚�4��YO]��V�0q9>�X�.�4��{�)�x�d,F�{4M��W�c��������R�6E�P:#�u���@���}��W������1.´�.7\b�i���<�4J3~"�D�F���z�hS[�.*���}�-�7,D�~�@9^�(���\pœfr�������_%�B�Y(py�5GE_ȃ%�J̢�Ϋ��v��f�ԮX?_��sf���5"�ק��̒v�s��+B�Ǟ]7��F�V��V���Q\z<P�����C�{c��-'�
;�bkd:�~֘m7�	 ��<��Zq�!ɏ1��$�H�=R��_��"S��g�=��7�	L�4�1Y����&;ζ�_��Z3���P@�V���'X�J�rG�V��䍇�mO��kG��hR�S���{�vt>��ߣeXFsX����A�K"C����̬��W���d?`��'aH�k	���D19��tSb��ld��s��T} �s���u�d4*����Chd�]�U1��	en1�<j҈RLU��더���vA'a���q͸KS_��Kv��k�0��.�?d�pG/���STf�A!�DL_g��0��ҭb�)�u��)w����D3����~i�<��b�=���� _k7�{=����R�%�z���>�`�3�Z6D�Jp8���P��z����Ͳ\�q��.B1����Q�ج$��U���=��Zfӕ1$�o��`�6�����d�F���&��e�F��I��jy�W� ǥ|%�2�ȭr¯���,mZ�7Ӻ�:x�)w��_�e���u�ə���6!5�ˁ�0�sj_o`,�� ؿH��hV�K�1r)��J����r�A���QB�� ����D�ՇKuyJ�u�Vҭs�̧�p�� z�ͣ�UV���\�Y%�1��颯���/;3��,�T�%���K�bx�1�c�>+"]s�[�:hT0��fe#��֨yQq�g�Ut�*��E��^U�j�)G��7��T����N�mE���`��XI/�vڪpZ0�ڍ�Tk,g���ꪰ�b,���vi~��^U<�&���8�,�J�%�=j�K����K����ع}�DU>�7�%&i��2��r���?()'�FG������"Ն�LxҺG٬̋6h���">)8mW�1-���ƚ�s�#6`2O�R9`���
�3�tI��-��	���9�<ܜ�\.6~V�����1���{a�~R�I�ߒq�5*p�%HƲ��"�Fa"*�j� �������Q��k��yEA��ö_ 19�%�;���I�1䝢����|����D�0��T���[���w���b'.�*�������>jC�,v=�R����+���"F�c�4}Xj��ם����2rϪ�&��O#3%ZO����>S�cl���Z3N����E�lƹ�?ӹ����m��+?�Ţ�~ޣ�ǳ������W}h�ÍX۸��k�m��q�4�흀sH;��KĂ�����D��D�o��N�i|~���AEk5�*�d���TK܅vmA3"�,��+��BUy�MOW��9��l��h� BI���İ�C�~˗����dx�:�ᡥ�ԯ�]�r`��m�f-W��Y���J��#O(��C��Z�2jv��_�\��y����:���;�>!��m�c��xbLA����4)�N�J����c�aӽv�̠m�f���33\��-�k����}�1�\DP]\!�m;qXy�Y?`�8�!7^Z9�
4���g��Q�j.�Ru�b���)�{�	g���iq_LA{�6- XqI5�N��̴$�V<����Z�ތ���V��δ�zO����"z����B���Ĩ��NY��N�{+�Ef��!��_��!�Ώ�v����o���k�y�����mw��3'���x.`3c%-�D����/� kd}���~v�V); n��c9���+L/j.��s����ܳ_v�ӥ����6W91f!3BE��^���;���=�(*2�� ��e�"qT��x��Py7BfFG��џ�&BP����
�xz��ח.�4V,йs$	��ĺ��*�f!xH��'�%I�ny�0^5"�^��������9Q���?D"̴�.{7�y�����j�;@tXt-�4l�pQj�P@<�A�����랖�J����הO���'��3�'���!G��d��dh�}�ߑ��E�%L5GT�t���#�[Zf�c%��oȪ����a�+6~�$�D����L�ԅ��2�9�C�_㲭�-V9�KU1�pof��C[sX@̹@a����Ǟ�DgW�@Y��d��x���6�aԜ����Z�/d�o��浆����@��ٞ�a#��Zׁm��0D
\cv�$�l�L"��bн�=��Q�D�gV׶��n� K� �yZ�� ᴿ��j����1�/\╓}�cZ,ord,�HH3~u38O�r�� ����}�����| f�o�?�o18�lոa�p�<W+�ψ|w��1�;-ٔІ���y�q���y��ex�l�r��G��Ӎ�"��9�M�b�|�?�t9���c���Օ$U����.���༉����(�U��3J��f57.��RK�e[��f�>$c	)La�����;۴�=:+6�1g�s�Ra.1c%�RGI�z�[ޠ���[�� �W_�����-�21Sٹ��k����u��c2%J&$�נO��0�ӛ������N�y;Y�m]*��X�>t���
i� ��V�Q�IlT�%�f��PA�n�	���^?���Oü:_ׂ�?k��5��W���ς��m�4B�N]|Y�� �f���Qz�Kt�;s�Fs�sfa�F�/�MI��z`ŀ,���P�e�0jRh�P��>��I$���^�,I�D�TG]�RfB���x�]���g�𭶽Eh�����c�X�����PVvڞ=R�v���S�X�G�֚j�7h:l)�)��qe!7�M|h�
#]�q�|~��a�W�1~�Dx!l�?E�߆����u��SzxJH%זּ��zP��̄�j\����b|u��ܦ$���������Y=k��fnS�i���N���|��ޤx13����Շ�
�P7���\U�R݆M
�o�"�����9)'}��[#=�d;�0�N�[ى�t/���m����*���ln|I��ߘ�^�(?bҲ�t�c��0$���̶�P�E�L8�V�lX��)�$�J쏯Soׯ�Bx�ݽ 8����~@J�T�5�Gp���L仝��y�����aC�at��R�۰�q@��)�r��,_��G���������Y{� ��Oڔ=�wڮlL�v'�U��D$|T�&�=��՛�Q�����C��^��ta�Q���FO��f�+P�@��
B\G�%3���IXTܒaƼK�w�L��m289�U�yD�i2>Fފ�$��EG��� np�z�r��	o?�hI�'(���d�H�#����B��b���M���|Q�h�cgneW�3eA9<�s�#�o�>]|`t4�k�s���@Mt�W������[�U�b��Ƙ\���m�Xҋ��d��kO��;����j9I}?ȵOk�(qS��m��r�]!h����PFN��R1�.���=q���nC��$��"��"��G��(yN��6>Qn'ro*���H���Z<�	�>�~!��O5�<k(�b +Z��֚�'�`��O�h"��Ԍ�,	<,{�i��YN�.�
H�+:����g�_ã�o (+Q!��0-ge�l��g�>��7x+�A�OБ�Q���_(�-}�������)�;G���];���2��ry�޳k|��	�Lnw����ª�ء�J�{,R��eIX��N����D}s�Q��t��B�A+^����H�>����*^-�6jdtN4�ӣ)U�U$K%4�>�]�z ���l�U\�`����va�r&#�f���Z8�kr�8���]x�L����sU4�/D�~�	k�	��$����(h�FX���a���A�=�ߵ���Ed�[����N�N>�|2�:q��'��w��
�Ɋ\�F��a��H��̈́�%�����j�)n`�����̐��j���W�#����
P��ȼIk"P=S����]�ӌ��9��� ���P#�����#*����S�P�^#��j��ڛ�5��0�YH��D5T	��?{��*����mD	��VwXM/�9;V�Ī��z��21�����1��64f�����ԛ�H䓁e��}��R�E��
:v�8ƹ�Zm����4�Pkڶ�N�<�G�s�Eޜ��)�iM�X����d�Jz��#�I���UZ�[P�J[W(�����G�R���uF�U7�|_8�Wʅ���j��sV���\��2]�z�����|�I�\C��4<�>Y��h�tHY��@�����K|a��S;�z�Z��5�(2⨁���i)���?���n����`?}.+Y*;/�ACfC���C\��l�6� ��B5.�,�4�R�V���X�0����z�+iV�e+�AJ�*`%/C㚥}���p�ԯC ZReV�ˤ'�d(UO�9�����J��@e�t<���+��Z���n� _��/��h�����Q�g���5>R�BËI��%~������T�r��;��޴����,"y�(UT��=a �
ܑǝ@[��q�3���o�:�Ǆ	��$��%Pv� ��L��SdtN�T��V��>�-K%�� ^a�Ci�$������u�إ,JDm��O�G�S��f�Xp}��N�����Kt�[��&�A�'��XL��4���q�^�ӂ�V́S�O#�Ebƃe�"n�M�;ɟS�%�����f����$����N5ȨBquq����=����5&�s͗��!X���)�D��s1=ۧ�w�r��.�~��ו6�Ec�i�������epzJ�w
�C�{�T��<H�A�;�����(��?�mxP�ݣ���Lli\,�>S�ʉS=?i�U����?����WHY�e�n� l��V�1�p���V m��!+�o��^z�V��6Z_y�
�6(0K�tj2gş����yj-5)�~�
�UF?T�����:��|'�/����1�	p����F�@e[n�rL���w�T6b�Î�47m���>8�J�	�O�͞�=��~��ֿ~`H!}*�L(�:Z���$��Ə����{�Z:q���������<,�2w���Ɓ�k��90TĔo��8۞��h�]�'z��n�ͼ�˨��-RtT��D�f:S��X�:x�u�k�?͙1�9>��*n��͞YT4�� ���͹�qu��p>���<�\h��ti�t^�mT��[��-���! ��Çj����H�r�&?/��p�ݪ�&��B��C�bmG ��I9^�7\) �hW��U�D�C�Gb�͚��k�R8�(8��@��'�n��:��^�#�ص��[��5SX�IW�G����*_m�Td�S�Z9cV~�C�%]n���F}Zg=�f715�˦&\�45HXǖ�jg@l��S���p΋�	��ߗz�/���!�;n����l���p�7�͆�R��S:�TO�8��9��8g�!->1����Ï��V�ed�3���4��#!px��י�ᔟ�O*ɕB�a.�C�Os�V�`��@ŅD�y"2��	K
���\�Q� �dPI�$:b�՞L���`�Ӣ�4q��@5E���`������>yy�~L˓&?d@�F{�?в�5�M�r��#L���_��L�bh!-:�,I\�?V�����#��� @�*��Z�k�aRL�jZ|�9u��t>�Fp���G�� �'Pœ�ǽ���� S�9�
#��~(9��3�_��:6�i�"�Zfe�5�����?���Iu�T��}���tW��Ro-]�Q2���Wk�j��4�=(J%r�����p�U\e�)EH�����M�lkK��R��в�c�6��³���j`O�^$�~��E#ڀ"�����'#W�N���RKzܕU�pk���nL���������"�&�j���
�ZD�Y���21��x������Ra�&k��a��'�V�6\�l:��/�p_�K.���y�{_�ok7��b3P�O�e��~}�'Ʋ
1����� #94][�p��y���A�b�)�վw������,]��p`|(��1�<�� 獆D.�5������ӡ����I{EM݁���?���R�rV���g�;��	Q(��bw|�I��Hu8�s�H[����V�� m���h�F&�< ���=�s;��;��~\��TK��� �F: �s�)�����%�!�vK)P�1�(;���>c�����C)��#��4��	���9�\�#>d��Ev������5�s���5'�jJ��@i4���?�f�4����a����v6��Ę��(�\4W��IK�Û���;-�)�q�^fлQ���`ݯ�&I�j���ɰ�<tញc��i�cGZ��ʆ&LH�룛Il�q}��n�����`Dz�5�̹Y��΁����M�B$y`����f"�V,h a��v��d�U2SzB@���RM΢K��EJG�z�>�G:�S�˗q����C���aYMN�>G�쳼+G����w0=���ß�7i���4zE��)�%�����I-�����Z�%�m�<.���+u0h����l;@�F�g��.D�L�^�fB�ݫ���,�I�6I��7���ȓ�*�]�d�i�7[�z}�[���m�_�:Qc��c�z)4��KDco�G3Nu8G9��&�JY�#śY�H�P�����Q`2�d��$D{=mn�ϱ��Ig:��_�J�$Q�aV ��6<�`x���1�S��!���#j�+̫�N��"J�������~�H�_S"�MOd1M���������8=0�#~�D���u���| ��όO���1�YX{w�1�ʆȮ*����YC���<���S�0>7�����r;Vtt��kw5�6ޠ���D�"��!�Mc���\<"�24q�u�FI��������WD�O�&�4�����B�rT�=<"?��)�K@�>��>�RW�ݡ�{�,n�{��!~�	*i<�ʶNK���Nh�{��t�7�S<}����OM	�����s*^Xo���E����H�xuNY�6�#V�⴪p!�4r^D8:�n��˻qZ�b�lM���D�Z���5������X�0��UN��`q� �s�g~�ܠ�������%�'��C���r?����UM\	N��b{}U��dM���.���^ɵp�hJ�Nв����Z,��cQ<�����[v(]��#���[1�4[{n�Z�ҧj[�nׄ���;D�E������ ��0�A�m���n�:�-Bm`�U��To:T��������KC��r� �H�r3����[�cĥ�k�w����e�#�-7�`R�Wa���B��k���jԝ����p�{���0Z�(Z5_��F%ZXN��v,� ��ks�J1Yڳ.�۷�?E_�˖�̨��8��*HƉ�D=D;�M���0K\�	)�-�a����:3���+�p#���⧖��v�.��5H�O��	���!g>���ʡ%�@9Q�Y��¸����zq�����:P�G)(���q�'�>�_���FY��3_4�i̾��P��EW^%oҸn�����b��.e���9���4Nߎ�U��f<�<���ʨ�+��dǉ����rV���8>����Mm�?�B�改���gQ7L�v,0��rñ���j��il��;w%Kp�3Uԇ$ M��-������
�
��Q0K�ↅ�9ݕ�L�k� #��-�����NA��5��L-qn R��;�MSE�&�k�xn�W ̦����,���)쩝���Y�?ZՈK1�<@H����;�-j�!�fG�2-,?��!19������m3f�*XTm@�Y^qf^�࿭��5
����0Bo^*�pF����/i������u������8.G�τs��Z��?~��z���T�"'�TPt\>����9w�M�@'*��!�=Nݣk�șN�'�۬eU��
�@}3}-g�E��N#�@m��H T��]5�f� ��^U��zQ��L�]��s�iY���9�.L!4{)fK}4�Kw
^�h
���[��Sb��]^����ݟzҼz�`��);L�a��W�S��ʿ�a�-G�ilm�O�GNP�o�كH�s�^Pk%ò�b��	�s�l7qLBX�j�q@V�B.����\kr�#�>eȒu��#lQGM�k�- <j���4)�_�;o�PK�4���A���8���CY���Q��X�e84�l˓�wP�tʌݾ��-_)U*/��s�8��:�Y��- ���o�>�..'����B�ķ�0N1�$�z�H��kx�����;Ⱦ�����v9���Gt���x�m���q��.g+��gJ0kw���R�9
{fG�^�P�̽X�; �x���.8_��Gu�<�����2��0��4�8�bV>�>,�ɤ,��^$W�31��z����Ap�Զ�؉��'�ߏ���m��)0GK0,�k� vz�0�3�jD���Y�q4.Kk�Cgyֽb������� F�)�J���R��`�s�FЬ�z3�>��-~��Z\{���ztO����s��{����8q�QXݺA�ٮ�y<ߚFF��;�n�3��x���|y����Չ�aB�!��o^�:.�̘�R���eb�p�Z?�� Y%r���+�����K_��ĮM�#� ���UZٺ�LP#z�$��%��vV�&ra�B���I�	��<�|/Ԧ�R����9�Ô���no2hLӓ;tb��	��$��-/tFNg�mU�XsN��8)��n�8��IՁD8�� eg"~�ӑ��h���j�l���M�����m{_>��8�w�	�ͭ�z��,s
{�\4�mtS�_����:x�g?w1���x�� [ aC����B�[�ҧ�V��� �W��\���8�U�>�5%E,�Ց�%��-�|ZpnNXrn�8��'�0E�C'GIXS�I$L�^m~02�f��=�1�KI_1��)JF9K����{i�9��y�֣��}�B\2W%���D֋]��z1ט�����"�aU���dOb˨6��J��nV�1�/�uz���@r��0��m� 6;���i�	a�2>�%�SO�Q+}R��~	��4P�������eJ3.ݱ�����{�6
���Mr�Ę�龫r2ٵ�Q`�j�S�Ȋ5fi ��v������~b>6k~9�����\�/ ��IDd��k�7�-����g�/���-�o4BE�~i�o}���^`�מ��h�|����$�~JA`Y+�=2�>$��8�F W+yI�?ؚ��c�h�~�"���t�cM)gS�|k��̎I�M�"�͡8��"��u��x�h5�@�Π���仚�O�p�����@N$�NO��J~��@*�]���(���C���@�,Nz[�j��9J�{��ӿ��̧b\��F���ӷ��M�>J���@���,aTj�+�ю�E	�_��7�߻h�����?􉲮Q��$����J��H��r�:�u ���z�՟�)E���r1rz����QgGi�� �+a�8?�p7ú�a�A]o�mE�~=��������t�;2�r��٢:��%�Qo*a>$�2�Zz)o�X��ȁZ�c�!�j��u����H6�d�q )� ��Z�x��KK`�ܸ[y�j,0˓K��fb��TcI)����鯞�}?>�������k+F�NŬ��T���� �Xy��f�,IS<���oys��i��v�4�Jgۆ.f�.m�c`ـ�m���M:~K������댒��O�-��m蕾�	E�������ڇ#��J ��j�SiR�O�,���U�����f�=������L_oU��{ I�hp0�_�2D��˅G$<p���i�l��� z�*$��gv�-��]<�uD�.�n	T�w�9Rm�`d��S��}�)��؏�~�����h�F�~�����%!-�M��^3��2��At������0�����������Qx��!�!�ǣ���i4�))#�.��T���/�p��Z;Db,֮�5���<c��s� �w4&��aB\��8�2�QTl)[�f�8&�e֖�]S%\Ǫ0H���G�myT�Y�n�؃�?O���a��J%S���W^�K5������V�m8��mҁ��L�0�NA\d|���Q>M�!��u6�7^�
�Xjgӡz����G�R~b���7d�LG�� ~Ѥ�\N�'�EP����fo��0�\NSӑy�y�ј�b�� ���'�U�<�kD.�5������?�0�F���L�Ƶ����G�2ϻ��e��a����ݚD ���j��f�#��u�WB�ĵՙr���^˦��8jB3�	��l�l'�/;x�p��;qu�5'J��L,"
b>n�<!ZCp�8�A��[�G*T�r|9º�����~��Ic2�3�n��Xd�vtf�~y����<��_֕94K �Ԣ�����s�a� ��L��Y;D�9��r��YHW��n�"s"ۥ��A�	P��zx�k��>@cC�T��q�hJiwp��#}��92Fya?�8�	`�5��Ϯ��-O3q�'0��ꎯR���3R�q�V��	�h\�#�T�B9���W�/M3��&0�!�~�/�`b�"Ne�d�����djD�R\����3������FC������E!�yp�I����V2"�����gq:G�&Z���i �s�y�|Wu��ed�V��']�0������~נ3C	�k {��^&���ڏ]���N3�$<\ ���@*��������-+���kc��R��^�h1ڹ���`�1�V���AW�9}��V����������Q�b$��&h&- ��B�*?�����3��-�-;6��X���H���n���M�g�ڑo������O�ı	� �!������L���o�����O���5��`B��Tc^o�V����\��J�����N0���7d蛜e�DQ�~�A6.s�K��Y	�;�5�X��9��w���d����9BRz��3�� tZj�&R�g&�o��ʲE����m�p�a�RCm�C�a�͠��E�����ժ�ӄ��	�K

�,��T�O>���/������&��܁�*k�=YLF�S�;]�z��tI�xһ	��t�x�tq�����j�C#�`�[�f��d���c̷+^!�v��5@v+���>sHN�8K-��n�p�.ՕuYx�!����<�b�@@�%!�h�)��8�pm�8#���S1�"^N[�ͻ)���gJ8���'Z��0rMǔH�YJ�|V��p8�)��qT)g����ۡ�����M�� �:e���ų����?,N��d
\��G�A�P:7"�i�/���Vw�!<�2В�u��?���@��Om�|H���(��Vُ=�v�e�I��BcU�(2�й2�;�����	"m�c5A-�R��*���JA����Ÿt��I��#�jh���"	q���@5�`�+Ɣlhu�~<q�� �iа ]��1�?��Hx�����r��Z�O��H�$��d���&@�����a{nneB²��+��*���H�/��z-[��3�=�#FO2�B��
��~�8t#�b"m]�iג����e�.e������A�lŭ ��;w�YKĺ�?#�9(��0���hi��QFg��&�g��iގ��aZ�����c�J��������i�S�y�0��a�����G���m�6['.͖�y�&�#��֏��Pą���j��*��䶺���Ġ�$�ĕ%m���[D���݈�0�ګ8���h��C� ��q��\�7�'L����|���\���R#i$F��v��mw.��o�#^��~[
��6�������/衿T��a0-�$D���5�bN�S;���pm:f1�J���u��t3Oj��*M���2O����>�"g��~�C��q�%l�d�D�j��'�UH�BSD�R[)�9I���ѳ���5��E-��i���.���ch)��:��Ȑ����qW�h���,�ULֿ5o�o�Ğ*�������F�Uj�}0�Vm�|E i�CS��8;��R,��o���Q ��q��pQ��5�`x o'�8�m��_%���D����M޽3�<�:<<�=J��jŏabp�CE˓�&=�]�o���tt����L&q�C4R�w��w���	a�_�^&�Ҝ]�~�_;ϐ�%�u�ρ����48�e�\�d��v��A-8M�_
�	�Ҷ��7M��ͩ���n�����S��=A�ՒD(}�r���+0i8��qԂ��*NL�4v)�wQki�I���b�,gѴ8�ZЀ�BZ��k:�7K��	K�1���Th��.�OL}�5�Yb��D�������ج5�J�B�V�h�;�8V�����p֮2U-� ��ſ0����r�NX*����A��/ϓP&�d~� G�b���r�h��ȩ\��a���?Z�s(�����C�X��<����=�AU����\��}O���o�ru{�D�.8(}P����3���) �l�3���$�a��cb#���p὇�C�t|�3tn+�b$C�}% %˄�mM��!�z�Z=A���Ic��K�Q,֏�#TӰ�v�9���pm�r�cp������s���Z�b�O���<a�(�z���$���,i9Y���KΓ�����ec�D��|�J��K8�I�?	��4�,���1�p~���n�┽��Ģ���4e�`�c���B��'�̬���L���6Z��dj�X�A��]fE��D>ЌJ�[}JL.O�@tSy_ �,m{��Qc���G��˥��b5����K��R��m���Ȁ����t��i�:���d��C�H��:�.���S�C�5����	����@�����S�LV���S�L]�^��}��`�&t��:��<ȑ7M6Q&a*Dx�?j.����U4�i=�һ��Ĕb;�y�CHL�[���_fT"���|C��C#*��!9梱���D� ��6�Sh���3I�n�C�&�j� ��D,���LhM����Z@�x_i�8Ed7���d�I���n�	��0�`Ԁ��&����f����Xs^���y���YTE.՘Fz��ɜA���^|�T|N-��v�I������
*B�RvVM�7k�.Ed�������-���=�����<I8GЀ�6L q礅Qs��Aԗ4������~w��8�9�����I�9m���V����ز2@s,�;��B뾣��2���1���{e$��e��[u�q}�_l�%�C�ʉ-��U��Sm�^[��X�i"�`���;0Lᇁ\��D���d�����{�H�ۤ���Uq�B���ؙ��\|*G�N��D#ż���06ɟ5��֜(���J�cH�#P���)5�dK�9�����Q��K��%4��䱿�IK�Eҷ'�*`>7�q��u�� �@�U�ѯ��IvFY�ï�K5�J��ι�j��|S�J�씘awŞئ,��N�t�ż_��@���KG~�P�u�E���bϴ���x!CRi�i���K~�c���X���a��pID��_n�-�Ky�T`���?n���	��I����cp�<%:%�'��Ր�i�%�o��Q�����]��s���'��x����-����`YAb���u�I%�A��h�\h�fuN���>31B UE����%��Ϧ�gM��9l�@�\M��I?��VJG��^̿���}��jX�׫{��\(f/�A^E�p��������x���n�E?BXS��z7��vUېڰ��8{��M��=�ow����5y���ӨD��^��b��$mt�#�aY���&���Æ�	R% C�x����t�f"~h�V����L=�!x��f2P���b�X� ��\;���H���c,_.��˝<�@�N7��"�N����_]EJ�qe���0��gvuB@�r�p����ˁʼ?o�\���)���g�1
zg�E��h�E���������]-��	��:iϝ�w�������A���G��j�Z\��r�C�u&N�|�^
��.l�͛J�jI������u5ef��0,'˯�޽n���LXZ�pև��E�*c�S�)C�,����Aޢ#k�/R��#	8��r~�N"U��>v=;~�m�H�kC��֢<����v>_���
g���ʐ���&�-$�wh�,��d.[�#]�r�9z���9I/�C�(�SƜa�5�8��d���6!@��<�o�Q��e��m��]�΁��$���Co{J�l��%���S�ia�0.!o�6-�g�|-Lp�Od��f����;���Q��S_յ&6�H�h�-]��FD��ʘ��G�b�[Jܯ�'@C�4���2Jc_�.���5.�vv��KM\}����n�'���CkAm��C�^�������8�r�e��l����|���X��ثਂ^�z�fP��;ȇ���dfzV�Q�������BT�Z)��c\�� �J�z/��!�_��\��rc�$�0�%H��pH{��uN��-��<��+������H����e�N���Y�
 -Ѭ�NkSH�w���9�����C�.0/��h�̋I/��:�i���� ���{����75*8@R��mz�($Sr!p>ҳؗ�v 4��J��0Wա��}�Į߸�a{$����X�ʁ�����s�=A��˭���X��ØR0U�)��r��G�c�c���(�������\c'�^#B����)�S���6�M��'?��;v�i�yN��5�h�1��ksb�z��`���7U�����w]\L�H��6�Z�`x�+G|9qRX=O��_L&�eʦq�_��_��Y@��lQQ7۪�	+i;ԿIC"�#Ã���x^���7Y�^����q�k]pF�Fߥ�ĳ%��Cʦ	�,�v�Hł�����O��-� Lo��&qX�����]����}[*�N5������������"����YPd���M%�bg��-E\��_�Ă�b�8	��^��`�B])6�Y�>0^�+3]a�l�	���ѿ��h���<���@2��YG6�Q�)z#��RTQ��v����{�uq�`�����RTm��'K>8>���?�����������v����S;����Ѡ_l[O]^�aႨ�Xٞ
)�,+�)���mE��P�7>N��;�gߝ�z�$��ϫFܛ��E��p|ܹd8�5����i���"�z
.NRp��2ͺ4m�J�{g�)�~����]�h���'���s��n!N�n�zL�T� �r_��I-���1�T����sP�����������P�����v�3���+30�l~R���Y��q��ۺ���)����b�1퉳?NϘ
z�:���_C3rP�!�>|e���dZ�D���i�V�g�}8�<H�KL2 ����s���}ɧ�de� u������3� �\�b�T�5�-4�tz���s�+Q��r^�;��V;���|���)��"ג#mڤ/C�˘�Rr�ݶhe�!P/s���r��V�F�w}���S�Q�Q�"	�]�/�5�K�aƮ�x��	H'B�7�I]M���ýg��V��O�׷�|��m9_΅�h�� �t�_��#}�v|s�B~B)���+l��p9��h�r5�:��-�V��R:	y�P�ŮI�Yg��v���Ʋ����I���4��/��.���;^'D �#�5?�\�`˗����Ih�䉩0q_�9�^H�q������)��7. �8��^�l�~�g�t"`zH�}�|��Y &{���$��M�����2j��6���֠��]h�b W���9�O�#��I�����&�1N�H���D�_*e# )#���Q�\4��o����Y{��Mw�B0K��V��QV2�2P�J�������<i�Hzl����'1�:�@� ��"��\�V�uEbn��n�"Jb`�?���x�ǁo6�o��$�p���^G�ڎ��&�Cxȱvj�
��H��vkҾ� V�ႈ�Wu���Zխ4���{�V��Z�Q_%�I���-����@F�p�vTTП}�X�S���1.�~��]43(�LR�W�|X�+�NRc���	����J��� ��[T-�x^Ң�?�>0g��n\sM���a�x3� H�K�����u�� ���U6�P,�ם*^$�e�p���
���P�-�?D�j���e���F�����V���i��\��w�엜� `�y�����Mm��V���.���A�I�����+4B{����!x-�_}'"�Q�%�&�z��X�ç�3�G�j�D�Ć�~�gkq�|�Q]P�#4P/M�' ���<&�r�m��2:�n7'��}j�k�}���b 0���7��ڦ˥�l�Ġ,_�ʸ0�����]+:�:p�\�l[��&:P��a����SU �=^Vl��}��Z�oFd-���D��Z�N��iB0/��`���=�����/�wf��|!����1#�fL}B�5�4��昻����3���[I_���c��Y��u ��U�5e�'� �k�����z���r����D�r/�x]�@��F���{������]��;ez��9t�>=��4�%뻻�e	�t�e8R3�* �1]�� DF��*�_�hn2��,x�}D�]Sw�I����
��P��Ez��0��ACq�>_i�=䯚��ڜ׳)!̄!���������U��Bk �/��y�׳J��w[��N�cJ�r�V{��Uo��r�*��{.Bf ^pM��ޤ�OI���X,5��ǫ�R�|I`�rm�B��n��U�>~���qA����6gb��W���dA�y���j�m�o�V�!D�/�W������N�2�K$F��^S�/�l��;��P�N��s��k]��]%�c�H�
{����:�����r4�v��ȓ�x���fi��m}�u9fh��N��׃�e�^h�lP@0����/ɽc$��+�+���� �h���Z���M��9x�?�!7&��!��?�o�l�ӷ�"9��SH`�]����#��Y�]~)��n0x��al�_xT+S�P������c�3>
���Y#���s�^�T�:ADs����
U��Rh�.y����2�P��Rxu1Oo�B��hg�-B�,��7l�7r _�B/�\��e�>9�D=��G,�y�~������{�{f���o�n�s  5b��G\]����|əRI�j�5��,�c��W���")�gG���Q���Xڕ�˨�CJ�z�֧�!��`Uw�_�W�\��o����s�Y<
Bm�q�{�Umm���=�>v�{=��U���	�x�qYF2c�6���~p�h�k��[w�q"�ǽ�����z��s���y<�yk0��]|B&v+#�f���/�w8!_Q�ğ�߼��}篏Jz���i����n ����I���<�%�����ÿ�8�~~;8�yB�Kl$��i��Ș��OJ�l��n��ȑ��3gt�쁒45�
�\�����aO�>e'>qӹa�b�Z��=JO��6_�f���
o�c��kI ��&^�)��� �{@�yԜC���)Xjd|pS�F�	 ��@g�yZ]�6�L ��5��1"�}<^����K,P������7�H����Us$$՘�&i@Q�y���$#BU��\I�셕;�վ�O�f���;�e����
��nY��ZR�[m�u㡆�\��b�%:���y����$m����A��n��Z�l�*� Kttψ��;(�}���/к����8F�3/U��ڢ����LG���|�YmESּ����\@: �-�Y!��7���Mi\���W��64��	�4���\���{Oz���G�Y�ʫ���	M;��x���e�A�e˄�5:j�4�!��ڭIc���A ��8�U-�p�. ����4����މ1�*^������p�C�,��_�����RU�T��e@|���g��(��EM�p%�	㕈�A�����"Q�Gcj�=}#�ֵ�>^����<MpYݐ%K��پQ`�����\�=�{L\�mBr�^��S�A:S�5`I�k��p+��y8�w�Y{�_HȆ�S�񔤥��ƹ~�l�!k#i�>o�N������������t�W���� ���B���n�>�enAMM`2����I�� g��a +0�*�t��C���5�,�5������?��(/Z�1��E=7�(,Յ��k?f��o�)���o�8]M-��R���#H���J'����s��!{�������^f�%;�������*q�+p�n��g�z���ìA����J���T�b�?��$v��E�κY���1#P?�;X1�3~2�Z��bQ��7�ˢg�1�L��(��V�˦Z�_c�M�MG�|�A�.��`�sV��٘�_l�/eg���@�i������8�v���l�zK2��e��[�שּׂ���R���[4���W�06K�i#�,�9���|��,;��"V:hx�e��P�K �+�d������jEw����X6�?����o�!sj�����Xob�j��O�^j����\s�}Υ�y:N�C����J���E��eFO��$��.mQ�ϖ�)�4J�lfj�O�&j	�vB��ZA�}�	�ҩ[�]jz�oߊr��[x�C>�Nl˷��0Z�����k���~uݛU}m��'Ŗ�E?O<�X�x��v�2����=a>P�6c	�!c7>�!�De�b�h�Ea�߂�Ѹ�#A��2����������⢼�ػ�۪��c��
��4ׯ4���y!��nM��l�������ϙ_�1L�J�Y%�@����1Qv�'T�Mf��R]��zt��n�B7&\l�:`��ޏ(�e����v��5����U�������wu�?bq$~uYv��8������@���*��"О��, �ruԵ�*a�ÄZ��Mp<�\�9�a�T���r�=`{p�)�A�wx���0�Fm���OL�LJ���^��l|`��}Ekp�L��J�`Ó�U!ۇ�3�r�a۶��9��ڤ�]�x��vZB��n�i(�Z���.v�<��K�*���u��W7p��1U�ؤ4�m��2�9�W���zii|�ee�I&
'��w�����^J�$�}[݄�N�X��E)r��H��v��>\��T1S�(1�;$�/���:� �A�Ԕ-��cT����x80�J�/ l3�Q�{�����B��m�D��0S��n�kb�l�p�����s�ƞ1}|� (5�mv{�4�2B������
�+聅.O��"�v�*�2�q	!2��!<�K��`n��4�X?����:�z��S�@�H;"�$:�0��z���bw��ٙ�r�S������%e�����G���_ aVK<>��4-L4Ѱ��|i���i��UBh'���V�`t���f @��P��]�3�g�V��tߎ��R��.�k�V)�?&@���h�@q:͗�!-C�s���:�S�L�8�1Y>��,Q�vtvc�l,/l�����TY�w��i;��M�E_Tm�?�_:|W�=�9�v���8� ���,E����}�M2��pi/B��<"ϢˎUЙ{�>��� toE�o|���6c���p;A�5>��9hv���u`d��[Y�@`���ռ`ł�� �g&�ע�	�(UC6p��EhiV�q�2*ݖ�+�s.�0�j'���%����뀇�$|���ʝ�xe�ݕ��m��=��Hײ���v��ڴH�H>$�dHJ�A�{�dX1xO�A��/c���DY��x�J����q��PQ(�\]|p��#����ϙQ\�Fu����!+p�Px0[�����X��ATh�z;k��a��Ί�(����Tj3�~ 	����~�A���FFY�9�	t�:Hw�"(޴�X8o{.6��<A�遊O̦._��lc[��3�&Q=�2`��~��*֦�h�ᨴ,�::c��ǀ��R�O�d�@�p���܉�{&���Yz�����[��sp7Ĕ��K�~
vq��2�G�%I6{��F�6��ҁ>yF<$������V�Y��+�N�vÞ��B��m:7n 5!V���g"��2ݧ���mSJ��<f�A��L:h �����b�F7��Ϛa�˒�-5˱-��h��a.��Nß<T6ʡ�)���볾_c��6A�o�y����1q|�m4�2��KJkq��4N�H?@f��Hy�N�zQ���#��B��Ez�E.b=�U4�M"�k���p(�}(B���N����YؒPk���5��΁����MԔK,ٱw��}W�aH�I���Dc'�ak����������~���xZf��@f��zR�{�k�f� K ��Ǧ�LQ�n�_U?%2�TW�6+��L>78.�z8fe(�@D�Z��E�|�.��i��,�#��px�� j >!��� ,�D)x�.���/`b�$hZx�EoC�W^K<]�Kj�:�Ю#��gSG��Bʃ:����λ1q�)���V��|@|������&������_�R�xH��2)��M,DJ�
��jG�ᡰ8�%�bJ��Ch���cԥ���"ֿ��RG�|H��VP{�����Ӈq��p�֕�.@�ډ�o�X�n,���#���8D�29��O�^��`�D���?w���f�QZ*pU�h�@�:�CU�&��9ӷX�h�$z��]���W����3l�2�Ѓ������.��S�/�B�[��r\�kx�z��ϡs����S�u���<����`���$��Ea��6x�H�r~[�g6Hc��k��bˆG�B�M,:;fI$�8>��w*�c %��@��M^�um���j<��s�gLk3��k@z�O�2R��(�Px�;��̉�bqj�&�\�Յ���u�i�,Z!J�L���V��N���7ϼ�m�f��XL����������/�G��� ���l%c�#�S=���I�I�4�n��%�X��8�4�u�hYG@��0��24���@�t�F���ܤ��i%st�,�\�=O/H��?R��5%杒�,�'���������o4�z?Ć��lYN+�(PV�2����.���}�1���ћ����1����-掃��A��Yʆ@���֎�Uw�
�n'�<HQ�ǻ�ת�X��zn����I����I��k\� =]wm�%��P$6�$t>5�5�*����Hl"���ì�����j�6&T�X�I�� z��@����ºF�Tlrz	�Sdzz���Q��?�Z���9����Q�9H!���#I�\���9��\���Z B-� ���Z9��_{�U[w9�pD�Yhg�g��O=^Dbh]�Y�nv�Z��>\ֿ�#�:�6��S���RZ���-�|cH�[�P��Ólc�	M�'�mt4�Ibg1%�W
�Y���O�71�c0u)��oY3�U�\�vk�������X���R�
�xƖ���v����,%�ɷ��.»�����W���88}�?b1eB�n�����p����ىi3�s��՝�s���|�f���.+��x�� ��2D;�ł�:mp�4�ځ4R�o���[l!�$ɩ9wm��ڤ��2<ʡ�R��
�7k)�z�D�f�e��6��@���h�d�������;9Z��S�9sԐ�3>,6�',(\���{��AaDnD��*��ԁ��v\2"ޭ�P4�0����K`�H�-�PE֣��uqY�4*������]��z��v|am�Ǟp$#�?��� sB���WQ����'���P	��u��Aw��^�Jj���Jۦv���˧8 �R24�w靭n��I832��;�&r�[�2�a3d�6c��j_=j��C^/�вq2�H���V��^VSZ̺���vT<�߇�NOe���i�!:��R5��S�i���Ǹ�`�^�t��ӵr�����S�<ڽ;�g���Y�@ns�z���s/���}nF����W�v�);���-��֞eG.h�`bb����L�L� ��L�z�I�JƠ��l�uaA(��~s}D�g4�P t��eZ0��Q>=�$����j3\/Yqhz5��Ax<?P6�5�����O	�,JGW�ɔ7� &��lG8�<�"Z*Is�#�ym�g�FT��̵q �;\H��G*����Q𛦻��s9-�ˎS����o9��t�U��!�-��Ki�2�zNgӿ7����c�y7�g4N��Y.�F����D!شĥM�Sl[f�U��7.���b3��cf#��<R��q��q�3A�}�}Miǌ��\��I�?]z67ڬ�X�g���J1��)k����oą�p�z.��r�!(-�U� $�p;�#ĥV�!S��)����� O0ȩ}$s|? �`��as��Zn�O�M֩_����w�i���%a���}���
�%-S
���M+����/�H����=��yRo[`Y�l��)o8�>�X��t&��`B�{�6<п39�ރ����y�C�G��)ӵ�ޚ��J�g,�����Έ/�Y��,�t��J�V����v!Y����%]��?�{��vR�jy��ѶWRs	���n��������]OH�U�{�Q?\����ӽK��?X��,��L/g߰�����i�)FM�����VD3Ntb!�a/�=�ہ@r����ݏ�>��C��w��b$XI�w���\0p8=�/yK_�>G.Q�i���f�;�ߖz扎k׽e���Ԅ%��_�_�����z�Ҵ��.T����p2Y�Tr�f���dhm~����&��otFmtHy�\�tX�a;��	���/ ���dj����ed)��v0��,�mcK���;�TE�2>�%ۼ5��sO�/+g�suY�L�z7�t�7\�%5hk�����P@7�[�gC7���d(/D���<
���C �Y���C������tX_�bc%٘	���>�k��K���WJ`�T��.��py��C�����j%o�.�冧�U(�$�u/�3BHz��7��)"�p ^�t'p��<Y��}a>��k��{����qe��_���zϡ��Σe?So&"*�az ��*��ݮ�:i���,q�%8��嫈��vK��\Ӓ��sa[��v�u<�",�u?�m,��B6�D�������Hf��?��f�����l���=We
���:��MabC�2�j�5&C��R������Rդ>Z{��Nb������[5ʙ���4�szSS.s��Z�F��od߁4�;���.�Y�eq}KZ�H*�qF��� �׏n�p��Յ/�I{�@/�(��LS�7)�"�9.%��I�)�`?�1��R�u��}�|����h��,O	ݓ]R�G��@�rhc�O�Y�Qn�Э�uy�6���F�6[1���29�{o$6 ��@=�)�_t7��!�]5��ez�l�q��-	�1�AkD��7�8��v��I�Lز©ڙ��W~���G�fv7�U�FF$j)��	Įʕȋ�������g�f����G(���t�k��~�ۃ�u6%.!+&nu�2_�j���eߺ���[����#��R`?�ε�7_ ��F��cR9ܶ+~V�9=�n�eF�$��ơ�Kd-�H�$I����h�oɬ����`��asլGI�U�*P�#1YǏ����;P����(3��|U�����J'�R���.-�%�����xJ�SA/mSh��z^z���cD��q�G�^�+R�ͮ� S�L���7Gn��^
Vk�lL#�4�z[d5a���`b������c��È�Qd]��!<!�-�o�>�fF��)�}�^�h����~1�洲�v�0�S����8ͬ6`ro�<9�R#��M����,S2D���ٮV��q���X�<N�t�$��q��I�����=���!�	�د��0���o]<�(��k�D������;,±TP�IӐ��z�fb#�I���	B\5���m�ش�S/���ͧ�9=C����r���fT�Aj������<�L�N���|���u|)3��5��[Y�h��-A�^F��U�����8΋���u ��o��=:v��iߴ8�MJβ�O��I�NY��^oe;���{�Y\9�v���b��n��G9����ϵ��af>p�aH�̇�
�?1���&[�Fa�:�EI��d2�s�����M=���Cg���t��1Ο)��4�Q����N��Q�:�>Ϋ6����d���A�۳���s/WF�+�'�����ą���Wp������,���{�&�KkH���BM�<	�\��
�"E�ť�y���oS�4#�$K�@��ӑ�r]o���>|�4��4��@9�s�U��2�؂yi�KC��2�U[�����Uцc[T�m�q��wL;�U���2��A:1vŉ6K���o�iH�Pi�B�!+��ˠ@75��_��u�f�M�e�A��A[^����.�g��-����vq�}^�c<��|�/T lX�ٱ9s�o�)6���e���ex�A#�o�Q�#�s��~�?K|�/t�����,�T|���eݫu�N6��?�wq�|b!Zӡa8D$��MB���@od/���9�օ�9��P^�Xҷ�4,Ȳ�o��P>n'L�bRC6�O�8ڦ| N�/�pB�Z팷��ԏ	g�����;:��[�㱡V?��SL���*��`�* ҢZQ<��v�N���0�^� b������B����0]w(���ԆwC�Bm ���ȻJ��D�W�/��csl`�)��]�L�Ӄ�}/a��4�!L���>�ުҺ�l"�M�]�_�CE�J���Y,�j*��P�#于;���>G&l���I�Q���fgǂR�����m�c?Gt\W!F���j8�hY�h�\�YϞ����������O}c�K%�{9,UE�+�AC�p��3n]�F�T},�*�lj��Z A�F�.S4��Zr\��~2�Ϲ��3�C���:���a�5e�����i0�X��eXR׼V�����`���zr�?̺��<�����(UMh,e1����/�N�L���őa��n�Ͽ���.��(�h ���n���]��0=w(�(,4�N��=�6�3�<N�M\��o�i�ب��� ��'1I}Nƥ�&�G�7���/
/
�b�c�$qˤo���PI�Hl�X�[z�ִ�3�e֛��l���Q^��E����)qh�2S������([\����P�|0S���<E�Jٲ�C�-�L#��bi�9��n��/V����5�QCl��5��*A�}1�3�:�C�������/z/��^���}��$��&����a~C$��{��˅�~�s{�D���3�&;XO{f��.V��+�5ך>ƋR�h�}�y�v��v�&>�#��=�a��P�z����[�:������jG��Og�]�|kr�K�ж��>���qV�����KH�d�q���R�>�ۄ��X�c�����<[���UX�/�(Ggǿ�\	l�@�*�b�Rm��{W�p]R|(6ׄ���ֹ*�DH@cw���f�A󧁰
���	�k��EL�Z}�prtR����u������)���y:�����Q?_�{��'?X�Zͤ�Ym5a��(����"���Qعa,[�+������3%�jA5|�N��r���f�a���;���`�
��8y�fSR�$?���g:��5N�T���1�����Y���ѯXx��H�gw6���;y��k�x��_�>c�C?S/�h��Su��ӞQ¹ѧ��� ��+iy���k���w������@����'7�6�jQ8ipp�R�X��\��[�@�	^n�����D�C~G����P��ւ4��n��x�.�@lm�~����J+j�N�lF�,�ȏ;1iU��	Uo/�q�����F�S������J�rKQ�I��]+�%����I-���K���l����bʪ���{�9y�:s=M��~���*ӵ�����'s`���(jH����m���;d�)T�hQ��M3*'���gy����Bl��/�\#��K�n1\x�ᒿ�[n�h��7��#��Y+�ӯgg Wg�S��6�xd�JU��W��D՝$��`��SӐ�@�=g�v�R�b?����(}BĸL�g�Ne7>I������jW�P�yqt��y���;�(j M9n�C!X9�f�)'��&'y/�m��tZ�C���4�bn�6���N��ΊT��t�V�����Mb��
�J�?�}c��
z��ag?�AgU��ZBL�x59��[pdY����9���G��"B�
��_d���Fb�p"�ɚ(������a���u�.���z�'ST�/8�l,�/��&�	;��]��ԕEd�琦���}����w/``��9�x�<E����[U7~D>[h� ��r�tS��0��(�����(}�[P�{�^d�B����
��J�ӭwe����R2�l�Hac9�6i��x��q��P��\�<JL�w��J��tI��ʥ��6�g��6���[������lc`r����/�g8��Ҭ-������Uw2��*��F�	�fVp����һ�v�y]v�r��T�ʹL�����:H����Y���t�[%,j&�,z����.I�6&c���Fa�>2�ܳm��Z�>��O��f�$8��X�/��������i�����%gY��N۾��x"0u�F� �ȋx/XÏ[�=v�#�Ǌ�������Ǥ�����KM �ن�����r�W.���>����������{0�b�Q�Wu�N�V�
`�4�#?���� 3p�&z	32Ujms�s:��d�n�ȋBl�&T�{*E�y��zËk]�qk���8>/h{��u3p�,?��%�UF[�d=}5���D�4
Ņ,)q�����I��e$ȅ���~��ش�E8iEi���@Ϋ̘�>�n�>�"C!�s�{���$�Օ?�]C�\恿4Q�BՖz�=�=��]s���ox�~&�c��ٰd<��/0Oe6���I%�0��8-��������Ν��_��ݦ����� (�r5���ׯ��W,W���OS������
X��E�.��)�	���z>A'����`�59�1a_9����R�{!�O�<'��+Pd�C� ��aA�钑Xa���?*����^Ы��e��%��X-9���!7�҂�_��&4��qˊ�d��F��@��i�3�.yGX�L��D���2�d��pa���&յ�O%���t�2�\c���}���1Ӑ��6X�#+<en�-b;3��9���g-~r,��ݸx���M52	J�����1# ����ĘΌ�Z��6,�sF7۵�8�V��-	_��O]w�GV�f6~��J����t��w�`���q�` _���~�<n�{�Gc�?W O���e������=�p�oD%䲿�w�l�_]�+�M%��mj���j�eL\�������B}>Әk^���5�\ �����p�ߴJ0Pë[6Яƒx��)���w��x�:o
���ntX:�Bve��<R�JJ����QԷ�oH�p��Z?e�zy'¡N�%���W�����єҨ���a��1����uǥ�n�Z������՛��W���E��fO)D�i�;cy���776�?\pe�XO�XfY� ��ܪ�@B�vy>����7����W*9/<�t��?��Lk��%&�& �A���ǽ���K�0J�!ˑ��L�R��ɴG�Xp�i! 0���