��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�_���v��	����}���g�GH����U�K��*Ѓ�!N�=�Bb��w�����9���\u{�R�8��E����#�)����.�!z�~���I -��ﹱ�Q��

�'d$� ��m��\�� �B�wd ix���L'á҄��w�_%���Z�E�4#��#zMY�\L�]�ph%s����Lb�h��-� �/����R�9��m(2�f8������Kkz�Hx�<����V�>7'��onM�k#��9�7Xי>��M�s�H�[K{��n^"Z�AY��ƵV�7�8�f��,�ov�]�N�-��k���fId����d���y��S0I"a����8�m\�_Qq�s�"ok8������qV�na��:����Y�!�I��K-�q����n �2��pm;�b�,��ʟ��hݻ��Izw�h�܊�� ��Ѵ��e��W�v��:�[�(��O�3��d�D��� L���QU�k�̽�S��KJ����W#��g�͉�Q�x
K"۱$6�a1ۆ;�#[���Ϊ�Kt�fJ���)����'��ti�A�9?o]d�߿j�1��쫩RF��fQ"y��J�R��HV��E.�F�a^�n9|(f�߫�~��ER��I�(V����f�Y#�����9� 7ፃm�ƸS���;�P�~�1/�����'�!0�݆�� T�I����v����#�Ōc
�#*���+�3��Y5�s��$&�����S�#B; EI�j${|���1�i@a�g$��/�q��_�R��z	����$�=lq�1�h��֧A) �g���@$Tj|	w`���C=�5�����<�ٸo�b���n�/���Y�}Y�}�Ʈ��u6�?`���?�\�揇8}�}F���ѯ ��K�q���Y�������p�bW/��`ֵ�l\���ls��g����H&��v�.;�����B��+�4q3n�Wؕ��WD��^g�IXd��	� dC�;{��/��I�����F��g���� @e~��w�:�`����*�jYK�S1=բIss-?&h4�o1B�^�NrK�Dogk�l����6m�E~X1�AnS�oWm�R\$�1��D���G}D�$�e^�*![���@��$}9�i3�M �!�Xp.�a�o�=��C�"۵3�f��F���N̄%���ӿ������m�Ɩ���Qv�@�T�I�Ә�H�q&�� ၭśUuȇ�q�PxF+UN�j���W�Ϊy�ص���t� F�x��"̦ߓ[�2�t���ޫy� _
�Wϣ�%�K��
�K� �������8��1V�4���(~�e%�f9�ZT�6 De��~ua�ϳ�\�1���`j����Q���H�{�[��Rf~��@ӈJ�^/g�y�>�JѼ�qft����m7���PV|�M%ȒKF�Z�
�'�v�)�/�cr�K�1�|������HM��2�Jty� MR7�D�s���r�/Bţ�������[S��0�v6��k���B;�H��|m�����I�WoҐ ОQ��]�ߑG�Fj_g��煘�S�nSx�çl�s1���y.��m�\s�rp��и8��̐LS/|��Sߜ���?��y�R�v\�/+>uu�����:�����eD��(��}���&e'�X%Aƿu�K"��$��<бc�Z,kjI�.|H�Ov�͖0獻����ɗqL��zZ�c��kM*�oI�s�����,)��ca�=�xF$|� ^`р�"��	���{��#��Ѡ�X,�]N�E�0���ޝ�G5î�}O��!�y�(��%�3������Ŋ/=D��܉�9�����h�w|O �p���;���BJJ8�h���2r0�����z�mx3z��~�y��p|�����])>p�L�Co��|pu�X�t�]�h�����}*�\���<�vf\�d���Ծ�IVx��{�z'.Z6~?����{-�s]�y�֔b�n���s��X��]���Ƌ��+� �z����_�����1��UNCZI
�q����Fo�T�GFܒ��-��	t��oV7h)7��qr��5\H����l�@vnL�R�n�@$��F�z��VA�3��e��� ����Jog�ۡ�[�^�����'����=�P�`�1�=>��_,m�aAb�O�g�S>y�|��\7!��q�p{%�6~!b�=�}4��� �ʠf|����v���0��l���u߀��g��|�`������p�v��J�M��*O����d$���{��%x*�ѽ�}+h;����h�����/Z�k�@��̠R2���\��FJ0+�
�NA��h�Ĥe8��܈�Xxtf`��sny�������a~�/� ��T��4�U/oߏ{q"軋�x �Vn�N���4G��.K�%f�����Y�0��b{
?䄏F�?e�_gP�$���bel�,TE2�X���<W;��'�=y!P����J'�i��E�&���z��H�W�a�����򜊢y(����Z��e�m ���h���2��=��0l���0B�A��F�A�@�ҩk�%�_��_r� B�la�����3��\LA�f�8�aq2}CYK-�ʜ[FS��B,���<���*홦M���1絬�����D�L��9`j�=�+�P���ES�ͣ(��@Xj��c0�����`����abqes�d<>x,��J"z���[ ���1�E|��?\/�ׇ�4�݁�b�B
�{��o{��� �5�Z���$t��Wi�&3�q��lUH�[8I%W�b.Ĵ�X	���$i�����C�5,IR�dA)�p������m/��E�쀑��YA:p�x)�aMGo6hLNq��9��-�Mn5P�W'I���Ѭ\Y�����2�W�e�b3�ҵ�V
鹬�Ik��O���z?P��x�M��,��t)>��i㓈	;e��YĽ�����������n0]���M)�'"1�a�9�?�]]�~�/�ٔo��S�����!��	C�6-��l����oюp�t�vOL�`�i��+��K@+������5��q�8	ۢ�w(��*��"����S�2�
�����<���0�[|�k�l3G� �6��D�#H&6�!L�q��Gw��X��:)s˲3-~r�-�3$�ݫ�|��o�*��H��S�N	����ҁ�i'O,�ݎHp`	��AK���4ds/�M�^�4����`ؾsb�'/n��)���}c�w��"�p����s[�̌�o.����OɤǕ!��?��+����T� K���7�Q���aG�1���`)K�۝)f�����hL��3e�����&� �R�|0�S��\��B��A¡ӱN>ݶ��bY?������l鈎�T�o�E�e<-��
��h/��o�װ�n<�VnR�z��)�4�v�?>}1�F9�ʡh3)��c�\6���<�'Siaڰ��#d�4��HI�|���ܹd�oN��໦s��k�$���s��I�Y����	~��"�,;�[�g�'��ekv��<�描�/�g�A)��%�u��PM�^��ǣ@g�&�nKj��:�t�:4ۃv�����jݠ>�:|*03{�K�*�� �v���2��0a8u��Ep��4���`
�@˖�tV���(�5b��f�m�I�l�u�r�r9l�O�&o�Z�^�H�RC���c"堫���\'	`��{)T�~D}�{h�Q�0	jR���H4q�O�sva��jHឮڳֱ]_6e���n��4g���©��m��|�����=�m4�b��d�L3cY��G>x	8ӵf�ɠ���n�qˮN�
eh�a;늽ӌ��%�;^@��M�x����`�.�Cԏ��\�]
�Zcsۧ��I��᫞�\�u�a��>�C)��+
ٽr�p���
��G�R�b%{ F�8����IP��(v�B���*���l�A(=>�f�%y�Tu������]�D�,�!`,�ðA]���-�=L�������l��+�=w���"T\��.Q��'�HA���o;�)gl�[��6��4HɅ%DE>��{�w�i��㙶%	�L��yL����dUݮI��W��과���,5?�W��i�0+���PQ��x�ڻ'���Xl�F @��8:��@�h� �֟�;�!9c�kl��Ζ��xf���@���Q��U�Ǟ��9(�&s<�L����J�*��^��Zx�1�	�:[�[��{}[
*vĊ�j�<�}�S.C�AQ乽\؞��^��a=�P>Eac���ߊx@[�����ipH�X�|��F���!"K�����K�FUXﭨ��r�ZV�S9j�/(�
����\��l�����o;L3���I5�>l^���<��x��O�3�>�}��B��0FT��b~�?D܃���3�hˏ��痟�o��� �\�Wt�|�t
������r|R��܉)�0O���A峠�F6�]���ۭ{�#9�}vn��P�~P���;%D���wl��9e�:�3{�*���-a��}����=���
R�ٚ�b牍�˭
Lh5�+��(���ΓrØs$N��E1���vh���k���� !��BmO4�g��<�b��o�!�JBY�J��$6P-9����H��-K?aF���/�J,����F�!��	 fy緶��ޘ�ƿ��s���[�ۆ�=��l���������q�CtZ����wk:zͧ������i:�kY��L��&䗺�b1\���P��Iu����&�S�~# �~p�Ќ4��'���~S�X:���qB{�hGd� ��?���;H�wn��-���"̹~t���AM�;�J+����6!�H%�}!J�('�0���[�zc�X�zk��PQ���}�)���Wѧ��Y��pj!��Z* ��82�^�з�~nU����7�*Q�v�W �2�C�>��}*4�0��X� �Za���j[��;	nH�z�U|���(]_uDJ�}���؜�t+�U?�m��@�����9�����{���p���!�����4��gx�F����:"*��!P$Yw2!yBnԸ����@���qFܽ�4Vn����"c��-w�,"�2�)bޕ>]�Z�����i��F{&Sqh�z�Ī��Ln���vm�e%_��2�`2�%)*ʧ9E���1E����8���^oJV��`�aG��Em�yXi����_�*|���ںM���f�mVo\��0+�\�+C�"0^�����0)�ʟbXbŢ>r�2��<�*�g�[LY��5�g��%����g����*ImS���|���d D��ծ+�K3;F�>�S�V�ckbhp;��u!
&� ��͖2�d� �By@x,v����AB	t�XOZ<�λÊ�e���^)�H�r̴c��#mb�xR�@�6����u��`W]��Tr��AJ����w�[���	_��?�q��]��(���"��?.�{<�߻X�#9x�A�������D���s���l���Y�����	<�J9�,�9+���Tl�6��'�D.�#��I��gzM�\}&���g��e���!�Wk3]W)']����dV/g�V���='�_�UB��6wAz���0Q�Ww0�G�Y�����)�K�ml��>�����,�-.�8Ńr�ݺ8��1�Ƌ�~����Qf��&_�}����[�����,�Y�lB��=��=�g�Yp�����1�^��05�#@^@�r�˱�Q�5l�����s�s���_�k��B+ґ��d,�T���"kW����F��%~x��0�Q�֠�}@��	~���a��Pݠ���>����э_�>k���BT�\vc��w�� S��rO��k�=� ��j� O�^2��;�v��ʊ�Ot�,m#'}c���G�jh�p��d@)�8O���Z��}жV�u���)�e���eu:q�fS�r=���_|�3�
�8��B���т��Ü�S�u����`5\T�!�ۜњ��$��,j�������U�Q�� 6�Y�����H��FI*��|�C9��HE:�҄W��M|�����c(���bws$3R+�3u�HN��K���J,p���H��9�I���1:�4E�V(�/K�����y̨$<�9� hMd4���E9�V'!i~&e5�#�o�$�9/W��v��AxrF?��&�Z�1���a�����g�rj���������"�����$U��D���^�Q���'�D�V��4F;�\�`}��V���Pjc �m-i�w-���������=1I)ņl.��MWpN֯�(����*���Hv����*c6Mm�Q�{fάE	��P*Ք�'�}�戻�R�j_eK�.����i�
y�,��i��t�p$�W�#��Z'��bߔ�%z
O�?#ʼ���u�E]�<X��vS���=uT��g*	�?�ߍP�q�t����Sa�Xp�^���k�]�P"����^=���/F�3���!,G��[Z�=�t��ۀ,�fF��j�Ȑgmy�Rs<��i�/�H=���K-9J�8�����݂�Z.��h��+����{'�_�(gÀ�o
�Ⱦ�!��%��!�Y�7Z�s��w�	ȟd"�%������t��UTS$�9�4�d˕�A{��>j���Cp%3dW�q��D��j���~H�ސc�-�{1��IX�(��
��[���&٠�`����1naA��*�;48<[���ÎN�#�o(�*Kj���M�#�[$�Ӹ;��>��&�b�Vb	��u�U$���Y��(�|��=1��	o?B���*9"�[�c�4t50d���M�����L���}�K��1�s3��������ie�I=���׃<�(�J���Tz�g栕����5X:�or���i�]���\1O7R��*<��9�m��I	�޲��*M�4��fBHc�Ut��s;��OC9�si6���}sUM�{ʢ�b�\G��ã�4(�+�s��ml��1�37`	o��^t,mjOJ�wϼ��S�*�yĆG��[����r�v�ld
e|"��9���!�*F	��@N�6�T�Ԧg5;L6�2�1�ԍ����g_�0�1�pr�4c����;���L���p��C�T�f|�ڃG���m5��>�(�(��G�`��5N�J/�S��?%�x��q�����R��|#,fD�B<��~��28��(7F���ptB}�j��`#'ٯ.��/6K�w�:]�k+:7	�Ϧ�ez�=zU����07���75�����dݲ"635�$G�[���8W.��Ai:���y+�h{\�|�D,��#��݄{
�B���r卑+EV��a�*v�É��ͺG}����	�D��Us�i�ڀ[	w�.OråI��$aZ�������	B�*k�j]��&�?�ց/[+CM�3g	RS��JtBn�-�XӜ��1��.r��CuÁ>lf�NW1B�P�24�
�~`�ꑲ�*t��(�z~z�s�� #�|m9XY���AE�[��]㾂k��N��g�(�1�t-t �n`i��,��ÑU{�o�dg0��A�+��g�3-I�(g��꟦d���0~������~�ݖ@���6���e
�h�/)`��-r��N�Ԩ���C-� �`���J��@?�if��){w��y�d���z�=�����r���L�r��%�-M�R:�^p�����6�]�\����_���0"3�{�
d��#��A�h�b������)U��*Z��Nk��צHN^�*6�����\X�w�G�ƴV�ciu�M.-3W��\Ӹ[��e��	n5�������G;�0�Bo�4F�I�����<M5^�19�G�.�C���&_?nА�ʙ��M�3�CbO�,��_/1O�����}�(
R��ci�X�`��y�c��`���()�Tf�beeI�/��|�m�� $��C�*B���ʃh�.:'�КN����!�$I�\��<��K�r	$e����	U_g�4����x�!�O�_�uy?	��r��`UY�X����,5��x��It��/���(|�7�;�]j����m;�v]��n��/�����eD����S�8��*T��'�
�����p<P�TV��eͧ� ��`�A�F�\f�D���?�ݖi����u��D�y?��w
��mqL�iF@:�*�ݼ9��&�	΁*4{�INXiT<�hG�Er���_N����"��}��}��̧Y�m����Y�B^R��x[��d�Hwd������x��E�+�$�cC����b~��7�Be�i�������V�D���rP�ksjm��X����ם`[<��썓9����r3;�k���#9N���4�$�W�[G]޶M3���� JAr]����8o4�XGȋC��8�h:O l��/�`c�xh�?�|�
�Aq/�{���YxP#����ݍ�� I�H�AAoD*/��D-��/*���y���C�j�Fs;qx���[`�ˤ��Mg=��;�QX�mi6��љ����65�:.�^>���5��WJv"5$��d�jQ���
�ꬸO���ˎ��<1:�x[�$�%
���2#�w��>��x�k����Ll��7J\�;6���)�7�)��5�	�ՋE��P<J�_�`I�?�.�%	�KbID�h{XV|w��U�M�o��}?��ׅ��40>�<N���c�������ʙK�%W"��~�h�� �g���b�8v��`*��:�����BN�75:�h�r�A㮅X`D1���Z[��� GP󽂠�B�T���MSC���$�^��9^��o�b����"ъEe�N>K燓�<����
y!4iㆬ���4����8Y��1�\�+�=�`^V8��eS���o��n�i�4�R�4 �)F`wA_�(�p�[^�8iU�p$�e����aR֊X-,'�,Ȫ�������<�8Ԅ���\XQs�D[��ǂ�K^�OL��;4�=�/�ߢb�����7Wgd�ʏX��P���1%�M�-g=�����seZ�XM�!�r�1I��(��ӓ��#9F���0��SȢ
Q�kY�7߳���z��O�P���W(�J�}�����P+�m�j%��zk����z"8÷3*����|��������,A���>��ȭX6�tL h�e��G�'�W끟��,�Dv���nT�F����E�4{1/2��k��K�9���<|[]� ��J!v�5E�3�gzS����8�Խ�)��l��,e��q�_ֺ�2�פ��LG�v�{�<�]Otxqa��"���bR�PG:E8����̅At���}Z%l�Δ��5�����X/�n�7��|�si���E/$�	zZ�(t7P��"�C��sB֥	�ZP~F��v�jMI�wkWK^���p���
�ٙ���2$�Tb����g��r�xtл���M�)s\"���.[��f?C��ij�$���̀X��\SscN/r�q�h�����I����j�5���"cY.],���N_��������-����2������ߝ,�Ҝ-��Z#��s�/���� =�䳩ajCR��Є��
���
ǡgP2T�A+�R�lÓ^����Rc���rfLO|�1KoV��=����,�?�Y��mz�_�=�T��GCZ���k�4���9�12x�ۂ���w{�J��0�UMg���x.M�^�S.߸���v�Ƞ�6��p�����P� J	 ����f�����c�Іj����1�$id�k���PP�@�&�BU���gMX����]��!������:Z� �A�@2S^k�næ`<�Q�H�V��v.��|=�i+@k3�5�/]P�{6��X˗.1Q� ����T(�y]~�H%|�g�:��@^��Z��2�H��7�%p��u&7��763@f��5�`@˨�
S�-)����#6�y�nCޙ�z.�Y�����Ĉ<UH��V�~b��տ+�:	�_c�sP��+�+�9�sgV�Hj��v��7k4�����ٿ��9zl#���ա[���ړ
L���<�o+-�gr�u�yM_��Rg�E���ԭ���r=��>�ЀB�z06���䮡��4�yq�I���W���X[ly�@���m�(����K' ��&za�L-��(���	V̑ډ}o�L�m�F>~�����Ng]���,{7}1����K���ojb�[yeh��GA?d6-��!�m8�5��Ҵ`���Y9�"7�G"��P�ɾ/�X4+�A
٭dcW�%W � F��A��c�7#�0=�]�DL+�WI�F�E�k{i�2���)}���(a��{�a$R�Ӥ��b��w_:]9'��Ё��[��+ܸ<��X�;Q�'Y��J��𶒇��ht7���y炎(�"��Nqa~9S����:�S��T��h*�-^H��K]���T�n�6��!�=x�( F1��[b�.�Q��fw¿jN�G=���X�� Λ�{~6�-�"PX�������;Q;�ko�To��x��U(���Za�T��Z�6X#�����[�� ��%`7�<G8z-縹R�C�Hw��N��E��y1�]����?��>�� ����X8��ݏ�o9�^���@��~&b��eCL���kN�@�Я]�J	��x���{���<>MTCE��@��|�pSkQ9��q��i��p-�����fx���y���U�k:Ӵ���S���[~�[Fp�K������u�eԤ	l����a��!e�A�cd\[�Xze�VȽ��/ڷ�M9F����)������{<-$�OJ�7!:Q����>�L��)���<��]��������O�M��81�/�T��0c�`ǝc�zdb7=�Dq&��H�Wi�Dh0���[���@�ժ��QD����R**�+�|�#��9�CP�Dy��!b[Ò6���U�=��׶	Y��Dx��Ͼq�Z��l.�0L.�K��>��P�+�WOM�_��X,�Qz��ۓ���kL� �1�p��{C���mQ�Ӽ�:�;5�����[D\�P	�K)��+z0���3M�6�hq �/|G_��"-�=5�Ǧ��-�cN�m���U���+���ҁ��]`��M��3>��)�W���B��h�D��A��0?���	��wς�fÍ����U��)��`P�6T�",�D��-J����e4��)R���+j,+r_ql�X��p,��6N�+�_i����*�КsP���%p��K���u\&�(F
�]��(,�.P,Ґ��'�>]F���y�k ��W���8)$r�u��@���Fh������a,��w�2���qSGa��8���P�e�&L�YiҒǊ�/��ȓ񞟆Mo��:�s�T��	�6���7���b�B^L��'��[�ʹ�=am|�n\%�����*u�Q�a�)#�|�G��nz��!��ز�µu,e�Y_S���BX�C����j���m�u��F_�����sX����̛��E��8�&�Q�9������Y�;����e�~���6 i�J/^[��� ������E0�ו�Y������X`�B�����B� ���>ȿ/��W
`A���������x^��zh���>vu[�L���˖��4�C��'ʂ��zՌ�@����{�q"���A�Tc��9�I9u�9;�&Q�B�	�(Ld�.B$e@���R\� �F)�P��2���"�c�� l��9�pL�Z�1U6��ey��׹�M4lt�fDx9ؿݕE����|mVyC��*O�/��md�QfE�p��(O&D�=�W�KO��[PދF|fu�TJX���v�E>­�GG�<�9��G\n�b����D��iD*��"��7����T~� ��w[aHxtl�!z9�5x機AKS��:]�n(K7Д�X>��.^��?�Iny�/��@�Y�L:r��zv���CS�v������^(T.��o�T�̸�(L7���Cإe�̑�[�p�x�k��:��"��nu�����&!TB��?P*<�N����KF'�@	l���ԗa΂����)���������#��$����~0I��(�_�Չ⿰ڢ>r'3Z 	���,C'���djϴ��-2�aP�f��MAR��1�\� ��i��͖�T������	F��T�-�25��* ���n�4��\o�25�3��dP!w����M�9���eЭ��јЏ'���X?�����ṿ�k��`���Q1��or�hBӒ����̽���9�K�єA_۸������ķ��u%-Eh;6P@�`h~H�6a��,��:�G�����P�����~<�E�l?=�8|%����.=�,�c,���Dg�%�-���8A�,N���7ٮ�z�D�~�fVJ!e@)؏DT#�?�v�6�vK�T/a�s���eH�[�jm�.� "p//�g�ޑ�j�%�Q��k������L�}��Ͱ!���lZ���)>M� �a�� }��i$	;ؽc%Th��G�'ր�|Kb�=�6�\��J����*`�b���fB���:�g�o~�(��7���Z����	��J�f�DXu:�e�r^�Áy����X�d���`�!��3B"��[Zr�ó��@�E�B~���p��$]~4i��(u|V���O[%��'��%���0���	�4�
�C��^�t����U#���
��F��r��`��y�����zE"���ݵ��/�K�/{W[���M\��z� ��kJ�ю^u� �Z�Fz����X���F=�@�L���O�����Sa��o���yJ��Ъn��n��0�h��A����c�v��f!by�O	�C��\�mi�u����+V��i�C�Ņ ����N<��d�Š)������Efb�}�K�j�%��9c��e���	=�>�6����\sB���i�\��>��p�WT�[�mk��L�޼@��:ܢ	�n�ب�r�DoT��%Gp.�K�c���X,�L���ay��D�θ��$]6���u{���^�|Q4.:ڸ$��[�']V��R��/g\0(^p��?���I,y4�S�}�:���,�
0�_�'�='kʟj�a�BM�g�[$$T��l�Q��� �R������b���j�JU�<��-����zf.��h�r�/!��b �o(�I�vkY%{�#J�Y��%i�3ܿC��3���RfC�9�y#t.*���ի4i���={�!��A����-'�$ �����/��C�ؙ>�L*H�p%�Q^�Ų�  �j}�ܚ�d��{���g��4={F/g�� ���/��>�}�!��#�3�ޑp���d5QB�2u�;5揊s��g�n���:�+�|�eZ��1_:.�>}ђ�6M��P}�f�Z|��h�O��&|�:��
�cڄ��K���p` �b�Q�1����~�-o��?/�}�d��j��>���٤����͝w�_J���Ѷsӝ��_u�Qyܱ6�{�4�e��u⃨b��,��ӼO&Հ����z�O�&��w���a��7�ո/V��~�����!Ƌ�����7��DcRCs��:rd0P������1���4�nc�Xk	4�%O��e�f!���2�R�������I�����&��u�_�)�%��a�M	����s�U�aD+���V��zZB�
�N;���BA��a ��8.a����C1@鮰��#� (u�>�)&���3�/�%�U�G\f�L��&y�h��(��ܶ���m�s�IE���r'��J��#,�@�ߤ'p�ig��SMJ���S��p���L��?ԙ���^7|m����o*aCڶ���
�X��Ʃ�rH!���c�]���z�5`v�>��:�u
�ϒ����yqHj���;�)`��t��(+rT(��������)�+���fҝ�t��S���O|E(��`�VB2��bOS�c�X�n|sD�.id=��z�.8����~P�&��7[���Eˎ!��Q�vu�M��u9���\ď�H@h�؏���^����Vp��8�,dD��W�����ā��1�0B��l�Z��l�˩��#(u���@��Fz�T�zl���L�v�_Kc|��������-z6�y����ݺ�$ ]!�=4JiĲ)�rm���.V�I�g7G�*��?���c&�xfv([2�����Xڼ��� �Y�|�0pD��]�/N5l��B�9Z��մa`w'�(v�Q(U
�dY�G��T�5hb٧|'���f[j�p���[8��R�34����n��2�z[4Of.��3�l�/�Oz�i����_�1�[.<vi��{[ �(����'��Q%_%��m��,�1����F��(1�;u�T.B h&c�k�`d$w|;n�_% 00�|�*s�ӗ'��xv��XkJ���)�v� ��|$�X��h���ސ5G>�<��%��~��|B�:�P�g�tó	�5g�����ٞ���2�������U7Fz)�/�#�o����$��2���%�n	,�8�"�V��v��Z�o6й�7��1�P�L�#BkS��$�,�&�M���ͫ����.�į�Q��,�����k^�)?�MY��N�z��n�jץ}�6+^M7���Wέ�������9Ozx��JvEZZΔ'F�&m2�S�P7fT����d~L,��/�?��k}1��·�C�S�A�^�,W��JIk0�ɣ��b��Rǭdo��ϭ�@;FM~�^��
�oާ�7���֭�I,��#A2����c.0&:��M1х��4`pѯ��S�ku�5���ϛf�2�>Sf��G�y5k='�>t�s��/���e�����`'A)j_�9��2~q��J���ʛ�E�|X��������|� ��A�6�F�����EhδFPܪy���F�6�zڣ��c"���X�~����xC����;F�1c�ˡhwM)	;Y�!r3�>e]�;�&�r)vґ�gC*x)*�#c�zD&�1P�2{=�m��s�^.)�d��F{�J	����թڊ�#-):��GqԐ�j�LY|���f{�+A�䲻S�ڳ��o���N�U�����B�	5��B f�����y�:7n߫�
����aW�R�����is}�Ѕ�|��6:�!�p@rF~��!>���5";$�Yc�Hb+7�"-���գ�ރ���q���ٗ���qeD��� 韝}`�����N���#�?�nh,+e�O�̿��f�o��i�7f7��%<��0:����*�d�T�C	LMP�������`&�Y]���>b.�U$hK��l�0 X�Z�g�x
���z��W
���_��#Kd*r�h��Ș㫵�N��,���p������0c/:�