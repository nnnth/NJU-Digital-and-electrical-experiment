��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o�:!�Q$�d���d����B�6H5��G�=����?���G�R�LvEf����n��,��c��\Y���0~F��$�4����ࠁ��W��P�ˡ�8c���C�EKH.�{j�x�c�ј:��DI]�>R�ɶh�&l5o��f`����K��c���&A�y�u��D�c��:�	W��@��J�*F,�@ồ^$�d!��q�����^F�x#������ �Bdr*Ϟ1@���&({x&�/ <���+�y��4y��lXa�XngB��O1�fd}]C����g"�7��s���J��|�4ͭ ��0�g��B^�v�F��#Y>h;!Tu�~���R�7�S���q�J�snQ�($��?���fjx�*�!H!M�(�~����[��d�'E�c�����[ ]S�}9��K5E �λ�]��2�:׉�6�F��; ��~z�x�4�u}C���s�t����=�r�;U�,�-����[�$p��l\��x��)]�6/|H�0SL�#~�-���Sl��V�Mk�عt���Vۇ�K~Z�q�}w�ٛ?v�gB9�M�t���h=���WKGe?�E�2/�{ �ۦ�?���l��>�)�"6�Ր�v�Է��=���}9��yJ\b����A��A��QBzV��P�g1���0ٚw~u終2̦j������\O1bcC;��ʗ��\��$��_�q��oEU��DW�A.����`��O[�<��-�}��ʝd��^	�J�~0Wnv�eVw|T��D�����`� �O�Ef��?t�-�=k�t�b�g��p7V����G}B�0�{�l�	�j�XG�v�.U�yLn�H ��w��-I��VN�Y��K�s��F�@5��@�� ��w�~������7~N7���r�(��v�� �3�W\JA��qh-�iq/�j���:2��(�u�R���ۖ�?/9I�?R��N��&h΄����0/��Χ~�<C���Fj���RӵcwoVY�Ѣ�B<��'(��٪��p$Z<c���b�fS)şg@��U|��z7�ɱ��Ű� �Ss@�+��S���՚�j(9�o�}���_��.=K�D�����&�h��{���]3^�;E`م8�6<���t�v��-?1TX��NOÌ%� ADJ�31�u�I�oIR�sfnq̂��g6���|�m�	���K�6-�J z?�=#� r���u۹�U2 �0^���f�j8KQ�6~BTQ�k���_8s�Q!`j��X7�VN�����B�JG9�2�;M�E��UW��k�g�mQAF}+�B	��ŧ�21n�z�L�ʍ{z�lR��aQX����qe��'���$�&��~%��?KUؽ�2��;�G*��f'x�Q��!���J{���@�k�����Q��w)�T#�(��A	v���PDB=hz���$�A�$T��5����0a����iQs�4����2)�9����������p�q�u�|N�OZ�|�9*��� ��@p�L�	��~V2VoKŭ���S)D,�97]f����1M��>�4=,�g��Մ�Ln�7��n�G- ��C�-ߟ�m=.�\tSUG���Q�=]{�^���9D/Ƣ�(XA�M�����l?me?��і�_���)&��u	�b��c��·�uv��%�p������C��5}�K-�`�?�u�~���!���V5;N����_!�p] �}
>�,B��%�IR���� �����s�b�)�ա��r��X������S�J5ы
)��j�#X��ϗ��`i���-?�́�ь�qf�J5�(
)|W�W>�\�qla�k�W�z�����egF7"v�ȿLD��8l3�;�Z�1�`�/��^�,wgד���
|��'N����3�]T��s�:�?�/�%d��T���4ȐÄ�����m�����d OSF��d8�bW\ʶ0sF�i�tI��a k. ��zI�+��]�J//��2��nE�>4@R�Z�ǛxX�#�]����N�*&�3�st�?���O���)?�R�1�I�R����+ɝl�=1�A�i!���D-�{��PJ�+K��U��t9��ٰ�)�x\Ɂ���4A$:����9 ��R��oKD{0 {0$MJ�Y(\W�m%��&����_�?�f�j�Kj��J��i�4O|T�Ut���ZѠ
�15����P���%�!����Ta�rT"h�00��6w�}����2�x]<2{���77�ES���dߏ{��ʈ�Z�S=�㌷|Rܹ	�O�� m�Kv~�')=���\j�XW�'��!��w��՟Na������ۤ���<�t����R⍸���8�I$\�o @{Ta��A �U�ȯ�y�eƇ#��'�5{�HU�ҝ�^G���I`a��Y�<2El1ھJX�{���1����B��<�-4q�k�����9moV�4Y��;L�x��qeDi���ϠV���
���49I.V�1?�`e2ىy9qװ(�g= !�2�Ϯ�1�X�(�����Ab���u8�K;�=k��NVo�ᴟ<Nnq���J���צ�jb�3u��@"EG��d�Ry�TC��dÙ1�ëJ�N*2�LX���iɜgf<�)zOF�H�~�����I�7�ַJ���M��eDE@u+ݲ$�)�ʙ�<ȓ���nEt�J��F.
y�������'�R�?ѧ4L�Q��6'\��DT]��0�7X�FJ�*���rh��	����P�"X����W >Bk�^�%;f���+�R�c�裡&� pr�
Ux���T\��B�f��Fxt��y4b�w6�v��"1�`M>�C����@��\�U�r	Fp��5&:V&jd=�1�f�n���y��D�7�6��/EΝ��}��Kn��dK�/���M���y1#Y��t��঴mF����7�nV�H�2n�i��L��%��E�u��9+B�\��S�➊*w9����M��XY�@�Lr�$zU�mPX�@J�K Nvna'�e|�ڟ��s�^=�&,5g$:l�1�{k��0k��
��u�s�K^U�R�Y�ˤЍ��򓧾��n)ym �)n��!��	�B���g�hAdB���w�jϳ��ɀp�2����"�k=�&Z�y��0ޫ�!sLeR,P5���ħ��&�hl���NB���/�ڰ�(��5o�VQ�r~����]�Ľ�O���v�X�4&��`��;��EO�~���	�Ԧ��Ɉ���k�n���#k(��2�l��5?����T|�w�E�!�n� �`Fv�5[�L߇��\��6=a$y��Vܓ�ɍ��.�D˔�_z�p�id�5�Y�r��mwWm������CT��5a����@��޺�@c�o��^���>!����_�|\vC�kq��d��&��+���u������i{
%��gÚ��2�Qm�1#"m���+N��#od��&�%8�����ݺf<\#rf0fH(.������Zj�XU�2��6(C���su�e�&�I��N�a�����T��V�n�99t�N�?��U�jD��(�?r�6�[�ͤl��hTMu	$��"�w�ܒPPY�a�h�t-tq�`�G�~\��������B�@/�FY:��g��T8�Zv�;J`����Y�4Z����Xڷ8�V�R�ѭ�S�i0'�_�#��D��E�:a�.�fbDJf����"*h;foh���@�^��M0��K���ADD��o/���YcR�,�-���-��1�R�k�G�J�H�}]s$O�8���#��D??�QwLq����.��|vi|�L� �KuL)��Gb�mPd���4�_Նw�����Q��x�}��4P�Q5lK%]Ya��ӯ������M��ٽ���g���*a�� �k�]���v[x^�?��{N��.r][��C��P��M�0F]�l�H��T�¡_�_�i�Q/ǿφ%b�d��� 4M�ZY��P͔�����
_���ؿ���?�6�։q�F�t�n ��b�LG�(�(��˙����ޤzS���|+�I��*ɵ>w��3���Y`G��i kQ�Ż�\%!#��S[��p �:.8��Ӫi�h��ƁM�:�eF�U;�
e1�S �ؽN[�P�S���ㄤ��,~��.z�ׄq%� �{�d'� ��_��W�u7~��cA�1�aH��H@yMs�#h��7�F����Uׅ2s8f:R�}����yiQ���/ e=�����$�^V2oQw�u3O��WT����M����p}����d�g��6�����'�$�gc�mJp��	��fzQ�,#�n��3ӳ�^����r ��q�S�a�M{�*����7wo��Tv���S�	�$�p�L4��`P�ވ�<���ėF������!U��=`>_�e�?�|�"Ѝ lJ�T��~@ܘ��O�}����$�u2��|��{ ��g�}�[�q�+{�8%7��e�#V{��a�qߤ|�}���]�a׆�sJ(��� ��7E~�mzXg��d	���۠<ԪH"�ǂ=Bb��?��`GAgv�S��5�M�֣��T���~g�X�O���	}i��*�G�t���nC6?��(0I�Q�����:.��8�W��W	`�4�l�?����jԻqƅa ���p(�(�c���!X���	��5�΀�iqQf[&�0{�}���/L�֋l�-i���k��}߇I�|WJ��2����䬓���'DL�r�W̚�ZNr�t�b$δ����h��G���{��D��k�[�����D7q�������'�U����U�o	Φ5�%`�m[���� ���b��L$��2�17PX�&�ar��C>,����b�'�Q]y8B>�� &�����)ſw�ko,ނ⧟C�><�.�����s��A�]�����J�zR�U5$
�K�2���*un�Xh^�{�G�1�vN�&.�ߵ{��ʟ�xc��b��sUp�S�q�5�/��hbY������s��� b��A��때����'��ܞ�`��oO���-ZYJY<T4�P&P���8�jp뾨8}�*��^3u06�@g�ڀ
�S;Qg�@"B]^m<���*/��:u�U4���y�䟰�l�����#��4�sa{�Z�4`A`8�~�Y�N����A���0��2lFm1´D~�!n�-�d��L5�[�|jwТC�i4�0!�nD�K7X��t/;Ru�z�}�d��=�z=5�qi�qf�"��**�4����Nz�Ѷ[E]ϟ�lFa5�ǞEW�ߓ�ߨO�/��*s��硝1p���a&J���Qutk�^W@�1/Ej�d�3K gh:���7ɧ�t�C57��hޙ�{	����%��q�7��,C��HQ$QP��)\��/]�R%7��/{�*���x�~�1��E5��#�
sT�h�M)>C�3�x!ɢfr1���/i�e��¯Jѩ�<�E�%��"�Ħ�yұ���xP������a�Q�ߐ��ތ�4��(�t-��Mu��|�?�h	�uHJ��(@5�>v��X� ���tSL/� �J^��>y�j�\M�£��}�KH��R��.��gOP�K��9C"�P>NM�
�Cc{8T��2b׮!~;�W�v
����֊My��#���}P@��D�9���w|a��iva8��t�ȏ�h9N��%���eU�jDR�n��|A�(��@��[|��Q�/g�Kx�_���6�߀�
��(T0��6�m��DH�naE�����d�1G=�dL~��P]G�
~��˯�`�`5�"O�6j�37Z'$ϓGВP����L�3�5���E�hzW)�_sn�\=ٺ��i���[IH� ���p�}�^����[lGɸ��K�;~ �����&)Q�ɵ�P���3Z��R�R��'!���2�
���,ƢA�(�7�吣(�	�?f���ѓ�s(E@�����'�!�PiG���$��a3�z;�;���;Sk	Z46YG������^��/��o�{>>>�n�e�Q(>ʭ��No� [�ht�῟�#���� �����	�ؙ�P�	�x���VH.������^���@�J���I����>Nl��	�8�#��j��(��u�R�MY&J�K	��N����~s{A>�_�1�׵�Ø��-�Os��Ѓ������x]GS�س�ĩ�2��䤓c��1Ġkt0P�'_��R�z����"y��[^����R��ك���b��S��%�=���яa��X���m�sG�N������gA9��c�)��0��z�i��T�б(�����k�:����B�w���5	�8��������Y�0��]�ZI��M���r�6��{�2G,����鶆#+H߲���h:��u��ۿ[숲�����$`}�S�*i�J�Q/aΞC{2m��h��U �R"­H�Ka趢Zw؎�D�-�dܺ�W+�|.�� 'B��r��|��k����d��bU�h@|_���[j	��]|�he��d,_>� �����G�� �|�1���24���r��#�!��h8���1Y�sbW�<���,(�>gy�ԞF)t��?sݤ�?3�������C��Z(��1�<꓂�G*� ��ry`
G�������ht�M�c[!Ϣ�i�"l	%�0�w0�]�Y���Bh�[�0�����+uΩ$i�7��
g ~��*dM&��
�c̖4m�h�x6-��N=�t �p�F�/4;���zY�q4��<�J���pP�k٥ꘌGm��7W۰�yOZ�6��!k�����%6>�C�xN#!'�f���Hڄ@-�x� �j�i\�qIcE4E��嘊+ij�]ZWC�4km���%��c$u��v�.��h>
C�s�I�����a6���xu�Q�/��֧�n��o\���DbV�`�]�	�B�K&�-������<�$!#š��D��@t�]��w���c@�mܑ� ��VSu!���������.����9�ȿ�z[x�A�S�9^MI�g�v��)b<��B*�7��T!�ee�/��]n��)��߻3�� ����A��!�I�������Zd�8���Z��=�x����U٠����a��ky�>,��;ܬͶ�RJ�\]��g�ܒ��&���wF�ez�"l{��w )(�1�|�7J�JVt�ȸ;����7�jhy �l[�u���Q-g�w%p6C��2d�����N79�4���׆	.�x�������X�^Q�;喴�s|+F	�C_��Ϡgv�x^y^��M���ב�������^В9m���da)��`S�T��:U�^���p\Xd�������h�I�c�<?��:��6d�)zG�2�
�`�#�w��n/�؋/��y�6$�g#LS��I�I�zl�B���j�_"�R�4ʰy��
ƀ��cO`�_��E��#�ABi�$G2��5*f��v!�`l����ޱg��j�AKU���h��mom^*
���;��|�R�ʫ�S��)�]�l�oe���ʁ�:x�q��������,.SG�_�����Y�e��Ho�~ۦL��������53h%þ�m?�װ�����D��V��И���H�/0�R͢�]����������X��b`εn��k������9������=9/ ��M�����O�yZr)������A\�.g�[
*DQ�dk��⏂��l���>u2L%��\f��FŐe w��A�z�$a�����Z;l1;�{#�lu[|r4�}tsC�1�	�9��l�7�m.�=i�?/�nЧ�r��l�QX�]����ݪCv�!Ƿ'@�B2��O�X�BN�?^�y��&6yUay~X�sg^`!�{�.A���#�7#P=�f�%h9Gb�m����@�w1�J����ڞ����F�;k�Յ�#��W���b�ݮ�bHI�u�j��Y�x��}�'�wa�����m!��t��+���:���EM��k�\=����,��w�$.ۑ�_�|�Z�y�^r�1�4��}̮�,5���ϊ��y�ԭ����<��/Q�k�w�JK�k���;kX+�m���0��L��$9��Hv,��3�	�h�� ���mo.���A��*��GH`����gq���n�\�D�t*W�jG~���ͰS�E�v6��8Z��(���`$ɂy�ѯ�`V��4�_~8z��G��5�Դr�D��;g�PG�m0�.�Y��N��lo��6�Φ-*6�X����<�Yѕ/����\�+<�kR��yjw�E�e�t��0�����T'H��QzN6�у����oˈ��q����\�L>!�@���6���9G��������� �^��20"��I��\�F�9�$m��&��������I�R�f5&lc��Z-� fL�w�PZ�E����~"p�;\�?ۻ%_ķ%b���Y�Odk꧙$T�o7��AiZ|8�5��+��l�VX0��N<.�؆���Ҋ�����񼨜-1��Ђ˂E��OU2�Z_�=)�ؽ�LS[��k#�ǹIIj�݂��Ŋ�׊�$Wߡ�(�G��F���]�3�>� F@gOf#��P�Z�9�H�i�h�d� e���
��"��{<:�EI\��O��+�[��}�5�j6��D?�N�q9W�k���K��4�Bc�w�pKƦ��˃� 6���7��%��
�����\���d�IZp?-��n�s(E��1�4�s0!V_�z޿˪��WH��ރ�aK�v�@S�  ���������[���Nh(���]�����M5R��tz� ^Q�#��:��"�'��RW����8���� a	3�� z�#I�;�8).;R	�R�6���ߠٲ���:3ac�$���%����5?Tĭ��U�Z#�|ƴۗ���(k��3��&p��L	�j�.S0����sr��\AQ��eQ �b]�A@�(	�ߘP�P���οY:�Q�)܁&f��7���m[���܊gH��"�P�7�4�A�`���/�������Q�Z�1���?�v�"W��J}8���<�����H˸y�u�c�Z�'"��P�-����>`5l��[<���¯�(�l�W�ikLi�;��I;����sOx��M)�&����X.;�%)
���E���33��ݏ7:��oj����T�]Sbz[#�r��]��<�%�Ů���]2�W:������ؗR#�,\�/�8���E���)�sn=�3�|�}�F1Ԥ�X�QK�(��x9�cJP�H},0\�#��-7�m������K#rG�"�@V�h��E��͞�U~r�����C��	䫸��s]eY��o�����w�U��_=��|���'T�p�L����|��T�?�q���I_��OJL�N(�G��#H(K��~��?"ac�z�y�?>û�f��������u$��bmiS��.��:�>�¨�y�W������� c.��9N&�))	X�P���dC@5��`�z���g �1S5�x�Q�.�鼫�`?+.�X����7��ToJ�o�\��
Q ��$��Wa�O���g,&w{t�� �Y����X~���A�����~��L������;~zJ'"��ab�֋��"B����s�I��T��3~�~��Ьĭ;����������ѝ%��J2���Q"��R�[O���ߋ��0$M�1o��ʔ�&?�/�Q��S͕���
���qtO�w{d��)^�!�x��h��5m�/j�>2����b��ĜF{*|��j�ިf�O���ܝ�����K�16U��t�Q��|VAo)J�xN"�E��ͻ�Y�^����yf��Q���T�b��7�`���WEx��9c�i���3^����&i��A$$Z�ﶌ|�R���=��G���b�8ڛQ��nM ,��}VĬM�;$�ksqă�%7nfפ��"�l�/p�6���"��8̩�"�*r�PR(#�+3���mY����������˥/��ܲ�0�N7B��54N_f�[F~+r�@>�	f��{࿴K������{P��`x����;�l���<��:��ak,�k�-�10�ǭ���~�8��m	��+%�Iw eObjPL~ժ旯�R���z�p�S`��w,+����_�+�/��t��ȋ�+m��iWa�F������Xg���
h�D!#6e�ͧ^��U�v�O�i
8q/��kef��ĲwK��dEba��K�V�껉��)��Ϫ��ɘK��#H��}��S���	򨉖6=R��\�	Ʊ<��S�;�?�'��+��j+3��c�LI���2�ڡy�k���ô0����� ��� ��D#��a��*9���Um7�T{����a���va/�^�x��[�'Z:(g�Rq���$&Jhҳ�n|v������u���}�W]->���jHωJ�K���
e�Sr�]�	�I����t�
XE�nկo��܊h ?㣜��_SiP���}��J�WAJ?�=�KՂ���8��Z���`7_����p!Z/_x�wT;��h��[��#�$/�ɽ�~6�G)��������3@�D�m���:��ؑ�ɛF�`�L�5�\:����R���y��is'�H���yXI�Z����?w��߉�oԏ=�=7/�K�"��^�s8Н��0N��ɶ�-���/qͪ��wS�e�[����`�s���`�>`Ҹ�?XU 8	��ٴ�h���+'�|���/���tW��{A:nGr���sӶ?t9,:W�<m����J���;+�r��?��e����<5פ2��Y������A�W���w��j�=�����$��e�3�
I9�<Y�[��F������7c�G��}��r�!CA���c:P�=��Q���&�Op��+���cG�:� l���.��dr���=#e}������X�_Fa��=��ġ�26��U�+�gG�#���쑣������PR?�0[�Zq¨����\<���T���v$�p�F��#��m*P�u�ٝU&��~�c0��"���.BU�c����,(�~����0_X�R���_�y��gxࢱ]��iRt�sD�u�0O��'Bl�zHK�`^<<Z+ܜ��n,2�=�j�v�ȶ[�r�rS�����Xf�C��ۇu��>yY }�h��B����O0{;�~# �]A�����[� ����[���y�7|2��b����t��[��r}|�ȁ� �Ma������{m��$~��G��B�A�(�Z�T���X�/u�đ��U+�"�AA��/q�}X�%���1_�9g�1t��<�=���K�:�S��߉i�`��"w�p�#�Cf�Mf��LHu�AHYÔeXM�̋�L��=�3��	M�d�PE��e��q�N~�Ǐ�w?��{��F�|���;g�o�=F;��#9*��]/Ss�.o!sl[�^,k�d��T��l�s�]@�郞��Ǻ<���1���<�d���v�̘��nE=ʒ{����L�V���� �b���ax
*����~��\������kV��0��������{�Q�
�kC�Pr`���pE�&��c߬���Nn�V�{�I#K��-^]�	������p:��i�r�3����6Sڹ�\07�'';sҾ�4����Ҝ�&��-�(���mQ��qJ�.���Ў��^�C�� 

l�{���s���X�YWk��\3��ӻ�lL���Pȕ�i1�;�>w��C�۞�����B�H���]��ű��_��l]��'~Q$�^K3�ީ��_1(y���� �.q��܂�FJ
��]T���3Ċq�t(��kʟ[�7��߾�Y�"��\�:n���y�Te������@c�a]��¸CC4No9u��.f]�`*�o��&\�O�)�`F���8�F�#0:O�V䧰e7>[ŗb�W�/��FǑb�j�88X�d���Pi������\�R8(,Y�w���eۃ#l;�H�K�|7=��z׳BjB�+�P\k� �K�����m�P�8�5s(�
:LZ/�}2qb��)pB�6�u N��s_H�2�`�%��WPp�n�7*B�!�-^|g�[�iJ��G~@�p4�k8�8`�d������|e&�'�/eIo�]��w$��ӎ�Ck�����
u����˟8k���Pu��RV9���Ei�fh���C��F���Y��Rh��Ϳy<�Ԋp��[)�px)G?OW[�	�3�=A�+���%�����4i��kq�!�Y���_{\?l�-��
�Ͳ���-CR<��L� ���۽��g����n��WD�B��`Z���j4�����<+���Ms1�}�����`��t�Gr5ՂӪ?_=: �� ����-��%C�7���ݒ���t,p��b7�"Z���`��N�W��F��"oCn�"�ʤs%�Z֪��T��$��?Z�Q/n�����:��9��I�>����/
CO�E$�����\[�G4�za���'��=�]V8JR���ںgv�B�w�8{8SS�e�K8��9�;ӗ�^Na�f�*خ҇�U�6��Z���C5p����$ iY�xO.T;�W��,���|�vCh��q�����;E��E�p� ԦO�O��TW��+�I �#�	�V���� {2=�,������7�}��|枷�y���\�X��Fi^��ĳ4P��qV�����{/9kJ��#7�q��}��.D2�n�?xL��kn��[p��0t��C����J���?pH;��(��8�W�Y�4��ƀ�D%��K���l���%6�~�(�>��$s���i�1	�qt�`����1A!Ri!{�IT2nk��\P�ř����kRLQ��%2�@h)��S�ʰ6w�1n���.��zA�z�;8[�IUs�ƍ����3uL��%/EB�k'�*�}"��(/H�����I��2�=�\��%����(�H;]q����}6����N�"�.�#�?�%��&������S��GJ����[�O�z�\g��/�d-,�m�f���]�ضq�A��¤�h�.�s�c�n� ���V[�m���_�J�E��`�1��������輾;?�������}h�:��B��uK$���))o~ ~�#/;0P����ӟ=�I��*&B����dװ�c�b�Q�ӆO`���@�����8TJ��|;�c�zQF�-���Xi�Ǩq�)	
��C`{���S�.�J�?����[�B�9��9���:^GaM���-	m��c����i�D���n��1��gu�d�p��l<<-s�'(ԫ2��n*U�r�܏��F�>'f���E�e<��
!�r~S���w��U췝�v�о٭�V���I�eۇ�H�

-Rm���1��v��2��eZ�*���k�� *�sw�f��V~Ls�đ�Z��������)}���k��ŏi�ea0no�m'��\��'P��N��'��^q�Ψ���0�b�Up��W{YQ�TFA{M��$��{��,�M.��+J���Id�`� �O�'�+o�{g���=���Y�L<��s��O>�Ϧ0"J�[M�oL���!���g��EL�?��@�(B!F����H�{&'=ĝf-^�K��7� M���{4����S�&��`���}i�E3��x��-_�'�E�i�Hr�&�P��ѥƌ+%�*;�Xk���-1�N�5#;�PF2�c��Յe<���Ӷ��`50�I�h���@���F7�X�v�5!��~E#PwV_xG{e�j��Q5�+�H�����o�Vl����m��Z�>F�%iJ펤Y���-\��r�q����
)��$ؗc��x���^�w r��̵�<'���F���3��hǏxt�F9k�����?I�#�������T���CW�����z��+{��Z|
M�<�֯��+����a<��U9ւ���U(�er�EO��@EG���L����Ø]f6�E�:,�_� xt�Y�RM=�q���7M�%��o)7>�Z=��������BC�3�L����ñ��^-K�Hu�a}�����^��#���w�:qɌ�D�~ځ4�l���j\��$Y�3{�<�Ew��H9s�� T����L[�N�$�W��Cuoh����?1Z�k����F�v0�mI4$rI�=c,F�c�n^2��8�t�96��3@�� ��JS[Q�G,�Bg��
��b��s�ց�ǜ#5�-��r[nv07�׶���"ę�J=րXJ�Fr&�k��GX���^��"�2G)�:UxN��"c�e�诸a,���B��{��qr7��M�T0�6E_fz�݊�N�ñ��ͼ1�0f�ŝ���?���-�/D��nh��(ښcT]�d�CNl����i++˃�9?����%~2��:?UϬ��9�h]��I��I��gA#g���4XM,|蚜�R��s��f�-�e9��;�8�<^ϲ�<��R�\ ��H2�W�zu�����´[�"7Lwm�f�G�5����sV����u�?y�ohҙ���A�����N4�m�N�{!�����!��՟��f���3�G�'֭._�>ݤ�t�} .��P�AŰ��"��F�6����4�vW1z�_b� -���U9��ЪYh�I�(	m����=�6��)TA�L�A��qB��RU<XK��Ѩy3�I���uH�T�e��-Ui��~>KE$�<M��g�o`#��a:��D�{��l��ڌK����ob�tS*���hA�
x��6@ٟU��ڭe�a�m�91G��$�]j���}����:�b�B�w򟻃���
��Ë���oC'	�CE�9���(�oW��8b��Iٌ���4����A����	�Ñ*�	�	'�7̡���S�E²gl�1��O�lRy[,yӮ���S��)����	�7Xې�_6�����eTt=�C���*֗O�ak������}a���C$���Fi�bl�/vr���J�Gjx���aM�K�1���j%E�k���М���"[<9�󑓁��e�_�<$o�Z-*�j]����2T��{�L�g.=��Qv�j�N�t�I��W���G�[�@��]yWL�d���8���+��9��1O'Oy�i*�⧠��6[S.�H .��xH�J(���pB/#1P�3<fA��>g�92�^. F���vf�
Y)w��@x��lR��
�{p�+��E0�Xkk��H[{�?j&8 y�ڄ�o4@�HC��g\�+�x���@�A0xQ��+/bA���4�H�卷Pr ��rW��b��KQ�(yz�\��[�rJ��U����C��:���;�%Z���j�P;GA�'Ѵ����Wg�QL
ߴ���:|8U@�=���	��7e����z�f'oD��ъ�h�U6��9�H$'|ڈr�(��7�BMK�~�{P��@�K1��!���"n!����eC�IY��`?�fB>]�ǰ�5�$�j2m�C����Y�έ�SH���>�x��BM���5���a=Ѳ�Qڸ�{�MpP��y�z�1�O]E�6� �&m�U}��շG��Q����ǅ����֑Y���5?ؽ=��'��xe"����z���QJ���C�a�����=��7���/#y�Z�{$E�'�~�Zrd�RHg_zc�	n2��_c�����D^6p�~̲'|8��d�B�@�NI����>������ ҥkJ+�	�:l4zh���V
��-P	g�̐��}�&''���X��R`��t�>����&=<��rޱZ0���~�/��^E#0���c���ɪ8օT�cĬ������z��/�z�� b)�q:�N�g���!󒕺!����
�R����r����O%blا;`Er��cj3Bv�]�=�]^�g�ޡ���hLU�	_�R7��0M�q>"�H(/�A{p2��H�I}"��ߟ��� ��)�����Q��Mږ��g�1�����۫���
�麐��[=��5��M���M4�Z�d�Ǩ]p�9O � Pi����v/e�̂����/^~������qmk[�D3��ݾ����Y5kmeA��b�v�!��+��c����r_�(�,t@�%�O�-L��޷���<a#�*w2��_N4j�]*�:�����)��z#�i[jH�Ʃ�� �]䘕5�*�T����L���� ȓ=�%K�%Ӽ�O��b�]�������3��p�)Q�8�����톛' ��ta�Q���rDVa��ł}�E�]��h�Ώ�D������Z0 @0�VZ-Aw�L�E;W�P<'&���5Z�����������% �ר�
�X{+��eK5���%��Q(��u�DY=u��гQ�h��/�𔸌�g��ԆV�vc�&��D�V�3[�J���,�ت�5yY�	�@W ��O���`
�r�]iȬ2��I�0�79��k�bz喝�����Oz�ʝ�x:��п ���1�1�Q�I���*��k 5���|_�e��VD>$���#�x��G�q�����T���C�O��A��a���x���Ld�c�b[�"��A���Ԝ��!��bnD"naz޾�o�^�>��9W�T��~ ]�����!�X�*�֢�c��]g<�C-Fs��|�[�������-�����pH�׻��zs�Z���m�}�G����N�������?,�&���z���F�}aX�
�'��h�I�Hƀ2��۲a�r�l����4+�A?�.�Vڧ@B�W��J��������l��T��w]L�n��������;u�9.����ٛ��`��%�gi��PR���σ���#H ����X<�J���U�T���3\�!V!5c��Q��ڟ� �h����^�r̢W�<U����_��nȢ1�d�%Zd��C�"�V�]��9�NE��9�S\	I�S�xF���P��d�9ʌ�W6�JB���r6G������1���|��\
E��!�{���l��Q�! 9#K�i<�ժ��K�i>;����R �(��2~:��>5ubB��z�d�<�D�(�<����;�����>���~Y�*_^R��~3˝��|=��?����N�)�l���|��$e]��mY�Q��#��c�=��ì���~MT�ޘ�zt� ����)�љ|�������c!Rh���u#NA/Ӛ`����<�(�f}��4*�] G�l���f6�(��7-�E��X��Yv��{��`�$�i+�9�u:�5ؒ���!��H�taO.Nk��ۿ��M�d����n�)�<�g��Z��j�aP��&��ܜ�	i������On��V{�� f�>'�G�
|%�gl����I� ����1�O?��L�f�$!*$�3XÀu�I���d��35�a^����t�6�N��N�x'<�X�O.E�HY��f,9�tأ�p�t�����jH��c�ڇ�!������q�Dy��ܺ�z4��B�;����b����a�� 	9o������3]IPG���i���4BN�לn'��{`2��O�y*؆n��g�lu�WB�T���ς���+.��:x��WN$/s�w���Sz�Q� ������,A�v%��)�DZ�M�'��,������9��ٟt�Z��	q'<�j�$�p�8n� 2Z�#���J���a;��\�G�r���g=��X���Ss,��,h}�)���"�$L��la/d��E=mx1UT��
֓8���%`��x�?봕�����i���?�1�$��+���0|S���H��zaٽ�-(jXD+Gݔr)4�b��D�]��Ҫ8l�(��.A��M���õ�f:/5��G�"���·G��y+�6	���v}?͗B߼�'��ɣ���е6�&'����A��s^7��Kr#.��R�7Ѐ?�?�go3r���Z���+�x���{��E���M���o2jy�����Z��D���o �m1|���ē�ٕΪo��(��PR��<��@t�-h.30��N�ln������I�Ĵ�o!��.�B�5����bb,�����T�%��6�^T{L��)�ȫ���N\������P�j%H���d>�Y(�ֿ~�L��7���{R�Z>���̶˚��KB���U]i&�����_�qr�:��714S<��mn�=��b���sw���@����kh�]TH��7O��O��2K.�Ё��v{o?ꟕG�o��X:���I��Գ斬 5(W�}P�F�����V#F���
�[��:` W��{�fH.ցӯ݂�%mB��Q�>���'����oe_�`�(�`��	� \�~���GR��JZ�Z��g!��{���h�j+����F�S+�O��C;�����7��2�: �� [Uc�h��su'�4���Z�t3t��mt��XrO�"�.Ȁ�dZU�k�Y��I�,��=��]�Iz�����d��#��X�hŁ��gكeb�p��S�����3ޝ�JI�&���L�5I�CA��3�y��@��5�3�d�f���MQ<͂��BW�m¾Y�vz�V�H+x�%�샯g��7pj^��A\�I�P{D��)�nm&(������nGI
(�6;�e=�=e0����TnI��!�?
4��,����Z�˹�5G&�y�4]�ܧ��/��:�<���n�h6Mn�p�̫w^ .B��l���g�� ?�.`JПV�m{��çi��o�<M�V����� $}&1\��<��cmx&�h}v��;>B���tlv8Qʻ���R5�,�؞�_b}���
̄�2QO�Ch�|���	XJ⮜�}��QT:����Xg��>&��v�k����ֺ`���ѶC�oS ֽ�������e&$�\DQE~��O���Ծ{��ĞWs x��ea8D�fl��J-�=��w^��\{1�\Y��b�i�/魄�8-�1(������޵����ņh��%o���~����YW��<���%
�K�8�.f�r0�*���<��*�F�eɦo1��٧QHy��s�]��5��0�.Ju������`X�_:�@�=�u����{��ӦV���ROD��N4�Yn��ڤ�"Z絳ѤL���}^�rTF3cV�.7֯!��C��r�k�dX���$�X@P�0�a�+hoU�a!SS�]&�e>
\�Ζ=�^���ᒋ��g�ٛ�x_�|����w��䴦�n�N��;���*�j5��ß�Z�O�оn%�r��(������)X�D�"ϲ��I}�d���$9���&�p��@�}R��ѶELkE�4`��ڲ�����<m�g�j�7��m�;���?��0m����㨠�7C���t���� {U�������"�&�zbŦ:��@M��Cj�dH�q����r~���Rty�啈�8��1]��y�B��H�������s�!V{b��a�}�i�ǓX�T���[�;���g�\N�/ �]��k�L�ԫ���I-%ш�R2�k'�9,�܀����l >0z�ͯ4(���(7u����~o���f�����"D�����<���w�1K��K�vz��v�f����W��\��Y�V�����M9(`�����˟&JS�z�i�{�g(y�gW���.�A;c#h8�u�֧�a�w��ђ��5i0܏Uk*�d���v�R�����RÐ�� `��&fu
�"wg_^�e"�}�3?Μ�ȇ��1ꐏ���h�C�gT��_O� ��w/�: ���G��м�;����*��djMi o��i���)Hj7b)3�֖�G:��H<�ff�Z��k	�˛��<Lo4�=��3��W1c�����_+E; ~�l)��
���e�CR�ڊ��l�]Ql1w��<C�|t�,�B2d{�kF���9���om��h�$οuL������f$�8��4����_�V�3ԃ�^^��܄?^/�>}s��e��ɼ�����[�x�F'_���Y%�g��/����t�Z}�]ဃI�vTm
A!-?�el ��T�3a��T��gE͟�=ॗ�����G8��;!�IBA;��V�A�[�ݒ2LPJpe}��g襵�ӁW���=w;�  �(d���8����p!u�����]My���ti�V	+��Dm Y~6bق����v�z5^P+m4���!.���B9WY�0k�Y>���aǹ5)~�XX@˖t�nz�5�N$},�5۟�W�Nk�6<�{3;�90�~�_\�wq߹��5+�����Z�"Qybw]�w��Sx:��3]4b����9�m�W�S ]�>M;L�?��.D���ޡ\�������?L���蟽
�b9�ܹ|�Yuu���#�
�� �G�()$�Yw�M@:5[s���+��A�뢇��Df]X��?J5��gD�`�X�7���tL��	<PN+>#Y=^��\���px���k`q��㱇�ƃ�2��|ÞSҶ��7����D�
f���0��p��?�Ң������67ݢ������hWA2�@�Is�-l��I��WXm�+��¥_xc8�֐=�'� �\p�$��<�ǐ���+.��g�i6y�h��݋_ǀ�^\�;����"����47Q$G�?�M!��⽵��iB��!��S��C��|�˙�P�쨂8�9S�O�<�@KE��YZ�g~p2��N/����L�2MGU:@)�Y�Sq�8Ω�0�p��_4���˝\y9��Ċ?��y�\�BSE� 0�膁��i-A����C��B�"MDw��D9��8���e.���xk� ��Iꑃ&+�E���W�����ׯ5��#1�w����2��X��2���M�CGA��k&*/���[4c�l�8�·�|ݔ�Y������sd)�
�Mj0"^��99��]`9��h���w�|�k֙��@���/�31/��!Q
Ok	I�pA��t��	ǈRF0;�׷5�w�4O������*]_ ��F�2��IG�?b_A
���,�*i���&�V����,ͱ �+^�RȎ	��up2[��Uț1`QI6�O��z��,%��mu���a^�j:ũp��ps6n�% ��J���=�Z<��JEE<�a3΀�v�:�i`=��P�ۏ��3���[��Q��S��c���;/�i�ܶv|@�T� ;P��;���Ξs�c9���t�+�۽F`O�>��=�,�;�����E�$�Ml��38���x�o�ؕ��?|�eEvm�v��T
)��/dJ^G3�%>0X�3m7 ���o)�A�o;P4��q����%�m��'Y�V(�Oo�C�:"���,�ȉ��̤b�ҧ�wث�C9��dG�1Fd�w��T���=8��"����ܳ���%��,A`�z�~��&_�Nk�u�w�V@�5p��t�k9Y?�px�kR	� �-��C�z�-@��/�
g����� )���֋��\�D���>~P�L+�6���6
��=��R�����<�6J�)����|����iޭm[(UwVN#�%@9iy��W]k�"N)��(}G�����2��}{���\)B�ME��X���nN�BҞc�>���9;�xΠ����1������I��B���K���Z��h��N?��'������,�+��+ܓ!�q��x(eC9lz�}cp��P�����~GQ	��-ȩp��'�$]HI����{z�L�Y�NV�f�}�����-�)��=��:�6�����<�v�?TL7z*?/\�7�2�g��Yu㴪K�O;�E� ��N��p��;�ߊ�<y�����`xՅ�I����f�P�3t�>�t�׃�v`�6t��n_Ri�!��MQP�i @�W:�o*�	�̗��(ic�m�>}&:���cM3愉����Eu3�(L8�3 �>�@E<��Kef��V0��H�� �;�gϣ��Ѵ��Fz�w��/�N�Y*bR���t�ru��nǴF�m&!�4i�h��y��Y�\�J�P����0Og\��1�,�<����%�����.+�ef�0�N��stszM�O�gW���w���&B��ɣ��un�#��"8-j��+C΍7g�ӂ�
w�sg�f(}� n�0�f�닸�F��	+��U1qq�߱��@�E�Ȋ}[�ʡ��)�~$xp�!��n��&�ז�gj��'�t���Q�mg�%z���g�F��w%^Ӯ��59.L� �  �6��-��I���1�S2e�_��G~	�PR~�b\����x�<�Ʋ���\�
�T@��m��k���N��m��0EU������/ w�(X�~�(�cr�*+ݲ