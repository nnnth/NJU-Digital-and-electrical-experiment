��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��rs. ��t$�x�P�~��� ��gϢ~�Z�n'�S��j�C:E��U,�o����(]�q���ɠb��FT3Kf>�b��p�2s���P8`#3�L���*ـC�0j�����lf#���P�RG�6,��-i:"|�y��F�u��y��j��#��\��]����Xx'���fT�g��V��l�e$�j<�B�ʛ�hF��Ϗ����Dt����׀nc�.��Q����#D��L3��1T���3i
�,Uv��2�l	�7Xxy��.�,�����0�'�'V	�{�]�5��ċU����>t�3�,Ly*��h��pZ��&j�6��~�{Ov��O��:��n��V¶���1���B`o���DO敫W"�|�t�L�*���:��l���x<����K�����ꉐ�����i�$G�hw�Z���	���yfx�\��mA���M�y���)���%�
�2���cA�:��<���N*럃ҥl�5����;�=�Pw6�9��ԩ�?��l�P�J�	Ѡ��;�V��Y�>���v��i����vj;� ��Zj�m����G(J�O������=6�~��D��3�pU��B��v������ 0�D��^<R u	�&�� �I/�p
�Ȱ���+��9���HA�㙀D�4:�Tj��k��>x������;�c���" �̰�5B�h�I�[��gf��C�v��s¢ě:��> �W�Z�V7b�Lpe�æi�b�vI��C�[�Q1��h���Ѕ�@/(�h��lXd 0o��mѹˡm�NP�v��ާ]M�Z������pHCPQ�%��kcX�$�ȟ��z|HRp�gU��꧵�v����l����z�TGX��:���brU�D���z����6�#��ҽNx��]q��MDP'^5D ]RO��>	�K�+�LG�%{)㉁}C�xnK8�⯶O���6� �����oܔ]��r��nWs�|�.V�_
D��pW�ݺ����A�=7�r������&� ���D_�N���2eܛ��wR�KY��z@'��{o���z]���y"]M�e��FD�h�$���}w�5-��^y}�Q��M=֡`�ꋧ����㏖��� ��h�E��&�j������N��zϚ�6�]��
z0����	>�3-���l���39w�~g��&���PI��l�K���l=6�)�����|��h�