��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��X[&-����v|��y���]H�lMI�C����e����J^�E�e�_a� ���g]4�n��Rz���	d���~ �@�����Ã��m0�X� '��O��ef��y,���r����q�I�l,7� H�/I��J��	�o���Ŭ1�;��"��� #:/ߟ�+>ˠ`��� b]�����O	s��"}�#;@�iXG�
g�0��x�%����zZf���ݣ�'�3��>?��F�_�ʹ2�O�]3��ED]4��t��q���{T�)p1����*f��7��P>XS>eC��e"b|��K��>�fBz_���RU�U��S��*�?ۚ�IH,��mp��+����z��ו-�@O��e��Y�[;���Sz���/����GY���$	yK�Q=C^g���c�'U���Ł��]cKJ<v����^p�"š�,VK�8g#&I@�4ёg�O�8�G*��u����mܿ�*v�t����O�ѓJR_XZJV�b�q�u�Qe �;���� �C���o��s�h�%�C��#��x9��u�C>��u&�tݘ~/GN(:=iy�d�(���%�X+�ñVfn�������a�@2�+:k��7Qu�Rݔ��
�d��R�i�����W�MZ�6b�I�%�������׌WrK��Fj]�p8�z�r	��MJ��매��x"밆vw�}��|d$�ua}j��9a�N�o��_��ԏ"ߐ-Z�c����70+)
��G�ӧA
?���+x5һ�l�t!�B"�2�WG����X�aAܣS�gɽϋ���h��ENT�<r�p��Z����M�9�9��_S�l�F��k���؊���$<N�L�վ)^�0�_�����fL�"dZ�cO���߷����/�FD5>��d0���9��I:F��zH'<_�'�X��H
+������x�����p9��5E�i�"���X�fE�L�R
kA�6r�d���sZ�Y�,7��K"�����F�A5�<��Hǟ8�C�@�n�@��ٜU��+O���p�~���9�?i� �9�aB����rrx\�~1�����/�XD��S�C	��XQ���2b�����*q��}��u���:�\8G�Ѐ"ݲ5,��j�O	�jLp��>[o#��P2�5�\*
�������ࠁIF���ߨB6�{����M�M��x�QX$�L"7ցc5�-=�k9��Z/e�;դ!��͇�&�v�}��ʁtGZ�ܱl��(v)��� �6H�2���J���6F����2b���į9,���W+C����Q\�a��1��'��:��zo��p�Xʁ6hFG2�E�d\�M���#�ˉv����v��ꞟ΀Ԃ`o�3�f�	n.�K�������=��c���[���y�l'�A*�;Yg���w���g��n
_�Q˚�������H��E�����|��˟���M̬>���&dXg�L{~`GIk��cߙ���Xd9����ܰ��]��[|՛m�_~X�Alf�z��&&J$c6���ɴ� N3��^--��q��8i�@��nW�K`��t�wx�yX�;Po���	�lk�>0)W:
0V5�p�}9f��9�jwdj� �Y4��?1۱$�x��aT�\y��!��.�|�wޖ�[�v���6�u�apf��p2=J���u�Hcc�������^�{¥NrX����j�`�/�q��B(k9�F�s-�����Q�Y}�2e;J�A����P�gi�7���9�x������SY��J7Vϥˊf��3v��:���d֔yO��^�;���><'5��-��2+�dS
�5�]ǥ�
���RX�R�ܽӣP��Ā�2]b-G4#