��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�ٿ�հHm��+���-�eG�7��	�b��O?�]	�����m���->�����D����̅������oT3Q7���u��F���Ot��MZ'X)�f������^牕Ǿw�)�:,N^c*�y�?�ɛ�qY~��藇nd�~�H�W&܃
�/�i]�r�	,��oQ����n�����<�?���&�0A�}���Gpj>���X��bc?��2��8��	A������Q�V�|�(
���\��p�~�����3ٲ|om���ԑ^{d�#�\]��X(p��]3�'[ �ӋfZ���*�[FB��}((���}�e����&�m������(v��9�����g�/[���Z
�1�b\�&��9����MZʥc�ư58�FO��'-���:�HP9�pv��>h�hG���yCh��`�I0,C�����xfi���=Q e�/����\'f�O0��U�'�j�$���=T�p{K��e�m�=�$]�oE͘�F�_��wܠ��ݴ��7�tqd��޻/3��2&�L��S�(Yִk���6o�sR0�����:ߦԭ��Q+���%�Mix{� W�vlՓ��𹥄�����9�+44?|�>#\	a8�G�xP��w�#���<f��4  ��j�F�$-�� ~�����������u���)�=�z�}o7��F��� j������BL���W��wT�>������̒�UxV(/� �Ő��՛�d�!#ڐ>��g��d�=/��n���Cn�z���.�^�R�����әِ���<�FU�m���J��j�@)����,�4g����x[km��D�)A����+�'��~6������.&ʷ�mQ�w,��2����sz��Ik�Ԫ��M�lg��w	N���6�5�eV�I�g4����kS���#�����Y��z�!�S�����jpsI�?i�OhD���w����rMe9��GA�5�u���ھɼJ��+\��ch�6��[ݡ�uu˼���Y����7|+�J�L2�;��Z@H�+�͍��GԹRnE��:�*���\���O]�M��Ej7SQ� ���~@͏������1nK��e����x��7(�2�pr7���>�L����6�o�(V�*�#���k��w/��j<�[�_Q_6���c]}��sg�=�J_���P�<��8�Fv��N}���P����CR�7ʧl�#i���v�NF�!da�ߎ�.X?�F_�7fH��=�#��{.�jm�����\L=��'.=���J�)Í���*���k�M���n�|�V"��/٫I��mS�;U��]'��-��j��-U�:\Jv�g�򼎝��T��L��^D=�A6�7T �>E���\���J���'����������yw#�Nkw��������ఽ������D5�r�\N�Ǝ&g��������P�I�T�k�o����Q��75�ҹ�Β_N'+��&[��`r�#Lv���l.�f�v��6XN��N�Sg���-��i��|��za��;��Kwz^L���Եl���WJm���G��,��5��2�@�p�+��S��	<)~�]._�e�����	-u=�[NP� k����Y-��G�ī`��G���@F�z�M�	������ԯ��i�ݪ�B�1�6�n��*�۬1�`[�����Ri� �G>���m���K|���΂��g���w���Y���"�|�����=��e�/��µ�CJͨ�f�s���l�����Q$��X*ɭ�2�T|��b�4=v39��1�������(*��E',EDg���\;#�1J3�	��]ah�V�ɹ��B�3��vB��~2#���@�O�E��1���^z;��1P��t��H�y�eS_�Y�4ܷ�!��$H|[����r���#�:���[���e~��������2%�p�#�l7o"�k���hH���(���U�(�f�m씘�0a�#�4�q�t�.���9��H�o����U�Ŗ�2�yК��K@�u�KP�m�Z����}I��8A��}��t�
K���Ldb�ݐ&�yr�=�����i�7�%�կu�"|fv�F�����y�(Mi$x�S���Ę���+�T�|����u0�)���\� �TU�@%�������\q�X)��QINge���u=��ϛhm��z�$du�D��������g&ٽ0
J�� 8p� 6�m�tc�� ��
.dV�9���CGsCf�7W�U�|ӄa�D{��ߠK��C���m�H�`S�=S �VU7y�Y!�t�ޘ�� �^f�]ĝ���#@17ڹ���р���P;b����VF&xd]��x;��+�0;����ȞT*�,QJ��Ї*s��^ R��Y4�q��M�D5���\,a{�q���Jk{�*4x�g"�Z9��b^���qNc��2�h[NM��\~�W��W�<YY�	
�K��X%���Df��WҺ�����H2�t��������¦i̓��.�8LR�Ag?�nm�m���_���{�^�j�a؜G[p��V�
��0o(PYv0��Ǔc�A��=��Q�ĥ�Az��`hi8�>���H՝� ���Z�n<=�>� �`��;?�>��J����7O�%�~<�^2�����Z9�^��1McT���틢��B,�&B�Pd0����x�T��;oQ	�v�:%E*��E�MyՕU�E9m}o�v��>4�H�Gz@��9�F�LV4�_�[X���0&F
ׅ��"�!�T5U�)��oe�N�! 44,3�8$.�1��<�H�\%'K������R\LԳ�Q��g��ۭS���Lp�mI8i9*@��Z'i�B�s����lF�(���bK7ۦbt��D�Lҁ0`B>#3����ڛ��TU_(b�f�OH�zp�������M�ދ�6}4�єi�!ª0#hoiȵ�(庅IHX������
[˒�sz��z:��>�i�Y�_')��S�O���]'�?Gfѵ�HQv��y&�*s� -���B���D���L��ڡb_GI��e:���-���vڣ=��)j�-���CD��僇�t��@*,"1z����Po�B�7O�'Y<��娆�E(J��tD]�C'���[�Mh+PP�qY���O��󲿙Y=� ��5(�;��7��Q�ͽ �-�ԡ���a����K9�Bl�3M=0�h,��6'��[A�&��Lf�~�iQ=L���!]KVv�Uҷ��I���������(V8����z�3J�"��M�*�5*ђ�l���HB�O*�%����$�"�[��Kch��OC�~sB�N�_�-LJ���)��<� v�=�{�<$���D<Y���(Q���U2�>C�{��9-��	�4�R��_^.�o�Ѓ��#9.�t�Q�KOz�/t�\��GV�=�]����M����Th�t� ��s�a4+�}��x�$�J{`����D�.�属{@��~d@�	һ�^XK0�tzl.��y�:z�!xp�7НS����&�s���g���h�H�8�r��0d�v��U��ҽi��������;pU[��J�%bT�������q���Kp_b֥*��xV�����C{v�ê�J�
C�'E����v�(�mO��'��*dp�v�퍊�E"A�>3�桤a|��=�&��
���
Ԍ��9�&� ɑ�l�3�%!���W%C�L��?Eŗ�����D~���u�|��������U?��]#����A6����s�S�D���)�j@�&⁯��D�3��C��W	9[��Z�sq�<
���"Y��~�'q3v��
�'uǑ��\�"��߉��?%�/ :�:O�t ��A�ǯE�_K�@H?P��W_�wٻ6s�o3�_�J�[v�6�/;�Ce��"B����($��D@#��8[�x<`ffG��p�I4��a����YC�]��!f��d]^+������������Kq3����|�7�#���8��00x��=���u��I����vٸ_|�r�� R���=��������������@���kF\�k�v������8�O=��A��r�J[�D�
�,<l���W׌}�r����z���B5���Vӌ/�4��G<(1�m���n��к�3��ҫ|����od2��� ���H�=<򺔇��A�U��l�.�{�"�x[��R�\��i����Q�R����N��w����E;��J��6�Aay�B �p���������/�� �W�n�6��A���c�ߧ�bW��c�M;�o���	\��d�aX��}��t��ud�#����i����Y�5�OڿUl��TL}c����lєRH㈗�N�p'`nvs4v���H�Ŵ�Жx���r}��'�BL��6RLX`�M�B��̊�������9=c�!Ե&��7�ck�.q6|�i	�����Ǒ�l%d���q} ����g�jZI�_d����OP&�=�L5�0e�ˆz�c���a<�Y��!�`so�6�0w�-�5/fs�N����Y5�6���=����%2 1)�\>T"v�6i�2��!xJb�-�16T�廇@��5�"; �G͖܍D�&��'I(��3X#�#A^.�\�ݐP!g6��]Ѳd���OY.2��dn�nx��7Y7!tR^$�iV���q΅IíG�lgC6OJ#�&j��#����2�� 2x+��	�Y�S�~Tt4�u썠�&��@���Ʀ�Zɶe)t�k��-���h
:3�2g�|];�^Hx����-���c�`g9�d��l\�X�^!&�O.&&�F��c���9\B��)��Y�,9�Y������;����z�K� X.��ޭ^��^e���&.���g$dL�|����T��]��x�a$�l�aK����P��ȑ��R��5�t��f��(c1Da�j�s^v�@��%��j�W�yˑܤ�8��\^�^X���Q$�js?Y�h�ƈ�G:�p�P;\���#��M�/�$x������֊y��uM�&��0�|x�U��o�#|��3�TS�
�$��Em��]�=A�Tq��Ӄ$G�i]$�:��$���§�n����]`0Θ?�a��Dw/Ou�����a���ds�ir���B۞L6Ͳft��>�P��	1o�>��M䶙��"��=���7�9�נ��d�3\�U�I��j呣5����3��J���Z���_�Q-V���#�P8�D�"|���Q�0�����<��.&֧~,�珊�Mv}�ܠk�TI�w=	I����ǁM��q.伽�fX�3ΧW��(�(b/DG�+@A�6�l��A���4!��]^di�����fV%�x�"W*���D���n�(�E�.������eB�=�Qh�#A$q�9x�;�丯y������ϓ��u��Z�Y�&�轿������2hl;X�J]�͈<M�Y��j1A�/��~� o�w3�C����l�z��(2�R��df�;2��Ӧ�'S[�P66���� �=(1Gx�*��F��?7�E2$���n5����fH�h ]�^Z&e#?�N�E���<R+�dP�[�!�Vu�� ���1�ȷà�+��u~�RAm�=�=ʅ���z�_-W�APs�'�V;�~����Z�FN��]8�}V;Q� ;,d:�-K�Y�
2���7�D���:��Ruq�k���njӈv!ζ��MKCO5ֱ@���`i����Mi���p�q^��=�6�AaBt�}9�m�^�7Vʳ���M<��wy?E�bH��������a�A��4MI�����s�]C#�j�>��R�[z3宧m�lf{.�b#����<n*�k?�;=���������z�~�XpYʂ½D���(��`#l���ŭ�7����2�{����=s\�]��|���-��ac��P���E"��������>N���]�J��xKϤ��h;Bji�x�,�~��?����
�?�/�TU��,Ff���.'����I8���$�nb�j*܀膸Ug�w�~׋z��,W�d���tS�u��t�l
k�ܢ�x�c���,������
$ou�|O��@(��D-��Q.��#�m�v{j���d�N��I�Ӗ"�1�/��y�� �L��)�!�Rrh���-c���WNH}��"��"�r	��=;�N�P��Ya �1?jQ:`3\W����>�$� ^�mV7�r���ʏ��3%I����۹K�g{�:�[���쏉L$=�x� ��ڋ�s!U�k�E��G�糡Vq�/��Si[M'T2�j��R��L�(��#�;}J<ռm������p��Q^x����`��]�##� ���js� ���T�(Q����8���9b��fw�OV�i�E*�A�SI�IQ��Z����N�O&�"[y�An>��9+��\��W��D1)�ZN���5;�<��h�i�"�E��8cs��fL������r��JiO�&�q��"j��k"ʫ�$��e��N��dб#�}���/�Q*�mfK<e:�4/��t����tKE5ވݽ�!��d���;
�b�����:�Jղ�9�]�x�E0%<��e��T��k�#<zțvCH��)���}�+H{��ɜwc���!�fJ�F�E$�����7�RS'N�=��5�[��oj���}� �O(��Q�r_?���1��dɻ��xo����sWʸ�N�кx�ʵ��K�ys�O]������w�5V!à�1^�9����`�"y ���^ٲ�'�O����2�1x�N�,�p)��%��K%��'S��c J~�D�4�^���v(j�Q}j�ѴsJp��GR��T�9��&���	���c��R��^������-�����j�D����������P��#3}ߧ�_����u`D�� �BA'��FVVUȡO����6��-A��-��KEA�{�V瞭L9^7�"Lڬg���CyUP�w.f�LO35��{q�=��()�Dx-
��=�X<e�afe����6�����K�a]���ǧ���P2]X+����:�H�kH)��}��^� CwJ�v����t�u'�.�Q�ϩ�oh�F(qmd�8^�M�nT��g]��ĆȻ�,�I�]��&�y4�� ���np@z�;�̒�I�ϗ���,&!dn5x�$���s�pH�U���ٿ�-U=�=�!���8$g�Iy���G�����T(��OW�i�'��5��6n2:��܏W��?�N��6�~i�����S�Y�����lNk�T���	�(x�	�����G��������J�k�� >��֙IM|?�|ߥ[