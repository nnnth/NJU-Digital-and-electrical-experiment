��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`����8
�2��'��C�%�@��.��ϲO���t@��n~�O���:j���t��4���NݑBU�XC34����EKߔ:�i��.&F��䚚 lM=� ��R�<������#�O��Y%�O��|K/.?{���b[�O^}`)��Փ�]xpn�PB%Sܪ$;Ut_�E-#E�s&
9��7���I����k�%z���I�t�f�KF���������f��"�I �ߔ��"y�~��`W�d\U�2똛���w�蹏���
��+�88+3���L��B��Qr����4_j#�����"�����eW�E��<�7�U˒�kL�X�ּ>���\�lJL�>�~"�
ޞI�E�5�,��5�0��H�x/��O���֫�w�0�d��n���Q�X	Ey�P�Wt�R6	y�$��g�^�u����ȶ�Q0_�����@{�E85�!z�]�o�D)p�:,o���HY!٩I�f����	5���ic��K2��y�Vċ=���P��̕�>GI���far��+�k�t��\���⇉��]!`T��v"K���!c2C�ܹ35�O���%��@���W �����O����NK�.~��;�ԟf�+^��J��,�{�<�A�(�5 tJp��v+�/Z�M7 ��RcE��Xl�(R�b4pr�a�u!���V�Ƣ=���^j��Fy�zT�ԉ}�?4ϫm6({zΣ�D��5�x1��h�e%�G�Rң��G�� ����y8��f����AƹT�?
��������c {ěb)k�r�Zh��>�SǄ���:�`��W!�!��;��� ��i�;y{�k��=�0@&�f�#%-~Z��&4�pE4l?H��!] �N%��	������:�U��9�/�&��*��49�J��#I��5?,��O���[P#0�)�N��ضoE�
E^��[�����5r��h��o=��7�hr�/�W��aP1�)��%i\���R+��2��in3~1[�,.����c%˴�0�(wZ��*9�y������(�{�q�����-���6ߎĽ������d�x�k�*fr)R��0���1_'�~�ؔw;h$�=��E��R�%��T���A�.	v
�	<Ϟ��WV�С'�a��R�;:"_��:��~��L1g�- )�%%4n�j�_���)�}# �\ǖ��"�y=�����^���C��+����?�T�;bӣ��qЮ����Ga�2x�����7-L��%� �|��z��@������kcj�8>�8��:�1~K��`��yQ�������b}�+�`��F��YW�Fr�_-P}�H��ڈ2N9*��$��\'���?�����?L��ڥ��[�6"��<A�P���W@�l��J_���"�j��H�B;�	�l�<���Z�y��k��qzֱ��@Ղ��?���!-�yY#\�\܏衭�/-��Tw��+�?���7�	Ҵ٦.gs�m�~�[��f�+��C���G,~!��kD�2$A�����@���A�$!�|��^TJ��fn�e'&-S�M����^�=�$��C���D,	<��������Q�.`A'5=z���E�>��Jl#}���S�Ea/Td��]N���F�J|odg���毑�z	,���6�k��^\ġ�25�#w+��/�]�C�q	:B#L�rmyX�Ń�	���cm�)�Yf�"��«�D�z#0���~�g>\��n�4�e�s����{�`�9N�� �8�����I"D���(��o�7�*���_�n��D�(�6$Y@�v�2�߶��5��,<�?}tv&��I!��]8Y��g�n�C�ؚ�.'��Q����������-$�j1�ۚ'
7*��N'y�Ş5���2sQ������z软�|�z;0�ɰ�����w�>P��LȋY��-�z������p���J�?�U�[�͞ќ�,sl����QC�J�q�<.�[��-��ۦ����t�!=_
�+���#�t����j9�A�Oy�V=W���h3!�*N��&�S��v�Ư>�[-���!|�jb��������)x/��X\� �׮�'$udI��пP_ԩ�;�u���R�N���P5��GJ�]zl�/}Tm�ݯN��g3��X��UI��'�[�Ts��X�d�����U���� �w7	B���3�%���?5�l��81�6�}kHH��=�{FS��w��)!����^K��-õ*�.�d�XnR�z[,G���Z�bu��He�5�_��P�z8{z ゗���t������Z.�z�D"�H���!A LYp<$2+�򍄉䓐dl�m)�T,�l ��=%�L�1���f6J��.���Sf���Iaj�8��q;+�姎+��!�eY���>��^hC+�.�枦���sp������:���odZV�N�s٣1 �
�#�0b�i��N�z���wY���E��2=�E]�����(d\�?�2�J� 洤kAM��5BY���'Ěv�b�i�6�l�c8�C��t�^����;6u�!����1}�Z]����̦����i����ߊa�K�OQ�(�4����^�2R�4��Jжg�_���uA�Y�B��`������RM�R�ݰA܁84�q��1�4&{DZ^�9�@�~ٹ�a����מ1N]%���t��C4N����z��ʱ�N��g�����|�!�^)��A���E�|ы
��%X������?��"0or�U����#ʋ@^W�����m������ؖ��H�5^��i2DB1I]](�%����lq���z��Ƙ甆��5N�ĺ���Z�Yz��L��5g0V���Ck�� ������-�=q�5"�.��зۼb��F�7D�4�y�Cހ2���Jd�s6R5,O�lR~�з�I�f�NӅ*>��)WNE߃��3^��|�s��t7���^Xj(�SW��x���7��7î���*X�n�>��l_?#Q�w��RGWa��p���� ���ݨ΁��X�f�M�(&��2���AZ=ꔁ,y�r��
�Eiˬ�{b��e�eͶȘ�%���]z�������:�f��r���A/�u�#0��7�(.P��@u	ފ@cڅKIچ�z��\��^����u�t,���[��#�n���,��;�Dj��l��vf�誌M_�\��ii�N=@1��w&�hx��ʑ.��ҵ�+&1���[��u�E��}fN2.����#�i5Z5�+j��6�<��/��O�E(�jf����v�]뻋3�_�_ըQR��A�!�o&�k��}Z��zu��t
T\�k};�0����ȩ�vI���	��&qq^}������:�f2������gjH���Y"Ío��}:�P�¡�r�
-Ҵ�KQՃsl5h�跮;ў/��/"�j�ކЏ�|c#�A򣎱w�o�x�IOe�uuy��4��ǽVd����H-L�Aޕ�/�t2����)Qf�{A�6���Ԉ�~���Xu�ZJ����C3�� �VLds�B�lD�����8>�8���������և�~VZ�k�\C��eÑ��l�B+kʦ��{[��i��[��j{rs���b7ƾ�:��{���ȍ�cz�a�(���$!Rɱ&�<�R6R�pa���'/]�'F@��RsH�t������$M��+Na ����.vb[�Q�}m�#S�#���x�TuӅB�G�e���	}��������;,�Rȕ�{_�%1�����|Gbd9 w�1�����s��㢞�s�+w-�Ti��L�yW�ߠ�g��R�Nk������y+���Q3:���M���afR��bq�$o�]V͈���-뎠b��즑C��y� 3q0��u�)t�du�E�Z��r!�mY���.^�烙)��E������p�7<����>���_��GܨY�)��{���ET�S�/�t��y���T�-��O��Qad��d����a�B�k�W>��
�X8@�I� tdQY��Y���{�����F��!�j��u�ȥ(���Wk���-�����e�:�-:��͔�k;��ł��X��`��F�Ǒ&$��,��
D	D�S�sAr�o�0��"]����ć͕W�t�|\\�O�����Fo��L��~�ٰh��p��&��7�KjCT���Y�Y�ṙ��N�_]�&KKŪ�qz��`^X� U���en]��q�ag�jI㶍�����^Jc�驡#�V�
�� �*l������cB�M$�e��J3��G�p��s�Vi�%,^h�;eӷp��dW�VI�(ň���>b`��}Rn�j���	������r���8u��w�¬y����t�b�y�]�a��m�#���ds/%ډ�Ms��a�^�q�������5���I//�۲�M3W�����덹FM�����$X�O�>�)�������~�!��y�)��i��A:n�z�Q,���æ�2X' ~$��s�M54��	(��bN�w9<�GHǨ녣u�c�N{�Tw�C�]�E�����"z5�:mdB�a\��?��pD�����wZ�Oz,��̼�Th}�_ج�� �������#A�(R3Q����Q�mj<$j2)�(�@��V������C��9��S�D:γ���NM�T�q8� NP̮���)�:�|ZL�+To�&���n��;�O�!�h��'�x�pׂ"�R�v�bie��.ֺ~4b����:���ˮ��Jm,�� F�-����#[����,v+jd����>�.m���zYL� �jr��oƄ�'u��.-J{���W�F�Us 4�n4�Y6X7|c�O>��6�=r7:�6}ޝ4H�	�3���v�9'���N ��9,�����}(~.��	+���#�oyh�~}�u��7HO_Q��0�)@������M�/Y�؞��{��ك�i�.��ri��l�"\w�6� �D�u8��8�X�-���cF]h"�m�a�n��*��R;h�,� �(2whS�q������xۖ&D`K�Q�2	��[4�l'ҥ�+	v��`����%6���kGWo������%�c���-��pA)�~��Qќ� �*�38zL����dȰ�$��Siཽ5��WTճP��vL\�} 6��9��Q�kҹ��d�:����D�e4�S��7����7����9�O����`f�xpo%�*�iO��o͘�ŵ�~��>��x���%tNZyB��N��v+����L��ҁ�B#5�ݺ3h��G��5�=RtT�®-�Gu���{�W´�p�"���ܘ	�6����w�
�%~c*S�pMPqu�sDM8F����	��j�4��!�1rev��,/��9/=���'(6��3t�������lK���h���w�61�R;= \5>�p?���x~�l��8�y8�T�_�^$�s�d^�d��H��d�0ҥv�$EЯ�Zp�G�1�I�pZ�|U�}�A�@�8���*�6��*:G��(b
`h��mEm���}�k�S�*�e"���S�0u����g�Db�ҋ+Ha\0&:�a��0G
U{�4ut��$����++0C ��b����CȚ��en��W�w	v���w��3�JD������%�� M�[y�LZ&��k���R�mו	n|��Y.����z�S�5!7V����c,^��Iz��_�!�j߬.��~n�.)Y�v�I��>�LUVk��M���"_��`_m1N�q)��+2xe����_�hr��h��J�<�kOjtJ�5�}d�[#" !oX��[��B������>�D���W޾f�C���H�rFz�%� ������Q ӭ_�Xȵ�0�[C�!ד	dH�^��WA$�|���&�7�� ��K�ɤk)�h,:��G�P�{FJ����n�Y�|ۻ�_��6a��߮w��Q��I��扇xb�S���Vp��^����q_>�2�g�.:ٚ �*#'=��,��X�ɭ�el@'tN��`�\>�5D�_��� ܾ�)C#��B�+L��7�"=�E��l��G�����Q8W]����yAͽ~&�xopl}��y�[���o'~�ʃ���+�C��ٸ�m�7�;�D��{a�Ãg֎%��x�=�2�#�p��H�)��)����f3�����J�8���4+Y%^Y���-rn�����3A�P�0�݈S������4]�����4�c����vh��I�;��Bc��WX��}n�������sع��vZ�2OŌ�h.���N��'(,�9^2u��X�5��P�N��0��kj�8u�)�h�Is�[=����N�Mu�	��	i��Ec1�a/ڽ��¼�~W�!1�(�ϓ�M[dkf��`��Zm(\��9<������.�������9qs�r�r	Qsc���nr8���sOg��1�!���k:M���)9�Ԛ��'���e%��w�Rc�M��2��ψ�O?z-<g]��u1$����>N�eT"�8�q4�z5e�1�ݤ2�VL$-hI���t��x��d�8��s0�!ٞ��CAԞ����b����3v��2��j�U]�B7B��
�O�Ե��P8zCJN���0��ޘ<+����H���Q S�qa����< �Ma�R|����ϯ t;���U<-�O0 �h2Z`��X2���`N�v乖͎��u�Z�zlv�@I%�R�̖���-���G���/$�m�C�ʕQm���-��!N��{G��w�|E�PJ�%�(
�Z����J�5�ʯ�?J���O� K|!*���/���]%���B�T�%M�˿���7�
zv ����
�&�C�����6{�X�,A݃�7Ь�u�(���`r��[i}�s��&�Ns��A��5Z�2X�)gN���N��_p4��1�jyc����%f��u�2A��K�_�]XV۫��6R�G�?|fл�WQa�/GG2�4ze6�7OD���t��@��M�K��E� e��%L�.A�nn���$ u��.>�k*F���ɯU�Yh�Ex��",k ��5�K}��h	pN~�a����kST��W3xB⻝��K���ga�����s����o�u�!���Jඏ�����$sč��֌]�
S:2���[m��m0V%d��HŜB������?�� �S*�2I��*��9�%pG*���/;༘7691���u�=�G���2(z��`��vD�� 46)d�e�@:j�������5�0�u�����u��}�Ȱ�!]��ޠ���`�qW��ɽd�e��@��$��v�<��Ykp�b��Bp��@q:YK�r��2�4y�-H"�d�n�ġ���h1�����L�����������N�̄�j|���>oň��l�(�M���]n`ǝ�8�܋�e�Gu"n�wnU��/�H�^W��~x��M�>@&�7a�n��2��W��}%���=��*�ݸh �9j��s��g�)�~�t���-�1��hu7�E�����aE$lB�������&�c c��$E 7�4�W���A��K$��緔\��	�kҦ�KbdS��I_ד�����RIA����1��3��z�"�f�_�l'�	�*覲.��>�H���Y�Dq*�t%{!�8�2�A2�BOY�r8V=)߿�ٮh��q�kI����N��m�od]�wBi�H��t�H�|����m��S��$%�;XdlOQ�Z��� k�v�6�&"X�=/�5�ۉM�0�ǎ�~��C���Y��6��`N�9#?3S�O�T{���2���<��8m��f0-U��=Xl�J�?+����p�Yє�ݣ�%�c��yI2� ������d�?�4&�M7ȇ�x�y<{G���ʵ�o`Iu�-���>��AF6��ÿ7DyU�W�w5�!u2}#��PL���ҝ���{|���(&WΚ�u��������v�b�$� �4�k鋻,FIL����(ڋ�_"�~_,�q>pP�?��\�T@�_�Ҧj�ۜ� �� �3��Szk�<��l�����YK()����������6̺�-�Z)�����Cjq�葉���Xޝ�3�Ru����L��Pa!�A�{�-竩��[�K2��RO�@@�%0��v�x���2�����?�'1���i��dr���R��?k���4�j"�Q�(`�\<�,d�=����뽢�"�$$� ��xX%զp�Muh=T1f�������8��4R��n�Q�6��E�x��in�"~�s��\�Bɏ�D�!e�)g����:c|I͚��e�t�0�c�`o���|T�R��'�63�^���5
҉=�;�k�OJ�C��/�Da�?���h;��My �5Sp��6~�֊�)��a�J��P�nbu.JF�]ڮ��.��xd�f�z�E_۹�6E¨��[Qpϯ���v"����!ǧU�@�5t��j�%H��C]���dX�
w�}w�@Wң�(_},߅�zX^��|X Z��Q�j��^��F����TI�L~+���]t�H�V�, o��^"Բ�3Fr�ވ��.<�o��2;�����%�c���Ğ1$R�^�|Rkvr��A�� ��͹,���ͺ��g�ny[�!�L]��p�Q}>,m�.��o	�9`E�l����bR��M[����rw���� 'q����o�sN������ �{^����v����i���g�W92�!Y���Ą����,;�tf~{t��P�
C�J���cnCF���d� �����0,pm�1;8PRi�Ycqg�:i$�R��F�6��9��\l)��bt������Xc�v�"��W��l�%�G4$���T����ܭ��Ϟ������������@MQu�ܩ�<*׶��M\���z�� t�2וX��� @%|EߊZ	��0�c(����3�_{˪�N��΢��!0�N��9��2�]kc���R	���R��t9:�ѲR���OE�V3�H��I#�2�OB᛿�5Uo��<-ï��P�N�nJsfb=b�֡��l��Ȱ1�a�SI��DV 'Y���S���M�#���i��gQ�<Qs�W�A	�X��� <��
�u���� ]�����Ȥ�.��.�������
U>
�J-�ɧ��~�~ʥs!�Q�`��݄o���6�܊%�p�:���ƞ� [U��y�Q�ǉ;�<�%���A�_�A$����!^d� ��V3�{���%�մ�4ڋ����B`�K�q��N��j*U@	�UO�<���%��$ĻG�R�QV1&���h����OW*t��dh9Y���.��S��T,=��@�[���0gڰ��I���ϩ��ͷ�^���[}��l8��R�P
g$n����k����ȊԵs:���)�|��o5���Y��5B������M��u��Q��U�yQ��O&}׭��Agf3:�h�����'��$�v��[L܁Y�6����x"(e�[�n�H�t҂�:͵t�l$k�:�u�.��${�.,�Cq�Y�"��
T��a�����Z�m8�o�vL �=[?���[X���¡��7�\8�?��>�"����B!4� �j{�@��?ꐇ��|��N �Nf�/�1�̺ȲVٳLn]H�hX5\�V�||��u�����
J�'T�-F=��5���[����It-;��0\X��7���F�Iˏ%_�dzR��@6+.؇��Eu�飷d/Xqz�����d�w3ĸ����f*��P2��@�Y۔���<N�Nܺ����c�v��	��s'���I������M�ޔ�����@+�c,��)��σ�#��Sd�-��m��Yy���'򣰣�"l��"�����܌L HC��4��[Q�DN�m]�0І���<�F{�{F�؞7��V�/�BT\"I���%���V�ФfԥI�Ģr4���~l�WĞ�ï�3F[����[f˸�ff0i�c���Je�K%�0�����:֭'=M!Wf��hr�:�����(��S���TN�~�Wl��a-�W4�\f4�F�3U�E���z�]�Or� ���萬TY�����a.�^��ȣvk�!ANRS�0U��xr�{4S��Iv�� �y����n[oN�0	c���P.��y*�e�Pս�'�)�%yў[���,�E*r��8@�p�=�s����^��ȯS�rm��DK�������w_v�p&m��8���M�l�r�f'1� ]ɧ����(=�j���QLK7�����m��K� ~��
�'M����m����u&�\('�gVÊ�u7�y�+)`�u����|ЉJ�9X�$$�Z�1�!��>���f�xu���%c��8`��)�����յ�+�t�;"�f��%���Ni祵���:�D%�do��z��-�/"p��:�]o�%@~�E��������j"=�Ү]
��y%$���r���%�*����t��h65`0G�9k8W�`�7�Z2â��b8+���#���iXU���uL2Չ��߲rv���"Q�z�����H�&0�:ϣ�q�bu.ݴ�1��,
��a���_j���u���Yk�gzq��\v��^�5���:�"���K���#�Q�&U@�x/�B�$]��c�`����Qm���-O`��l���cwV�Sk�Ni���9��.M��]y��ld>�eu�?Ę��.RU�i��\B�d*�T���p�?��hb4��`�%'��̥�R�5ڈv�I�q ���H���<��I�o����zw���ᬱ@�;���Hu�j�}�8bW~��6KL6-\0��g@�0B�������<b���~�1*]d�7ώD�ِGͰp��9ۍ*wg��O��E-m����~���cI�E`	���_�@�2��:�?R�.���ָރv1�<�l�g2�W�G�Oƍ�X>�t�n��R�-�<t�$@u��
,\'L̈�?h5�ؙ�K2e:�`�<=Z���7I�GJŇ躠��N����k�&�����?�q������W&�A�4i3�EX�O1���	����WX֥cG ^W���6G6�
��',�6����-�"'����<$�s���b������~h���֛A��G7��X`���D!}E��ߌ衞?��81�+~�"��>�f����F�����Nm�P}iTi�[���d������XJ�Xй��?�ݕ�-��>1I�%e������VT�GL��n NT}j���T��H��ܦ��������+�*�iv�Wλ�f��w֚~Le�DL�Ҏ5M7�P]���h��]����AY�i�Ѫ���dQ�cє�Q�1�����%�I�m�����߉��̔U�L�D�Ne��ӓ��hEX�O{��Ǒf������~�r&�h���X�%�)��Òc3|��s�u���
\=���?
Jn��TǏ��5�mn5��x���� �\o���G��2Y�����b��~I�L<-S��|&:�O6��m��ݾ^E��\��&�&v�����$)���@� 9���\��R����)p_��c���i�q���.�9�eE���™R�Ok��/���6<��9`2G�4�����d��2��(����AW&���6>�UC��W�u^Ck�-�E1X�~�!��� @
��E�����y�!�M2�'\=���T�-��}��n;����c�̩�؞�Y���B�`!��1�hݑ�Lge=Ei����h~�L�b����yF
LS�T�E�ޡ��G*�k?�$TG>��Bg��� [RwZt�heB�Gn\��~F/�
��Tw����:k]���]g����貋ȃG���m����Q<�w�q 3���E?�R'�0n"L���t$�:�����{|YǝV��zI��A�7O-Ҧn�x�G�%\/�s�ڷ�!�yK�9�O"P(a����H×2qh�vN��BK��s���_��s��%�����������4@E�~P�0L����Q8���MK��F��8�`d1x%�t�3��:��,[�@�}:L�oE�X¬l�!=���+�pVۢ����Fe��Z ��;L�_{�>ښ,j�:c�,|�LN�9�Ү�z��G�g��Z��(-��V��@��� b��A�jc�S�`�x�( %xA�R?1�-øD^��=ٚL�D"�
�(0�n�c��Gɵ� tD	i�Yv0��"���a�8P�ou��z.Gd^����cG|���ܹ���SLwp�'';���\�1�*KӼ6�-�����7�z��ը���;rk��4���v(�����y��TP?��1��+�vxm���~����bA2�!j#�6�������(���*���<�o�o��^����۬��y�S{�eM��< H^{�_���}0j�������Wԉ��;nT)����~��,��(a���L�+6�~����)*�q�CZ�(��X���3&�}d�s��������� ʅ�a��=T�:=�G>�X,o��ar�OT�f;�0��ː/���nѳ_��x���NK`�4�>3�\[i���#2�Q����1��h�DO�0n1ZgD^<�����s�K�o�܁�M�ĺ��\H����T���ҽ���P'P�� hD6��V㵾�Ci$S�9V@���E �W�B� v�4��<��?%I�Z�{��_q�^h��˰�*�W��#%\|� ("a�8 5�����aű6��ld\ƃ�ElOw0��ˠ��U��)7�_�7�py>�_��	�,���e���	��� s=�X��R�{����0u�wC�(:�j�Je��	�2�E~�I,�u�i<�����N��V��Wa���1(��?j�Ch�r�9:{ŝ�[�j���W�����L9�k	QN��W��Jd��!c[�- ��먼s��.�u�^� ,OF�U�EoE��y�$w#t��P������̠��|k�}�0�b2wq6u��\�.sD�v�m�&�b�� y�C@6,�Oիד+��.�[K���+W�Y���KG\�:s��m�;�5,R}^|p����j5i������W���9e�m8�K�K^�S�B��_.N�Κ��l�� QW�t��n���R���H�#^�Tf�1�c���B�����D�CGO�~Ϲd��~c���>�!�q-�ڣ��Ĕ���ϋ�i
�u���2v��"�|�H]�IH(�����I`;�c���$��y�b�x~���!���=0�7�u^��1���|`��'$�P�@>�O?��!^/�8i�z����ل���{&�
��4A��>����CA��b�����v�A�<:�Ah�h��x��s�
2#���~�A5��EA[F)�%O�w�?�QxJԼR�ɽV�G��JR�y�����W�*5�����U�| z/8����"��@U�a�B.���ZS8��<�O��@����|`�U�sI=Lļ�k�=BvQ�� _�� s�f2�`YTr6��@�CD D%���"v�y��<Wq �`�Q;CJ	k�!IGSo����De`��.E	Κ�co����������
�" S���1�Y*������J�;�J����e��LD
ri�b&ž�����8PH��Sm^(xr+�n�%X�O7H4.&\�;�T����ކ�T�i�+r(�8&�K��9��2!	�cn�҅�����Ʉ���~I��'�[Mz���谡/+h�or�;���
������Y���ξ���%��T���(�诩�S� �B�Z�KN(�
&,�=K�l�/�%��;rY����#Wg*qi�E��W��jr�����eb	����x1R(�y�Q�3n����ISY�s��{$C�\�/Ix�i�.,(�v�R��y;����U��m�<�5����w����%�;�@&��g�87��Ӳ�{��W���NM��A-n�ٺ�_u���_h$>�5�]l0u�q�%��tb�$�����0�5����_~�@�dO�l��G���[�y�n�d���L(�RQ�-�?^ʕ��pK��������%J7�`�����{�o��T�p6����3�5�'ٹu��P>�/��M����w	z��hs���l,�_���d���$�FA� �L��J���IU�u���#�\dL}�!a6D6���*~��k���%{Í����j��?<Y^��? ��k8K6��8�B_)۴�₁�`=��>m��ߋ؎1� &�S��M��m��큅���w��,��X��'�_���ʤ�⯁���[�Y�K�*��Zϸ���6���E�^Q�*x���r�V=�r�t���c&���[5�_
d;(�[�%�)G����azgr%����f���:�p��/��@�L�ow��u�����F���來�H���jIT=����\��h=�V^�s4���^�N�q�
B��SxF����r����A�}�	pz�F��u��N ��BSØ�>s�uq<�N(9O�6U�LNp=�C�ް+�Y/؟��H�,��$�PO���k'���N|���ј��fx�ph�?�������LƆ^�H5����G�"��!�}��	�L��/r��x�\�������H@A���H��b�_��[FՌ))��=f��Z�R�	�0��zuH(�>_�|��5yO�&[t������U��+ҫ�A5�7t}�?���8e���E��iMƀC<Ug�<��[�G�&h�B(�b� ��m�@&F��｛�]țҀ���KBr������=t�n'�s�P�ͯ>��z��߶�����g�̲��l$g�<�B�������e���6sHah��B˰p���96F�вq���Lx��=��;����#pFg�Z?�/j�!�Z�%�;q��oY����	���Cڽ]E�zI�!Ԫ%8�0I��*zy��w�I<�c����dibΓl��V�))�(����	Z��/����Dޘ�d��vA��i+�V$+������|qD3�*x_rc��p��9�d���;b�}����4E2Y���B���k !�A�ut=�lT�h�⍿�����{P	�V�6C��q��I��NYœ\4�\��l h#�6v�U��຾ETl�՜������#��ni�)UT4gػ@n/ۑ�r�#�4����V����?)�Z�j��P/�����=��ե�x1��[�Cv�̦f��D�`��4�Z�y <%�	BZx�zH!��!y�s2����Z6?J�����IT�	�oT4A_��;P��W\�YE�=�GIz@%��73���0&	����$���*V�o-֨�E4�z�J��*r�#���:�S�=j�u�kb�"��A�X��m��.Z�U��]鶀L~f�%���s�fx�C�if6�_ޫؕ�ﰯH�h΃J��G��m���s�/�ԙ�h�0OI����a��-D���_���+6�j���N�$q���M�w)��. �0�?�+&��{a��o�Q�|&����Q�0�1��Mva脅{7՚���u�wڦ���5�)�ݓ�nV-�|�F j�v���I�q���:�Ȼȳ���g�&4�m��w��+��d���N%�����b�S}5S| m����E>�Y���w;t��#�$C?>�����YcО1�?�hT�}p5CV���9��c��$�J�a+;��f��7Y6f\��?�eūG�^d��W���Ѐ��l����"c+���р4Vy�k�lb��d��W�v�<TԻ`d��\]�����p}a���Y*.�r���g��.�p�6W�'f�i����N@�����NM�TO��8�ְ{��G`[`�W(��*����*5�_�
�-`]�#x �G�$e6�f�L�*�5 ���f����NX��&��?�����&���n�Y�Y��E� ][�����49�:� �-B��9���ECK$��v"a.��H�cp�-��}.���ݸod��Tu���!:?V�u0��}�at�/���to?y�0���%�J ]9_���)�2��S�|Yð�)*��T�@[L�:����kؚ=1+�a�N�S�®�U�_��L��|�����s���S�z���KN���j��6�X��:v�Me-���y%�<��鑸:X�n�z�QE��oB�ݍ�@~1���(�[+����4+<������on6r4|�E��8�c�jo�RB{ˮ���0�x�ڴU� ��:�59��eo�j	(�U����j�"�c>�'-�[/�NҒ����+촄'����[��S����H>�Yh��.a�d({:<%T�ڥ+�s�(�]N�R�<��T�3��>ߩ	��k	��k-sZq���`.�i�ʷ0 �9a������P��۾F�%��]�IjG��?��;t�?��6�� ~%qoj���|4�s�P/��!͗��j4A����\?��O4e��:œ�u��ђ��2KGN����i�᪷�rI�q��Rv�A����$+����9I�C:y��j�+�����gu;�jr/9�	l�/XM^�h��H��������:2��)�3/�������*]G@2�#B����[A��[���	���W��a�W�JI�̷1��}���v�3Ԉ�.���ڲ.8v�r���(]$;�(1��:� �0��ƍ1W݄�t��[*3����b�R��`��ں|�x�+�T��w���yQ	Q=6�w�ftQ���m��� ��R��f��LSD��������f��;�ȵ��qN���EPg�-�E츾r+���{U({�+~�$-�����kN7��m�ra�
��`�'�f�-�r���V�Zi^`��Wyw�=Ý��<aa����Q�3���ւ��i)�E�ؾ�}a��D�I�㷉8収&Uع�u�?C�E2��Z�� v}�QlY�JW����k�T��b͆��r�ޟ��b:{	kd�NE��ou���vE�Ʉ��Au==ʭ�W���Cg��\�P4��p�3;���~�4�z��N��@����9��c����v,6)~�ʦchY|���=�`j�򯲫���F��=k1y��~�����e?j���텊30��[��]�{Y�����e ������5�1�A&��ې7� ��^[�{�;����v�&)1�G���t�]j:�B1|����� �6���9�j�+ҕ�Z���ㄍ{/ë�4���M�|��
��C�`펤!��&��5(2ҽ��25�h��fV%�6��uO᪘yQ�iɇFr?���<f-ܧ�U�3 �4�Lڃ>�C�7�����(�pr!��4$t��T|��5qR� ��v�>¼��(�U��z�gP�d����)���M�p�GM�گzG�k�x\����H�ǉ� �1�Թǆ�D����������8�[�?�<�c�D�![*�9�X�`PC֢��y���G��uz�2�����j�'�+\���7��R�2�&k���~�����Pc݆�=�oz�EG/j�������twگ@�_�c:?�]��c�Z�p�bɕޡHN���;-@djd���,���+�\�6�'�*e����kA��<�l�{i5p��#g��Ye�`6�Y�eؠ=ɏ��b`�P�(1�-Ʀ�IB�Uj�LPyw��ԫZ���ܚO����ᘲ�;�)���8��|�e[q�s��?q���9����V��"�ݕ��$Ì�����p8���Ȭ��� o�de�2�(v�4��{xT�\B�X�βC�~�޳��p�X<OAe��M>�E����L~��oסe��vD9���,�5Τ���LkЏ���+	hñ�tV������ɜ1٫J �a��>��G۬�w��K B^�� ;v�g�ۧ3�f�L�"{\�S"����ڳH!��y�G0^�^�}�����U T����{/!^\c]>t�Ɨ1X���v���|�����!u�1�����fȠC��iX/G�տ�������<N]�O��np�������?�M<Q���z�G��X� �^�Z�n(��%���	1�gN���ٯ�����*����;�d�E�H��	��t�/���2�NH�g�s� �g��1"0	CU�S�*��l�)��7�7Y(X�w�^�(���&l����b��e���Ǩ�?�L�E�>�obb(����Q�c�bM�6�*���j.1P^�af^�Ϊ��ܢ��&�CԤJb��3�,���3Bg��n�����3Eצּ���+w����a"���7i�9t��4O �3[�a�PI��8|��"b�E��B�p�U@�՘`���x�-�/g���{����|K�,�WV�cf�GJ��*rs�^� ��C2ҙ5|�t�Q&4��0l&���M̟����?k�>��8�Y�j��[C���$��EQ^LVU�	��j�ه�\�o���9�T�nf���X9���˗�I[�"&�c6�}��F�u�u1��(�!��/]3s�̧׶^�O��DI$K���{g�t�DFU8qa�^͗�%V^��m��a���d���� �������)랱���Ӫ�&�9��&քK ���Ӑ�(S�`u>".�R��v4�҄�_*�㐩�D�$�J��q���[�4�<�%�I9�3-��~�4ץ'����z�\H�>{jPUN���S)�P����q1B3®������Z�\|I��ЬnfM�-�N�b�z�r�`-�?Uf#�^�w��Ǔa�ljW��Zs��U�CCC�M��/�El=Ռ��%��vf��>i  F̦ ��b��I��;ͪ?D�/��:v-ލ�����H`�>�s�rڡںu��*x2�0H65�Q�WX`9[��qf�\,����?Cc˦�ϳ�T�������h���)ׅ��#���F�ϙ�d����*bx��i����g5����(�x�
�C�Yt�Bݧu����۰���KD��w�״���J�RX	�� ��WQ_|��5n�M ������џ�a`�m؆�w�J��~u���]�|X��Xp(�!C�S�^#�E��F�>�E�%|�71u�!��
��A��@�(Hߑ7�G5�*fc����Y/�(�|������'j(�e�8~C�������/�܇��r�������9k�;>&��E�|<eM�0]ʥP���p��&\��!G�OI�%e��7�&A�|�p�K8ͨ�J�:_l5�����vT���s�����$�̠�����#U���Y��[��le��xDߖ/ϨFQ�m�'�&�i����m�yc�{�Y�&��,T=X�E�F��r��ߏ��	;
�VV����$��F�VX詤M�����]��}2�ت��N��*K�&R��Uk�r�A4��&�A0����m�Ħ 3E1ѯ��K}�mU��C`���������qV�J�[��ȶ������� 8��V��o���&��)Q��G\Q������m5�hW�zl���;%�3�z�����E�����޸2MҾ�{C��6,ω܏:��0�Ԛ�!5AM����1�OQ؞���Y�:DT���+�v{Aܐv��4[ji��֙h|1��3�L]cl8z�_E1E�mY	$��J��m��	|�5�T�\��L���^����8z]^�5���v0�,$5\'����~7�n\`�V�t,�p]�@�,6Sa���4�P��B�]���#5L#h�!�D� �;�Yi�����.k�4��j����4��%c��H�lN��iS7G+��q��P��v�ķ���$E`�����2���A�H��|aAG�A�vA>r�������v8�Lb6�bI�}=�].�`9-d��(�0az�B�Ϳ�c�8d���,�)���%���.e�}o:�e"�x�Ƃ0ܛ�H���F����*��Gf�;��V*�$*�rY'�a�l�'��vLʟ~�4���6=�����"�J�p:u}z����=�Z���q8� ������e祴�
� �="W��[�\5H�#����2����s� w�Z�]QI���x����g`'h��q��Ծ�3l�/2TNY�&١��})�l.@�7q���?�4�ꀼ�dټ%Z�j�|���p%�!R�f;��6왷�^ߣf�N�`������93_N�}`!~���{i@����߽U�ly��M�^D�:��V�	>wuᮂ_�,%�-?�'�,�p�,�x�9R��9g�9� (��G�^��\f(�V���ìK�VQ��ӡ�S�'���!Y����.�-t�yw��%c�ؒ'���4	E��exu�1��Y��t�`T��h��v@`��"}��VNy:h�l�=d�r������!��<�*���F��˴���_�&T2���VUa����_��#���ޒ֨	ԟ�'��cQ;a]$Q��rڼM�J_B(�ˉ��Z�u���~<F�耣�c�'��^�9�h:��@8� C��}W��%�I ���w�_����a
޺��������Q*+��f.5��}�\(�|>G�aV!�I�_�KId� �w�G'�ܞ�� s<N)"v���N����e�"��r 
�X��|�<r�vK%8�x]}SX �ݯwT�{�:%�-��v:c�8�$*❞\�����6���5�M�b�2[9� P����:��d~�dK]����F/d�	��*�Ԣ	s|
V7�\F�c�E"W�E���G@�H���}RӠ	H���=��@�٫�:؇0��j������Y!����/a֠���U'
�t&�c�������~��q��-�`�E���G,����>��`���I�y�d��0��y=JȔ^©f����������P�RV��v ���`��f��Mc��^�jW�2A�
��d�X9V� �kJNaK�]���U����U�xӼ,f�!�kr�j��lJ����I��3[�/�z;wZw��dYG����@�s�
Ǜ�ʟ\u9��B]�e�`�48Y����{�;��Ё�����K���"�U���˟�Y[�B6mۊ7�q�5;�z �ID�*�ؔ%n�r��0�8����8�����o�rD��am�>u�;i��c����k�W�� �o��vw@Bǜ��9��[�dU�oa���mU����g<mE'<�m�,�����e�E�:�^�.�>��?��)[�sK�㽒φ��GH�Q���؇��0b�a��<<Uޭ��܉"pF�D�>�K����ס.��F�����M���`$@^2) �s�Be�f��g�R�|a�آ���hjBF)a!���L�$W�*�B۾_���T�27p
�1*�f�uQ� ��݀6�?*Ϻ|��ī�@���`t60/��A�MϖrFJ���^b��%a�����[��M~ϓ�
7�ۀ�=Si	�?��1�iK)9�/� �ʭtD���^0)y�9�q�Ď��]���������,O�·���&���o��~���D���[��6�sȖ��W�߉gE��Gw��v����o��z��z����gޱ�&�&]�.B,�����:���,�	�r�h�Ud������)%+*���_�Aَ�6��5�ZDZEj7O��j��atOى�	��452N�D���O�C%GNs�!K��,��7�J���j��5Q�1��_�\3���I�~y��}&G*K�4��A+�����U�)Z�^7h�"�F�+�`^�:6K]r�6���4k� d(�U��zB��
k�e
`�\iw���ͨ�Ƃ��#��ӖV�V���TD���0>�"_�u6�E�	8���f��[�+��	J�>&�H:_�XE�$:^��V�K�b��悧�[�Ջ6�
XK�bu��4^�U�ɍEg�������F�Q�̮بr�%���(�"46���Ox�S���$}A>^o>Ɗ�ӃI=+^�'��0��Y1��d����p����7|G�}�>��w����Ȩ�^��G	X���������j�B�m���<�G1����`k �N�˵�da�g��D��Q�҇���U����!p�f�1���z���@U��(�tչ�'{�����G^>'��� ��Eл;Sd3���ش�)�#I=�)�sW�5x��=��A�JbGA�Fy�o���4|�KR|MI�;�:y�^��\��W��v53��΁ܖ�!���� �/�N5v�C����FI��4��ř� w�b�/��k��i���@S:,ڕ�^&�šZ�h�7"L�F�c� _*$2��lD��~b�*�αv�<m	�(��0�!nW%?�9>��%���-��t���ʹ������fyWBG /��L��d(�s�q��I����A��e�!
�u�ְ�_������'D�ɡ�
� ��9=��GrX��5[�%���,[��Իr�C/��LZ�7��^��=S{)�F��Y�5�Tw=^�m[k?�J�?n�.���_K�T�Y�� �HQ��4���ޠ�Eo9���xYt�3����O��Ē߾��C�Hز����ď{8aK�T�y<-h�$���cg��s��`���/DN�9_�S��Y��<5S_����M�Rf@�c!u��J�?5>-O3d�L��GC�ޯ��D��l��d��X�h�U����x�-�a��薌�#�����a,[` ��gUy#�tR콋ޘ�7������0mt��P޷!h$?v�@% �&~��l�Y�����ß�l).ddx����۷U�Q����Ձ�����#+�!�^h����뉑6&�Rc	�92�e�}�\Y���K���/D��U��ԸX���]z��#nh����5���&bw�AڢF?L�?������%�i;��ց^�?A
�z�T��t����ڸD-����b�7g�#��qc#��I>�&��ZV)X+�5;W��섩�n����Sq���c4�(;/���x�\91�����'Y�U��ݯx;�8�~�~��(�09g�As��~�.k����D��|��� eJ5%� k;�E1{m\tT�L���Jm�*/�ˎs��H*� rﻐ� D	��B�v���L����և���i.�8��:%CH�����_��]�7<���,pgv>�o�(c�0����7Eo�����!ʌ��3��#���6kA��h�_v���=45BP�+d��8A�#(X�F׍���-��Κ�^�$�-�`����;7�B����k�#��l_�F��mGtX2zL�$�5�o�֌J��&MЃ��<�([�� i|мk2�l�/��m��׎���͌F��8�P��=��H���ָ�e4w�m��]����3C�	B�1�b�>'J�WI�%R��$��:�� �Үa;ua��1���xB�](���9�Zͣ��L�v��ŭ�m�{#�Fe/H&N�K4�S�h�����M�,NN�&���Jz�����4�S'VO��Z��0>�-�hM)�?�ҽ�0v�-6�(���;��;L9m������V�1WXu�+�:��E��)7�#������G,�z�D�l�E'�EJ�YNBɾ�i�G�pGd�a����V��;��D�o�� U��+t2�=a��H�e�t�ǚ9"��_��Í9Q�
�N�>3>nvh^���ς�p���b�e�v�A@��1OL"DPS%!~Cv���ys���w6�~���{	A�����9gr�+��@���r�y?B�T?�=�C��DAt�7�J�3P��[���g��[ٯ�iJ+���b�(ԟ%3qP٬��Op�0ފـ���?��Pu1��K�LCx�0���a�#i�0�J12D�q_��T1q�����IL�������0CmlF�J ��$!.Bu;�ÎBU�WLߞ�_jgr�*N�ԃ~��� ��rVTN�
��F��:�p�v��"ܾ3R��=F�l�b�$�C�K���>f�z+4A(�� �cr1�����~ʹ;;��C���ˍ�M���B��=�ĭ��#�5�'"�;QZ���F�x�
2��?w��-���^~$@�1�|���
T�`0#2�6e���^�]�	?�a�/�7�Hiv��v|䕙C���Ȉ��9\?U�#*+c�BNM����9#;����m~�^ay#�	��4��@�WC5iq�;������i����@1�X�o�r+1�W�_�5'�&�>m�QV?$�I�'���"+�-��F\D�^����ˆ��q4�*g:���(��'��G�ݱ=�3-�Zg�� ZS���lO��^����}γy�9�*ˇ�k����ƨ��wkk�Mv�&6���I[<q5�W)>�����	+������'ItZ4u|������u������J���Ϣ~�!����??�i!�d�]y���`�M��r�ݢ�݅�4y��=�Ɵ<���d?��B��Ӻ,��Hx}�hKd�xT�\G�T��e��]��gSf�f�������Jad�򧺔�*S�(�_ղ��b����_�A^o�C�8�Q=����{^^(� ��;�L�D��l3 �9��y�;ꨏ��ʖ:8O T3�|v/�*���	M-Q�ݸ`T�]�a�A��J����i�5�0��{����[J��۝7 ��i�u���l�9�ǈ:R�����|�����?C�(��F����嘨�r�W���*�w7�.�����o-n�6���L�w���mՁ� �������k��.����Y��ެDŇ��:]uj�k|�n�f���y�"�A�����Y�.FKl,X�rǮZa�fJ��1�������"�'�\�B�Q�Z�hg��=������o�T�?�s��+h"��U-�{�"���(�����>,�K��]��<�`�>��#Qh����6�.�G�L�"���Q���
���0C��r_��ck`����s�\���j�ѱٝ����B?MB�1.D��&�(j.�����i(e-�b�PV�eL#�4�B�oH���v7TxD�����׉~Nl�̦a*�#Ò�	��|ðݶ�Z�8��%I�"�}�٤wK|��m~�'D7���h�xz(г3��Wxz���F�u�M�z
F$Ю�1� �;%� �`2��9M�i���Y�|w�=c?ڐK�x�F�%�u�!����jA��+
���ݱ�G�a4f���r`4�yU@�R�3#+�&�)����@���۵p�z��ȅ��NVKw͊��X:��>&N�?Tи�Sm�a�*M=�^�)�@W��=��!^t�g��><Q������~����CPL��`s|���=EB�`�6H�>����1�%c��s���c����r����A4\����b�75b�>���DIoЧ�=���%r�<jF�J���F��'is��������֖��!��JtYu��с<��f����ý��{&��65�%���d���k���G���U�W���f��u��f��zQ>�����:6̉+��I����h�XR�+�ݰ��c��J�J#:��/�^k��!�/Y�W��T\o6�9
�D5�
�g���G <�#Qf���y�n��,v>�%�W����~��>�b_^2�oP�s,>X���?��˸��T����f$�Mx �Vl�vz�:�������ǃ�2�TI�ɫ���ukx��{���0�.�t�$�8pg���=_ƶ�\�$�?�&X;d�9�+x�|��Gx�ɾvѮ/'y���~��S3�G�-M-�<l�x"pq�
oJ�;ya��D��o���	֊�lxZ�H�vp\��,�VS� ��D�����C(��x�`X����JD�s O�:���nz{E��=�c�G���).G�<�.~�$�9���d!��C X4AG��}*���u �0oʤ��1j�d�����5��H	����5ow���z�ԝ3���|�����Q�~���%�u}��.6�� u�չ1��B��?@�����t��m��8W0�Ҭ���5u�W��^��;��0��!01�if4�?��W���+��.�j��L�	�!R1��{�e��qp�|Yn����#wh �+S}��Wcj)�ʑcMz�Y��cu��$�G�k��ӧ��	��V�9���@}�%�p�
mD�B���yÛ��}P���p~�>"}�K��d� [ks�������o�.b�(��ƒ��4~�|:f���{�xn�Q�1
Р�+�W�����6��tԔJ V�r���N�]���w.!����e�	����0�`�ɚt	���V0; 2ϩ�9�~�H��b-[:c�J#p0�Rs��iX�� �"l��'m9Ā]jqR͸�',Hz�<}�a�:}G�t�S1��(�Z<��p�V����	�7�;���?����1�Z��y l(w�\6�` k�m���Q��Xb]�uB�gx�-����Y�Ç�:q O��Uv��o�?_!�=�$c�,# ؤ�G�F!��rs�;�+���������m���o.�tؑH���c�4������! �0�Nۻ��<��X�'&f,r)����NH��b�<yf�(������r���V�x����$VV�V�r2	#l*}�4N�J��������~�7ݛG�ϻ� ��z>8�,�Zz�I�S�w3����%��c���N���ƙ�ƪ�̂��s���&-����t&y���C�[Y�#V��>8��{�_�I�5���ـb��by䷳���~�+kƸߍ��c쓛������YI���/[�EO��,T����ݐ���h1���`��D��4e0���������_� mN?F�����"#9���t?40T�r��
��,�+�yZ�7�f2"��X�"�䕸��a�� �DZ����~�U<�c�җ����w(T5�֋�󨫭�	�?#77r2�Vm�ɝ�q��Ux�����7�6:�q�
 =��$�Y)ZaOo����@jT�;�G��vGf	f k��>���A�h��R5v��VRDE�s�	��@M=��=R�7@5�%�]�&��Q]䒋�$�+\4K�{�����JA��;H8./�Ȯ�Q]/V��q��,��'e<��ȫ��9��#���!V{؞�hǲ��:�EmƆr�h�Y���AL�(���G�� 뇌��@�Sw�3�Yþ��5����� N�.w�WL�.e%�>C8	�dZ[������9�0�q�5�0;VV��9�rށƦ+�V,���`���y�y�7�2j�+�ͣ�>��\X�&��r��|Dp�0y=W*sŢsr�K[���Ÿ�
�{ֿ��QA'/��%�X"�r��e���[��Z�P�W����w��m�k5f�+�8�����o���9v�N���.�����9Q�S"u����Ce��e��N���T8�:B"jL�D�: �D��<S�dA�)Xw�χ�x5�(د���pEv� ��D?QiA�'
{�
��ۍ� s�|:���T�qЧ��T���u�J���h���߉Ђ�ͨ�������������k����(W���g���$Tۘ�/�k���|��V��|fx& �2~a�0�>Tn���������kC�3Q�}�u>|!4=ع���E��l�X�Ō惌2<I�3�@f�'� ���u҆d��(�8��Bv|�b�p��p��m�����j@���H;�繌��^%EѶ���1ǃ4N#P�>W��͝sӫ�8o|Y7Zq��yو�u�1�#Ur�Ŭ�=$P֚~9UϤeE�P`��M2e�W慏9��#{~�Nw��&0�L32oV��Y2(b���B(�n&�����h�� ��Y����7�'��3SŪ�bW�7||�ж`�x5�����4���h�J9Od�,�|�D��n������i,^զ�<�'�z<�9f�L����M?C�C�
���;E��m��.���Qb	�&���ȁ0�p%����	_i�]�kaB�ZI΂_n���$�����5v[\�H���s;�`a��}27�c�N�����f������z�~EK,�	1
��$@+�M�^�w�+�E�U�S�剘��v,�hs*�<	DdSB;�kܨ4�]�m5H��S�4ǝ����d�=0���g�:�j1Z0�#U�Ո������>eD�8�&����y˧?�E !ƺ��q�7.��Q��bz�ڨQk�MTz�B�jj*	7���ON�z�i���M.�(�&����nY��$�S���;���`��G��n������|�*"J��T�������إ��o��=��_�>���x~�,~���l��D����+Lz�="�9Q-EJl��d�_HxYAj/��W�����ݭ�:��Yic|O���?.�,#��x�n���$p����%�J���it�ƚa���_f��#l˞�F+���=��\�<TW��%(�� V�w\���[T�����Pr�@���g���������I����5f�j��!"lmR��o�4�x췒�\�8��w	��7������v��\��}��P$�W�Q��pD���s ��_��H_�u9 Ź:�����Z��Q�,��q>䛺�@+A#X9#���;%9qz�y���)`��<�m_��,HdeyQ�J���g�Ǉ�	��q>�Ȝ/� ���x@{�F��p���<�#��~�H1��ص]�R��V�;Z!���:��"��K�1g*+>�霝�;ƀ2U�q�ˉj��<6.%��<�ɱ���1b@I��a(�����Nvh���X8�"	�Iʇ���Q��� մ�1����W-�r���W���.d{W��9��-�_K�%���wI<������X�lXcCs�4߀s�/ʵNڢ6�AP����n�ez|����F��(�Cw�ǫ��a�2����HNh5���Rɀހ@�Jv)ndAt}���#nه�/|�v��g�����JR���J����&��� ]=l��"���7�/���_J���Ȣ�r��+#~.�~,{y N�d/������������);��5��sg� Y�&}���i�E@������.�W��O+��׆Я�f�#�C?��� d��������&v0%l���=�"ېֲ/ �l?�b/F�K�<r�۝j����*�p��rV�:�`36&�L�}��\˜zL&�k�)�Y��l���r�a��4��P����"|����)��A��(m��&�*N�������'���Y�ܴ� d�%VگAGJ�Iμ��qE���8T�\YC��|NJ<Xoz��.v~K͉�o���ݱ|!�S
u:�r�be^��1��<Ά{�S���&�5^
ЖPn�
������h��h�w��v�x��i[97��í�m�wzJ�'�.���F�{$A��}���vF����DFQU"*Z�T�W��C��w�j��̲�|���T���XNZ��I��OϾ��*X��5�5��q(Fe0,��JID��';���\�x�{�\!�6��~�D-`L�;�R�iw�D����;�j�1U���ؓ���R�Kw��6��Io���t9��ޡ�����T6����9��BQ��v�uRL\��f��h�=��'�>��cF����ni0��>�
�s�q�9Z���SASz�X�)%C��u33�c!C���"�:���}GeC���)��"��k�ǃب`Qmnl��-5G ��Y��?�nP@��m�~�&h���L�Ad_���;VQ�	�k�1P���D乛�7
.���+����d�:�}]��SmV�=h*P4�q)�+�A cUw�C;�q��@i�*m�N�WcՕ/���W@�ӣ�`����ap10Y96�U�o���QV�C�N�����{˷�C�o1([�hQ-a�V�c�d�ۓ�%���"�M1��禼\�c�ч#�/�!��3��R�i�����$x�X�zᶙAԡ�
��
��Q]2)O�:��l�4���5�U��-��F � e8�ˌ20�(�Wu�@��d��_�p������C4�x����l|����]��Vjt.'/,��pYx�ճ�!Wq�aU+@WP���,�����=U�}�T�8�1�*ѝX�������E�w����wu��g�zV��/���]�m�N�<�����1�*��x���m���¢�Z�̥	RX�'j�����$O�'>�E����	���ʬ�F6��9�?�s7 �/<�"��pcʏ�#�'׏=x����\܇T:[^
��r}�#�.����'���/+�<RU8�f�_(1��C�%r�n����#r[�R�'�B��UH���u��ט�ݡ�3ͧ#�mܝ`o�20�K�`�I�m?F�&:��O�s͆v�H�ZJ%;�m��"[+��i���q�@ <tXS�Z迋3�B���� w-��t�3�*�Tn�Gf{Z[b��2z��[8�w�UӇ�j�Ǫ����8 ��ydtA��%�d�Z��DO�����sR��!��� �Si�>��U��e��Xi������2�e�5�	�.$&����0�P��_�܎m�\�`�kM}�x� ��!w��P2�<����	��{�.D*,�ҊHL���	$�D��:AZ����hwQkp�ж68���JwCd�<�B�?~��Mn��en!&�?��t-Sd�� sBF�����Qҋyx� �4zboP��H��>0��A�����!}B�(2��9�9'�D���|��e	%jo{��P����"�<<S|�^2A1)AT%�ƹ�ڎ�}�Hp�Q0/�������2�Q\�J�WV�{��Ȧ�[����f�Ih����Їm���i�7ӝ��V
��V��W�W���j��C��ȅL��o�7���Z���	�g�HLZ��y�̓%�U�~)�A�Zz����I'�w�2h�[t[�h�� L`>�Id�}k����D�5���b	b�bUM����c�3�����*R�<eK�s�V�'���Z�k�
�hO��j%j�ٲ���;�A�;��܌#hG�T��1a��Q�v\�r�+�㼨�'�����&:��E�7z �e]͟Άk<�$s�;���fQ��>��<�ݴ�/ �[`�x��-���8ʩ��pT�=��p�!bh�
D%��'��&��7��k�������f�r*]�YC�����|C�c"�v�m!��9���L'����*W����%1�v�|��yC�e���f1i<Bx�ü�Q֚����!>�}#�?ԡ�vo�r�� �J���c����キ3�6��n�'���V��~��۱�	�ㅓ�=Z,���cF_3��ɸ8!JB_�������'D�@F�G�f��ML�b�c	��Y�ɵi��#R��dn��
sC1�Q�Ї�vj�/���i7X9f������\�=�����G�+ܶ�'�aS�A��a_��2i�:<P1��w�Cb�y�����p�)N���|�Y(���#\�Xf �!m�%���2'��=لH�����mn�<j��V�f�Q�WM�?R#�ZB���=���%e�u�y����8;�=4f��T�����3������� �G�#|�t?[�� ���z(���Z�Sk������k�~;sS�-���n��µ"�G4�L_)N:��C�m�X:-�7Ȫ���F��ӈ*a8�@����e)z���o�_��M�]!�V�i��?+g!�v��j�p=h��n$A�j q�M:�7m�&��AGk�iw�zAX��4y�l�=�]���vX�%T�2���%,lY c;w?`��WK��g� �A����8���K��ܳ�3��6�*��w[���NSO�w��ۂ�P�/_������v�<�R�f�D	�v�������ӹ;% I�.��Ƌt�/�cY�}�W���;�ٹ�!ފ��2���'Q!2���S��|,�<!�F����- g���gM'o����E�iK��Qt�῕9�z����3���f�D���F�F��"�^U�����O)���nG�y �FʞV_ꊃ��*��z�|�����L�c���'��[�O�~,�pSYq��@�����2S��O���k�{�	��W$���Ƀ's���9���?b��Ņ�����U'o��YC�O+�EHy!� �Yq��j�&��.)�!��`��7�BM��>���r��r��;U���6g��S��Qe(K��M�U��7�Z�R}����D�>o]�45+���V�u`���^@h�Z�,�"�,97Cx��:2	�ӽ�����z-�>n��^]��Ч_H���������%F���Sli��E!�ߧx� n~����j�}���:�u�gE�P�t�;l>���gs�#�Ѳ�s[lC�O ���VQ�-�i�����7h{�F4�:��[��؀Վ��}�a"j �s�b��<PN�>��48�mA�����;9�����t���T�0�v��~����Ӓ��8m�JM�ܒ�8>�.�g��J>-KD$�~Ҹ!��m�1�����������
��8��ww�?�Ϟ�?D9��: �᥄L,e��y���t�g�I������%���Zh��?.]Kb�7�X$3v������kL\h,7�����|]��3�\�{E�����M׽Y3�s��k�Pa�	�:O9����r��X�"TJGۢ���8M����݀_���bC�O߉�}w�j53�[|���?2]�A�~-�Я� �U�w�GP
���Ɇ���~R	��'"���?����Bx GEԴ_B4��غ�7l�[#�����������c�K�a�3n��p���~��@
�`h�{�][�_��|�O1xD�_C�0�����z�JW*e�s`��$!6}8����ԆA��>|��l���కS�p$	������	Ca�+�K�g�)-_��yN�ԝ�YU�ؑÕ��z�
s�*��V6΁�-��F�U�p�]� ������!�@I�����D�������Hm~{�{W���J��x�Ʉ%i�_Q�Ch�K�2����;S��P}㯹���	�%(�O	 �R�g�g$�
�Q����k��=,=�(b���ěV�g+�X�����d>$$�gHs�\[�^���+[��`�]Q��wCG75��jF��ړ��Z&�䑯�_V�a5�H��y§�ؘO}`�����G�,wa0Xu��<�mDlME�'�*�,�f��	;�YD�ҵ+x�;�i��żƜ����ږڧ*�XQGK1�#����ܼ��Kc̳\p˶&n��������C&�&6[!�6�(�+�m�pn�l��D���#����h�%N�]�,��/<�7*� ��֫���0'f�1+ٶǹ< T�˾�؅�e�AD���Gd0��jZZ`����Ļ�t���
͕E!�����W~���x=F]Q2�r��	`�<���\ Z46�Sa(�!�S��~���@s)R�F�2yu4�	̴/��Դ�$0����ohz��*���?��aԔ� <�9C>����e���R����8��+L�ӷ�aZ"��
�A Z�ʠK�(犝�2W���Ƞa��������ܧ�PQ%�h���v�:�ܚ��H<$�]���j���q�?if�v�~0u�ʯv8���U?�-�~R%{ٓ�/�e��{��~�f�}��G�}��ɠ��š;>4�=�������<Ai]H��j�*�o}fy
~�S����1�����9Cx��!�Ta�v^���ۑT#E��B�Ky�[��k\���l	/�'f�^����9 
����oy�B:�z��{y uoU�.�^+/������U2�}Nq����/�.��A1�5,U���l3�*�6iL��Cq1q��7q��`�+q��M���7tzZ�������x�I�1�Gs�.�:�����e9�:����ʅ�pC�@*ƙ��1���7:����4N*w*�=1.����vU�˺ ���{��!�.�z�:��D�d�(�� ɡCs(�p$b�oHYf�	�nE�&8]/s��Hp��]������fʰJT�}�xA����ȅ�B:̲]����H��_��b����u�¿�����D2n4�L����5�,u <���\(�_h׎4���V/�����邲�G�S�G��}?����ۣl�J@��,9kb�2B)�BfaZ�=\� $_O����5S�BS`A488	NgE�Ԡ���iW��TU&|��&{���'�=g@���)����E�� ���dΩW(c���(�ɬ鷺�,����