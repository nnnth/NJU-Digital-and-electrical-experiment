��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��op"~Ϯ�!Z�	�����0�q�(�q�S%�z�(Ha7y���k�Y�1R��lK{�T�{,{��M�ac�@s)�-�����'��ㄐTce�4�0@e�t���X�8F�δ��7S�Й�Ee�30!ToD�~��(Ub�S
����:x�myDD��r�d5��,��9�9nὈ�Ts��G�I����͏��>kK�v��g��1����9C���aR����n��x���D�7�n��Ń�?��И��[_�g�I{��u��\�Dn�b��]Q���= ��;�]��c<�7�O�!{����_u�MJ�o�1�
D���䃡}͔i��aB�O�������:��X���)���rV�4��W]�cl�����"�O�Hc�Z�Λs�+���o`&BG���K恋�x���Cv�\-��x^(�S}�\��h��_��'֖{��1�$t�ݤ��*�L�V���A8��=f�IQb��X &��E7"������چ�	MT�����v�l�&��G�YNbx��J�D�������\ q�~���]k7'
��� ��.�!+�e!R�$��P�N�c�%@ݪ!�d�э��q�m.��al1U����^*n;�w��Rhzem�����z���2�pHW��l�L����/���Nq�g�������(��ˈ)�л���ǵY&���W@ٮ�?K�F`��3`�G��϶˦Io�Zc.$LC� d���uʟ)�$�x���<e� u��s;6��&b�Y6�D��PS7P,�k���ԍI����3�;{����*tq��U?�||��L���	 L��C�Y����m��YOv�U��L�^[x�GJ(�~�ܨ���YG4�-�Q�東49�0*��gȠŖ�$��&�u�F�l�)�/QiW�!�I�ryA��<,��8�Wl��ȯ�E�N4�{��&�0:���]�~��������3^>0��o`�Z�D����V�S��6�x�	��������h9]��`�i�H���	?u����;,�y<lZ`�R><�q�lO˄w�'�n���}R�A8��rG$@�f\'�B�r|���ꌒϟM�� ��E)����u!�n��s�uu�5~�}��a>�p���d��tVz�����* 6��޿"w��z�R��H 7��̛��{��N|}[���9�E�\�c�u���U��Q.rC�0��pw"F�@�t( 3Lٌ��rZ2Cl�z�i���4#�X\����/5(L�`JB�M�輦-k�r
�8۠͋�6�z|�!�->�/�U�3��j����W�X@���Si)���:6/y��}y�:�!$R��-����"���U���'�1�a���>qv�lJ��N��"Ϧ����4,���# ��-�X���ڐ��;���Z��&j"��F��I���e�^O�
8m�y�Y��V!���I���I��?�j� �-���J���׼9e�\呪R�� ?��
ȡ<f00���^���'�*Qm�Y��	9�ƛ��	�l�u����K:�'Ұ5u���VX�9=�Y'���C��1�-��t��aN�f�*܊-X�h�������X��f��� ��7ğ�0*c�`H�T�=��8'����:2,�# �+u���:ѥ� ���/�cv�u�,��g�+�!BOT�8B��T7��Vl8Mw�X�G�����A����P�˜Z�/�ǆ�"|��s@R�m~zMk���4I+Q�������J%�J��e�V�zF��n�f�[?LrA�&��&/��R@�Ѹ@�G*rH<<���Q>	aF��R뺠�.D�r����m_��ׅ�G� �RPx��4�C���_{����$"��1,��uF��6����j��wOkd���9?�Iԥ�٠��Ry���}�'7�����c31�$�>� ;��ʮ2\�LR<I?j7v��B,j�0���HT��.h�g�$o�{��]�=�b:ez�U~&��w�6�������f��\'-�$V3I��E��5�w�'��Y^��Y�Y+���kX���_)-y��P�w5GjG7^���D��%�|X�ޣ��?���@�J�34p���Țc��7��L��6w��LN��$��jf�++&��bt����N�3�
"9/:���s4ob������F��×�����Lw\���37��m���S}��D�7���+��]m2S�M֏�Hr���r�ʏe����\�Q���?R��J&�{�O�
���AG#� i�#'?�-e�I35����Ѳ]~b�\�g��<�\����J��,���|�/��t:��y��Q����.唉���ԥ��*����㻦?�z��:2;@���X�`�dn.�r�"��:-�ɉ%NpyǾ��7l����\t!*�T+��rfo޾��@3y������#�cVS.��^��!�%/HR1�Y*g�������i�a�(��N��`K���<�ԼK�B���*��B�t-X����	wB���V T%��QC3�|IN}���]	�t{X;���%���`�Ǣj���u�<�]Q.Ă�[�q�0�i�k�l	4�8�.x�]�=�x����۟�P��"a�ν��4��D8R\z������6�ey�Y�ts%x'k�_3|�C��\�Ҩ>9<��Ȃ�V_���䧼��B�2�
vož����o�5*4S���I��6&�{�g) ��TM1�Ʊ%&�v�nN(ߕ�����c��`���t���y��?i���l���uRE�n��C��� �-!�V�fc��zɐv��Xn'o��FKq���z����R���yʋ�N9 |�>��2~��P ���B!��Wӵ�]��d��"F��K��>?Am�d�����g�H> �"��ힿ��0��g�������E"]M���j��ꨥ�OLe)��"�H�a�m�3�C�Sְ�����n[���|��<Ͷ5������ӕ�b��H{��o��Q����	쐥UUZ�(��J�z&~Z=7�55�3�v���<f�6�Sx�]%xT@�4@�R޿{���
�*�=(��n�q��+�Sb����ܖ��8�dp$  ��c�A�(���);!Pb�{UjL)@�!o��������R3��
5�=qV?�_�"����rG�n�N�ĭY��r�e��f�s�K��/g��*{�c-3�oW�_����!�W��Ӻ�4�.�N$h�<��������%�\`�p�wU�?�Y֬@<��Np��Q�O�����*���H(��a��lt�w�0��w��1�~��w���LZu�(sFx�0�!t��RQ�c"a��$����|��ąq�|��-/���0H�8��Au<O�oB�3�yT����7J܏�}���7�*�(v���u'.�����^���J��RK����Z�G�w����)�|���;�3S����\�mܮ0��U�6�R�q�du;Y�$!Ԣ|����-d�ռ�شy&�I���WBdL[���i!�[�r(�FܙOQ�����r����=t������?|����m��qU+��B����p��菪��	���H
*�$%��P^�t���~jX�����F� �;w1�&���QP5��ibv�;mT��G���,l	�mkG \x�w�Щ���|�h���p:m2��l�ЛX# W:�D �7�������
���c2�6�X��>~�⇑��/��`
<ӎ̃&g���_�R>v/?��Z���^�<���9��a�U�k�#���H.j,�&+�2ׄa�ؙ��$��SGa�@���+}]F�Ǜ(Qĥ3�PW�AV/�"̕q�4*�Y���/�J��CZ%n�[�HM &
_���3'so��
6O��,��%�ߣ���T�D�I�]h��\Q
��XS�J���mC�?x���<Y/�㳼7igM�|ת���q��`����&Y��T8��Y�.(c�����qBg����2rV�u�u��#�=sBwG �:���ۛ�g��jh��x�\�#=Q%j�D�+o�^\���v�U���+m�����.�yv�oJ�Gu��m��fO�y"l����('����y���Ꝛ:@{��'���D�b�,�"F֮u�n������H\�cī~t�~p�^�}X!���HԲ{S�=,�U}I��>(�tO@VsH�n�s8�1�pNc������NX�=�@g��+O��Y��|*�u��Pe/Qv�R�!��z�A��Cxp#���a�T��`�z�y4LO�Og�RJ�C.k"WbPA��:���K �ü0��;�wl��\n�42��r���Y|�N�:ݖ�(HXy8+-\V�DV��s
hy/���k�5l!��ju�]Ӌ88¿^U����g��Wǣ��/��n���	�83�B�c��c�T����RG��u/?�:����n�1yNz��,�Z�`j���ƋG�F���S ׼*��Zz�q�(5�F�'�����rݎ�s�6VC���2Y��S;�6>��#&�`�sW���c��A)��(�ZB���'�x���_�O�m�gag�E��
��anJ�6~��]@�	L&�v�d,;�ɐc!7��w�Q����`�$�JD_�G���
$(��.�	Ơ\��Nzy��y�kd��,`Z��!o�pf��P�xE�.��PPL�k/��	O�������e�1�9�@����v�������yiq�x���+�8��(YLɬ�)��<@*��z��e)�.�:V�Z�Y�G�^*-c�K�jNUwJs"[�S'��+^� ��Q�##��*��4���7Sq;�#$�Ɵ������*F����m�D�m��穼L�ݾ,��$��ʥ���Tօ`9�*��.P.�yM�D8.�%������D��r)�n��g�󛎗-׉a)�NK��k������ͮ-z�m^	��"�&#��1�5mk��T�ᤚ�/��UJx;��r�&����#��9:�{` #��E+hA4m[�|�HJ���~���M�����Ƨ�-6�^ؗz�<GX�JD��).�6�n��Y0�~ة�Ujbۅ-�E�B��7����b�RwZ�'��2�� �^��
���{�1ᓝ-P�Ԝ�,�Z*�-��+��j'I��6������sI���p͟B���U�̇����9��P���������+ƛ��/�`���:���2���{�N�)H�a�xe���}F�����wx�3�oV
����G�?*�_�N����r�g�1��Lch�(��Πߊ����H=��ڛ�i���u�wz	�N>��)�HOT�4�B�q��,]�Z�[w���^�
��g�O�Ͳ��]���������n����!t]E�X^��l"��B��1'D�B�#�����_�Ex��ъ��T�R2�2^�?�)$AO�ѯg��i��A�6 ��[ɯ_�)�n}�:��J�yQMn_OK6������qE*N�uI�5��4��Ys��+�J��M/ph�sç�^=�-|���D��C*��[��Z6UC#���zUq�U��gu��ѧ�W��\��n�n�3z+O#����;���=5��f���q9Iӽ�صV�H �7h%���ш5SiO�������c�����p	/��0{��r��Ӿ���v��`z�v�������î}�TL�\���}M���f�Z�;-��ǆTv�Wۆ���W��RE��e��y����d}��������q����fr�0����;�H{��87�������i�.=7�׷�C��w�ʹS��\l�>���{�&E���<���P��"�����<y���8u��Y<��J�)����4t&ǒ]��j��j��������w��=.�ݬ3�����}u� ��+%Řͣ�p\�C�}�ힳ��3L�:��m���?7�sϜӧT�ih)�[)h�X���0e��p��g:{�HBtĠ���C�H��iAЖ�}'��Q��4���\r��{q�6�ު��ϧ�~E�ڀO@Wle�2P�]��z�)y0rB��A�&��l}G���B�O�He�|F�F^�)�^���j��ɞ^�������֕��Eχ�	���)���X4,�a=y`��Y,�~���Vt7�"���c��t�^�5pN�H����wG����'T��.�ۈ��S�R����=6���8���l�l���<$i�R����� v�=�;\����%.����FE�����Q�����1�P�e�f��xQ���+�T��,���9��p(gmV7r�_,�i.b��w�f��hF잾�r;����7�-/�e��R��G>"lySl�im�±�'�O�KG=t�.p���!����JS���+��޿�Z��f��=�8YF�a���,lXf� ���n0����;�7��y�Z�91�]�#u"�-��
��,�o9��XK7��ը�F�j ;������z���	3�Ww�ۡ�i����5�3�}��y�Z�	��HAN�!9	���A��4���4�T�S���<TB��s���n:�2G��QL+�i��2���Ťѳ�yh��z��I��BK��=t�X�M�>����DQ�w��Z�Q�x����~<���3�7�̊����	�I%���7�����f�tk���Ek�F�tj��T�;�&yY�ޚ�� [2\8�8�Îq5SQ]�ٰ�}Qn���D�ӻ�ȲɃ�dߝE�� �&	��Y)�@�X�,�
�$_��~��{kż�uƇ�	���ƪ�0�?	���*�j]Ι�
h#�G�@2A�3�<z�
R��,|�t��ip��%}F�.4��4������<��d�.˹|�2�%�e7T�Tk@�FW�T���v�U�η�I�����ww��/�ʙv���~�+�c��^Sm:�ּ4T5�b��ߺ�uo=�~#K]��>��)��Q <�U�̫��a��q*�>��bCm����UR���QBR�h���ֵ�����lEɝ�Rf�) [&��|IZ���Ι�%�^Ad�jtR]=J����g**`7j��c�{P���з��4��<�TP�H���3�		#JJ�����Q>�w�����`R�{?9nG����[�E
��
2�%C(�l~Pt��I.�p�=;��L���`%�Z��DHț�$����U�V2,b�W0�`@{�$E�|�]�kĐp��Ų��O���i�[tv���� Ab����C�xj�Y��3��1�/�U3���T�O��(J�䘦V'O\�~$��f��&�� D���,��$p"��_�u������m"ּ����3nf����K·�D�{�
�O�>ZL�qฒ�T�^Ο̵���"�8����K��K��4�Vvq��H6���G�Y��kN)V�Q�WI�Ѹ_>c�B����Sfi�����i�ð��%~\���2]�<��t\լ�kѴ�d1;��� �ޮA��$��A���h�Zte
�a4����E'�s���bƧ.B���ؙQv�{^�5u�a��>|(A���9�,��˒{��4��spVbv������k�R�6q��wQ�~tCh�u8A&��z�=�<-����A���*M��v�n�p��)pm��c�D�8��`�'�XÙDO��6�k5?��3oDiB�U�k;M3��m<�)��W� >r=O�iC�`H�&�4��E-R���N���� I3�/���q��v�3�83�����t����뙘y��У���Q6��2����l<��}X1Nj�K��."����Y1�b�����V����2� �`]�V2�[��7'b�x�鬻U�z�J?��	�"b�� �9���DͭF!B��k��o�e3��.�5�%)�C�J��Eyj����
\�ps�����ֹ����>�r&�����b0~�%��x��%[\f%�]�)�� 4=�L�T�_W �j>�5R!q��w3��o"�F<�N%%�@�5�F�~.�1<���E���U�R��+��)px��fy�5�� Id;��p�X�Y�{����_ ���o����Ӗ[L���f�{�2?H@����l�)���*b��$�W�T��x.�D�L1-fK�2 �"���Q��u���r�m�=
��f�dE�Q훘�ɂ���ۧ�,���x�ߞe�bL��C��'�]9?�b��^���p>"K��k��_µ���W����{ =�P[]�N����w9���e���(�_I�J�k�H\ՐP���<,���g(Xn2`IF����h	�RR�N��6]
{W���&YE[��9[��Z,� ��G|�CW�_ǭ��'N�����<W=���o���aG��xn5�u)�$��>�:�u��T՝�g1��xYb_����$���ϫ�Fa��<���:e�K6�2w�BۏČn�%^G��a�����Ч�P����}8	�(���ӌ������!�[|Mb�#�S�_t��# ;eCX��ӓ���{^A���{s�g���Ơ����%C�������$%4�CE�4��.�3~����޻���[�B�.���\���џ=�DI��ƻ��߬�#��U�[M��ꎢ�Nu�\f^hϛ���g�`b��f�k~Ʊ,+��Zv�a^�����᾵��&[��٢d��4���l9�>��a~�4��y��RJ��ҠImUT��Ԍ���o=�j~2�w
0D�R4�NjZyߓ��9c��BJ�J��jYw�l�9jٴ2VL�9�����r) �FJ2�A�©�B������77�'s�m�Rij`)��� Z�|����fW.���L;��[���b�5b��E�DK<�h~k<kA���L[�Vh7M��q[���r�-�7lq�/{�A���16�Ip ٥@�T�
������l�ڤ䆟���ט�+�i2{um2����Nǖ�O����a�ڣ|}�,��ax�ߟ��B�!ڠ�4��.F�&���sXţMYD��f��fV$#����m�f;/;���jp���,��e��8G?�*�;:Ɯ)J��zqʥ���BG:+텛p���|�I�o��)'��5��eø=3I��a�x�a[Q�����>p��-�?eD��+¤B����/io�	�]�() ��%A٭$�:���ď�E���RR�<5���<���M�L�V>2:�c��_�s'L::���v1A��G�Z�(�]�=�q�DA�����6Z�#Gɱ�n�����T���
�� ���94��y�Θ����|��|EM˿W����%RW E�M��4
�R��ɪ�݋���%뙿���G�P��2.�ĩBU �ƶ�6\��j:�DgD�Dیm��d�J���q�8�u��sQ�1$�7&nA2㱷t���p62D$�,md)KO˅׉�)��L��a��h[6�
��,���=�{wV����ϳk�#l�\I�^�٠i�
����eS&ҁ��?#đ�肊 G/��U�6n<7X�vZ��
�u���1��G�c��B�T_MW�-�<�J+t	|^�ݸ�@:������N���0�F�V���i
���U��(��x���'������oE��z��7�˄��m�[��,\���݅VQ���l���ӝ٠���/@I��r(�p�m�� 4Kζ�1���
�N��9�#�/?�,���*W`��
[�Uۄ�{=�x"�k�ct��u��UT�	q�[$x#*� ��:�>E����J�"�c�����ê�`�'1"�PۿJ��'2���Zb�?�������.�/p$M���$�,$r�
\`��#���M�c�����Pn����#��Fr�q�O��~����R^����,btyoz�?��ϫ�!��	��1qI�ѓ�xU���X�Y�@?�g�>�8M0�ɖ���ÈD�:�xJ��;%��?]�f�@o��S;;�S�Ϭ������1�[�1�ыo���JqmK�/Wd���Y�A�rM����˞C,͖�g+m)vW��y6΅�yVmښ;�& L�ؾ����d��M�}_����mV.��gA!8�]!I�3��ؠ��:��x��@���`V������TCUf쀌C�p�/ʺ���g��)>�/B̈́��o=<�œ*�,���:YI��|q�wVn�iIE��0��!�$|�S_�h�n����P�u��H#HƆ=N��kqb��	�Clްmظ���(}�_ʬ	�&����@_�i��of�yz�l_v��&�H���c������n��?+N��c�5�^����˵q����_��O�t(6Ya֔NP�2�����fLT�RO��uƸi�%�m��&r�'3�r��X5E�=�	�	(.���t <Ic1|�t�* \�Y�N�1ڔw����
K��X�;+Ӻ���i#sf
��6���I�_B�V�	.�w;�	 ���FړR'�C�H��`Ż� �2�t��s2S;iY�\3*��a!�q?5�p��Iz�ȣ������,�J�y��|GFȗfF�&�����f�Dkr��q{�u_���|�7�d��N�+l{��6��L���KV���R.hd��#�!��P}|趟/Z����6�9���(��+��}��kQp��+W����I��uHV~���¡8K�$�<��w�c�U���ФJ+I����p����C����E��� ?ky�̮����v�E���l���y��3~��L+���Jj�c_з��5,\		f�ʱ ]%a�Cz��?>t�O���/��K&0����͛:Q2A�)]�G�*��(	h).�.�������+��Y\]R�w0J��I
�ai%�3(���9�*:	��h9ܓg�Ch���&5����[��D��I�p������B.9)�� %��G�	������'ˬ�`�'bg�"�"�z��!�)��?������_�w�)�g!�\�;6����q��m֭^��i�Mb�E���^���]H^B�[�gg�+�;(���e6sA+����`J�4��DkC� �=VaF��f	=; 9���Ǔ�Ns
e7>9�FE.�/�7���[3_��`�&��R]�f��~,҅��O��#܌|Hz�������UW����D03	h�V�<�F��̚&��3�4�4;!���%S��x�*���}?������R��LM'23�8�s��F4�� ���t"�P�JYE�N���Jf�q��s�{���-�Ǝ�Ο��W�K�?��e�is�
�k����ƸxE;�"��u^	AT�)�ֱ�$�(�票�J��KK��� <�?�]io=	�c�Ia�?�:��f��rzd���;� �-���v��Z�����&��-����t���1���0q�_zr��2mnr�i������n�H��_FB=x�������C-��A��)�c\��a�$�fX��vz�H�:Px������_�8�$ѣ �#J�^�Ųۄ��b���z�`����H���W��p}�Z��� :hS��tMs��'.b8FF�{�2��W�J ��hEyeZ9�u��b��Y,Gy����g�̸T���-u��Z��y��H��7aQ�K�9_�WE������ܣv��] ދ#����0ԩO���6��w(E`r[&:�����tv���Y�m����wA�����4/�����pJ~�����%A���U^J!t�{���6AƼ5�,�Z�{��Qt��� ��Y�.���&��o�ٹ���*�XF����:C���qٿ��/%K�� ��8��"i+������%�B�M��$�/0��`a�885�k���+��߳�M��;�Q�b>��^�F�#aҞ�1G�J�M��!�ǳ���HA�����L����p�����=�Q9��L�E)2����Q�O�f�t�^��-ֳ�c���+!y{����e��Ң�ǥI�����&{�	�����L/����%&���:�SDa=�O!^6M@� �1�z�|"
�ml�b-A�bz��hk��D_��F*.����NV��`���$�?	1�8���+罐��l�TǞ�}��%q�æ�< �y�3���H�	��Y��k%�^�A��߮�Yd�u�<�V�)���W��>� ����'.�¹�|�U'WЦV	�wTr���s�:i���ۀgp�F�@��v��>�(�O�_,���;ӎ��v�
�f�`+�(H�п��^�Y�&�ΌD	$ӯ��x�z��+$O�DKv@� �H�����ѣ�1o��6A)���vZ���^,�U�e ����#��Nx"�i��I��2?��߂����i�8^����:G�	�W�@I�L�F#����ERt?
��`�$!譺�I�Ox�Q���_�y�r��� ����XAt<Lnl����6�a��V�*�5��v9?=L�6�'5NUl����Vإ�V͖�!L�x��9c![���66�y���iY�����TF9��x����8��ƏJ�����վS�5�ZQFfS��Ư"�Qư�w�9Z�j��{��ӗ&�"^r�� �6��w0V���y�gLYt,J���D�lu����
Zo�Q�,����^�N��:�kh�wT�s��R*��B�+zs���k.���fi�,ڀE>�I��h�\X�J��T��Z�R�8��V�O��;��9��B�Z���f�T��.a���*D���Ԁ̆�o�����w5徊	��8��e_6�1,3@7�P�^X��%�]/�����2�Y���q����5a�	��jx�Sg�o��o�,s�p�o*t觝\���M����5�Qm�0�������\=�7���Yx8��_�q��%���W����<�h�?��ΰ�|T(gp�c4�G��o�n�78@��gƖ��=4YIa�@h�����ɕވ�L�vð|��N75A��a�
� *�ّ�=�X�3j��*b�`�1w�Y��+ڠ?|dƿ����3��$�M����?�[e�Z�C@��2��I�(�i.��J�|0$��{]%^��Es�n��*��2�g�{=k�7![��{���!{GB���!����֗�W,\� o�ص0~���;������K�}=qL�pz|�&| �o�Ir���K-�u�c��m�6��P7q��WUVp�xє �3�q����풄�)J"?�Fj�a�[;$45#�V,F�E��j�a��eۉ*�+C<'m1�n��5?7�Uo#�r �!�&-`��Q\|<�ػ��H�R�k� Uta�:Fs7�}=����c���wʀ)�YT�%�n�g���K�F��/5��ӝ.�wZȪyQ�m2[�R�J�G����@bZ#:����v��4f/\"u�E�𸽼!��w^�r�7gO���]��c)�8ۖS�K�5K*��qڜ��\o�0$#=𬘁�7���;:�pf}l�=̏ˈ���g��2$e�:��MR(A�Ǣ(5�4$.��3�;��젫ơ����%�m�²E��tQjD��IJbL�)�~�|��YCg&S�0�'�=�ej=r�G4a
��Tڗ5]���|;2b>��!�8m�Xj��EC?�d�>��S~�!�
��ⓢ���۝|��5�z�Z-8hf5�T��ն�]M-���
���?�@�G�#��>#��e�C%$����.Mz���A�2��4ڎ&�_��f� kf�����n���B�(�ːS.�l-W�����K�۪�p@�裓���pyG�>Fm%���u}�B��v	��ۃ�U, J�yQ�T��Ԙ��r�c�tz�O��u3r:	������t�dȝ�d�ѿ!����N6*��;�0��s; <D�P]IS���x�fJ�7��`�L���5Pσ���]��U���db0@WCS��~��2K�h�l]��2ev���Q�Q��-�2�G>Zd����6B		,���"G^��Ր�m�'62�`M�L�7�IaK#�F&�[��~���R��"ȶR-���0=h�W�Km���a�����Xi��bF���e5���慤R��b�������+	$;C��GD��*����%��ob�K���k��I�Z��6��j�{>�� +e��Һg�ϻ���[v�3��X7�@�&����<k{[��v3�o���J'
����rx��� �a�55�I��BX4���2�ط[0�����6�̳�TC�~gd�׺�i����f��)V��o/��ę��9c�����AT���9t�5�������w�{Nzg#!�ؙ?�N�֪ς�^T�s8����
1E-z�l����R�|��ғs}"�P���Qm�`��1[D��'MOH��sQ���?���b��w�"E�%e	�{�[/(�R���а"���^�ox�ʿ�����-�?Q�va�\(�'��6Q1��K��f��f���3�T���/�C;5��I<�^��>j]dX;Ο�/D�s�[2��m����B���Heq ��D�P�%����6R�����Կw{A�^z�����D��#�ekC�"��c���N� ~�E����}&�KP ����҉�6��+���l"��I��-��Ď��NR� M��b�	�N�H����C�K<�]��_�D�f��qT�n��1��~H������R˖����/�9o[a��;��U��7����q������el��sƼ��
'�w'�-��iuע�"=����؟�[�?�!}�f���-�6+�}��~��3��zo�Ih��/
R���8�FaKma�w�]����\�y1�H1K�TBOd��D;t�=��<is�B����y�'�˘yN��fc�(2�����Jo�~��R�C�����2kM�kwNE��W���/���(vo��.f�X4�{�H�n�s/�/��h��-[�Ɵ�[���'��sk/���[��sc�{,c�Y|���������?�@]�/���:`�Z<[X(��mtM�9o���\���Qw볕��qo|���p.'���ࣖk����W�x껆��&p˄���p^�2��e~Ao|Ek�#p�W�s���ꐮ��"I�;�w����fS'�ou)�����!�R2�(|0
Gt��8�i�l(��q�����
��9�Sf���-��#v����e�@h���Ղn��ְ4���G	�٤s�=�"�D�1�����iF��O�z�	.A-�Ybm�yuzu&|��;���)���x~�5\W��d��!I8n�\�"Rsā?��-?�J���q^�ڍC�0����=e\�л���I>�Q7�������YG�T���s�ƶݤ	xD=��}_�C�[����H��K(P���U��$�����1jf���F9���F��N(ڒ����làk��F�T��`���_�'��Tpv8��WEقh���h֐E��AK�׌0���=��\f�2�Z�C�2�N�KS7U���[2����׼
�v��	�w���R3ef_,�:�D^N9x<%��vЄB�h\V�ۂ��z��k_�;�61�6]�	>P������\~�"�I�j��	�=��&>ڂI��U�����|�H�?m� �U8W�c��+��$���hT`�k{D	�3t�cr��$�glZ�l}��]�
���Ȣ7��=W���];�o���[mRK��T�'��ņ�!o_�,
\���[��J���[9^�=fs�0pz�ȶ��� ������/�*�<:H�04�c��bw��U�*��A9^��e�C��]r�2������O_}9y��vw�
S������C�U�7���9��=B��sZ�e�ȧ"���Zۦ��/�/sVTB��MK���B�5�IN�I���l���N�Cp��`K6�_�O�Cvv�_�}B���1ӫ�%r�P��E�P�P�'��=�� �5�Tܿ���PMKvb)�.80�����W�>P��n�����Gz}Jvv�*A"�|���qq��>�Uf���=�s+e��kݥ���[,�:���`&��'[��H��P��膨��&��z�@��1�3����U��(�Zk[�#&�,䧸b������[e	p�b_���?_�~p�]h� ���w���vW��X��fE&2,6�W5�ǵ�k��7������-@Ķ�R��T�J@2�2��/��J���4�I[[�����)����D��� o0"P,�����D�b�\�"��t�q*�^�9	���`��z_�=��[��K��tA@�/]�`+k���-�����L�'�j��=�޹�̰�>����ܤ��}�7&F�b�ح��Y�Ȉ
�F�YdW�����~��`��m�lq�Z���*����B���~�_w����߁n� t<��\���]�a#�.���R�B��}]k���L4�m��t�����	���__9��~� �B��ed]�'{�ۘ�a`&I$a��YZƙ���W�6�����x�]�:��j36����a�4��[�g-������ao�5��E���#�%��
-`�?������֗�3���
,bZ��.3!��	H��)�4Z/>pܹ/�P��Ȅ7�8�ª�l���5$�Lt̅��񰙺m͙�|X;�ȷ7��y_�^K�9f�Pc
�t
��c��S�+ɮ�ߪH���<1�s��9(���Ƚ�T�4��DYtW�n�i�u�W~�Ҷ��w�$<�K�,u��}Qj<D5���~�*M�������6^jې�DlVT��)��[R�3�/N`)�PN0�UM���[��$�+����8��~Y�2k���'Q�c�ʵ�y���N���7�z~�4B�ߍ�N$�$��dD�5�Yp�?��H�?��!5s�bU�O���i�|��X�Vs��8�Ny�{���tna�7��0
	���6�^��U�$K+�9ߓ�Fq�)漼WX)_��8Ͱ�P����:�jQ���㒤n���:.�,g7�#OjT�ʘ�7�=�:L��P����	J���w�`��7��;h[h�� aK+���h��<��J�Q�j�Xf����]_V1B'���q�-�ț�pL�@9&!߯�w�u��X}�$eǽ���91�w*W)(?��{)7Eؽ�޳�����d ��]�=@W*lG��G-q�t]d����J���F�;`w���Ƙ�`�O@���F�a��73D6C
?Q�e�]Xr�lc�V�ψ<��7��P�C,N��:�!��}T���$S���$��-	��NyC�n��R[Op��K?����ZI0Bp�buA��Z�|P����e�]�~�1�	�)��ظ���p��%֏/GU�]�Y��"%@�	�q��7V�
� L�)i���ģ���c����˞{U)�գ���3��v�J����O���f��m,y�\gBG�g�8��9P�xE'�l�ƭ���Su�=���v�����?�ȗ�nnW3_*&N	GBH��Ìc���w������_�t��o����aC�2#]�o�I��-�&
Խ�ns4���ѱH��F�gGɒ�`P~��	#߼]5��`/	(�@�¡���	o)u�i\�z���$}-��0����������Š�v�LV�)N\�wt�W����,�p���V`�����׳Qp�8�H��dfx��*N?W�p>��,8}� [_�������6%�^���2O�Ke�2��,�枸u���Y5QJf�ng8GL�EBz�jy3�r^����*��\r��W�(���#Ák��K9Ӓ�0�1���dL���ĸ�q�^.��Yr���X���a
� <A������CRP�9�1�q>�f2\+]u��!?5dտK1hx־����ŷ�Q�M7�^`�ĥ�7E^�ٹ��QGvѧ��;f*���+X,����`�W`��Q��j� rQ���4����Tw��b�!�,堶�rw�B�=�#,8v�+��K�Қt)n�Eʤ7Y-����0�T��?.t9�z�43�~�(�fnE�ґ@��e#�C�8 S�X��5%������aQ��P*H�����|Hw��E�r����ҥ9q��̰�/t�޵�]�������#���r�$o��S�t�,���A�{mD&]�C`rA�~����"� �R�r�B�{�g?,�͚yz�2���$FlK�J�;���	�&�ph�O��g��>nڼ��N$��Û�jح��8�ˈ���$��Pn��lc4��"/9f��)�%_U�<���T`�����wʍC;b'G:�XYu����>�xc&�"������Z#jOº��;kd�ٛ.H�h%Q�U!;�4߻A���N���;}�;<>^�Rw0�S6&��uN�Z{�F)2u�dL��@��y=�?�YB_���?�4M���w�E~Vx��Y�0v�4k��b�S��u4�]$,52���� �l�!|���Gn�R����=#Ew�<���~��T�HJ�e�� ��\h��,������Ƈ24�9�t���v�}�6�XW�y{3"W�ë�����rl�;r���^�wҊ�IG��Z���Sw���Cq}�`2�$�Z*��v%�H���H{PS�w.��\�( �܄��Q"1�@�K��	g�n�;B�n�9ܕ�L����I#��}	��y<�9�b���-3�d�����j�3_>qd��������08�USI.W6�4��(R)���=�o�L�0_�X��� ��� l��ktb�:mWW����$�NW��[��w�7C�HuaK]�i��@�����^�⾱��;�� �sc�Q��jC�cs�j��c�W������AhG�b�ɼ��4����g�D�g���U�<�i�۽ʉeY4���H�h����ލ ņ�u��,-E�B���/]2l�~���nN�Y��حة2��~��cx��i䳱�!�Q[8��DlM�^�Ŭ��	��$�+�ea*�^�`K&�(tѾ����yh�eHF�-�����xK��O��ˆ"A�ġ��}~BG���=�dg*R�*��ćdhڭ�8KK��5�yp�#uh���<���u��P(�ΚȾW*Tb{�7+��Ѷ?[FyQe��%��<�`�R�UɅ�s�!c;OQ��ni���>)C����c�<ژ�{M��mj`�<,=�L��eB����]�E)i��I~W������|"�ٲ��	�u�Tc���}���$#/6v�a����|�`/>�3�7�J��V�����J+Z �?�3�Ő��"pE��{`� E�6u,�¤�G�1���嬣��d��TRű�9\�(����c�W�9�l0zxE�L�Vَ�����,�AȧtD�>��
cTx��v��"�>@h�c�R��B�ɠq:��G�_k�~����Zm?��Ԅd��x3�Υ3��?(Q��^p� X�3�h������s�j¤�~i'F�bDb����6�#�Կ�� #��˼R���UdW"��!g}����~HS��]~0n�Ģ�h�����d�#[d�@:�8�R���hhE�1�i�i���u��4��D�G�Ly{��V,ù�Atڣ�G9L��_��*�ԅƺ>�8�m���d�o'W�k��-���>�}�ʜ?��z���毫x9��,AF/�^��̡��od�*��b4s�lԳ7z���,O5�;X�E����[��XF@�lkN0O�n�2�y�pP$Ɲ�__�%|X]p���e��s:��r�}�)(�%�9�����K�7y"i�q_�s�_k��l���B�	�t����x[ϻ�(t�l.䶖şF�%�{=�X@��j��ٓ�X�N��2yV1�y�b⎼~U�&Ί���k���Ǥ�yN}�����e�9�D��e_'ɜ�Z�9	��~kJU�e�A��6��GN�^n_����l�����@��T�ֵ�?�T)8q��1�陽��>�1u��g��b�r������[����uʃ�>���ܲXl���������)�+���Ǒ]����&�#Vμ���2�����h�c����� ��f���~5�O�-M�������O�Ĕ��_F9�E8|�qL)"�C��8�����.4k���&zz�5�����}ѱ��ܣ�^����kQ�؍ǥ+���G�d���D���V$!������
yOI�u%�BhbՑv���B�JH��HZ������0�-���%�� %)�nR�k����!W��ד�l[���a��X�6v=V�ua�A��`7���������c�Ū�3���_��G�>�ͧZi�l��p~"A�	���P3h�����yc��/��Q���������
�x� �!;�׷]����A��&���*��������f\ӹ��iQF-�|����Փǭq�:�B助�C�[��]��u����E֤<"�j���t�-5�L�Y�;$�i���|�U*)a߬o����M�8���9(���R4�O��d��e_�ubf��1�1"l��� aM��[�	�K�H�{f���37K�lXf�� �*%O�&���k����-���e��� �7�h��>�p$��o�C����O6�>���o���%N5
qZ��J�/�	/�f|��O�1�9?3"��&A�s�@��_��ٖ�^��!�q�m5���c��Y�G��c_1���q��A�fN���!f�S����Z$��u��F��v<�%�@FF�T�e#���@f�V�.d(�F$d�Y�^��ɱ��9��,a0|����8�V�՞�D�Q�[�������Q]��8O�ƒo���N�����a�%b\�z3��̔��B$��Ꝧ�d�XL�W��,�ޏX�����kgڰ�4�w܏9���F�ƕ�b�)�K���MH�Y=�w�i��җ�߭c�{A�T��Ls�)Yk(e����0�*8BMD)��ϊ��
E�@��S^��
߉X@�(�N��bFii۱(H7�Ƚb�r���+�<f��Ot���}Bng��wN`'Kxu��E�~�xZ�]T$�ɩ[I*%���
��[m�(�:B�ޡ�?�C ��5EY�c�y��5(���/?b;J�
�Ж,M�#v4��r�,�4���n��8�3�Zi�M�"B'�'Рsk;�Qw�r���d5�N�p���59r�>X��ﺐ���X����(�/nb�c��$c�Oȅ�ӑ;z�����w�����@�M��ld"z�;�
�u�]*�l�;���|�P�s��;Z#pi��n�$;�k{��#qq�¿�.�0�+3#ע��i4��L��_K�yi�����ai�v�m6�l�����#gxό'X��w8�4��0R�w����+�n��4:.(���"9�!h�^ƆE5����K �(�2W���f\C�%����g�� MJb�R��k뀂�haX��U���Q�q��-I.�ӳ�Y�.7�)�7�G�n^!�!�4F��QK�����s��o�ΰXg�H~T��炎�R�ُ� ~8�Ӣ7Zkt4]�hC�D�2��Pg5E)so!��-S9�n4�-MR�=�f�rJ��ı��*������5.�W��?W�Y��"���-�JR���� ,��]������v2i�u0�MU4o7YM��χ���Ѽ4�f�2%ء��OR���
O-`� k����NB� ���$jZ���sWNP��$��ފ�ҕ���5�*7���m�T��ӫ��R�z$l����7a��#"�X;RU�����1�R�t�CX�_����3����I�}N>��#f����Eb�Y;v�"�,.<H0��(��/�р�g�݀��	J' ��X�%�r��}��Gc*�DN�N��x��5�b|��	��e�.N� �P+���_DR��v]<�,�K^|��?43�:���4%O��ؔ:�
���gO>;P��,�׮s ����i6�l�#SZ�ݽ�l\Ƅgܿ�[�Э	ܭ�un�4�:���%.̄�@��&h��Cw�n�p�&���
�XC3`�5��8�&x@���}�t� ��πaR@h�IY��8��8@vЁ�� �ى\D��Ъ�#����k�$;��q�Wh�k����.'ε�sֽ	�E�0hJL i�Y6'�E:(����?_���|�/���s=�>�}_��_�+L��ZXFH-&�͘y��!�Dc|�W�ޙ���N��z�=I�2���K�h8��5�gr�K�!��q���W&0�^�0n����{��u�%a���Gx��ү���~�ƲC�Y���S]�q�S��(
�s�L8��S�C�傞����I��!4ۭ�d�y2���%��Ԡ�v»����/{�y(^��?"<UN�4�~�gHvy�j�z[.0�Y|��R�\�α��x�K�W�7�#QJ�yFfM���HN����X!�a����1<�Gp���T�L.!��Հ�*t����Jq��]�*ٹ��C��G��=��ΰ���T!���<��*���V,(FN?y�-F�5N��^�G�ׅ&kC�KD+��wS��u��,iq�Wj1�4�b�h[\�T�)<���^vl��8b�l���S���Q\.�Wf��=G���yVZ�:>B3�*s�潀��-�$#<MJ�6ҋ��y��ww��A���QZ�u詆�:
6]��-��tz��?���ϙ���WtX툯��Y剗e��3�V�Ox�J�h��E�"�<,�iYK��Gy�e��K�\^*#�_A��/4�&�1�Mc;����I�f�ؿF�+s�	(���i�"4�Ï����*9�į�Ζ���<��Z�2l3�g~�}�	�노ፔ|����F*�����F��c���Ěʨ�]vED��J��ٝ�R^�����i�ݪ.�jq� @`�/������V�:�@&��f��Q�B��+��(]��'��H]���_�����1����L��v�*z�\�,/�� n1KH^����ܾY}��^�����Ԯ���%M1��@�5�	��DC"��C%�� #�w!�p��KʒH]�����ۦ x �j��<hi,*�7ӗ�/��@��܂#�4d����q?i�uRj3�Uߴ�
�f�L�*��#�1s{�Ӝ��������y����
'�D���[a��L!6�8�����چ���	r���:�ee�qx2�b����kH���U�^a倌��mK�u�m������H���e��L���(_�+p�
:�s5�ۍ7�W֫���M���� �c�>M����{s����.9��S����r.�Sk���Tw-�,)@*6 
Yח�������jp�7�-Nb�M�fP�d�d�Ւ#���!(1��?�\�?L勉�&=O��P��b8v�&�t/!n2�T�*Gٚ�Y�I��3d��u�S���.�۲$�6RD�>����R���߹:�����aȎ�~�r
K6m�׻a�6ɹ@�Ԥ$�*��ͦ%��P>c�a�S�=���{W���h��$���f�O�-�V���������hx�)L&uT ��{s���yq�w����;�>8է��}-�v����T�*����E1Q\y~d�f���|r!bK�]oƗiod��{��]���N?es�,=���#U]��� �2��:Z��s��h���`�D���P�dxk���.��n�3'Nom�"Ý�!����v��>���qO�Ph��I����"
1��L
�+�{ �r.�ߢWz\0'5{����w�ܨJ�I	��<�x�a���6��:B��*Զ��>A)�����~1�"��S]lm����b�r��a�ͥ�F�O,p��OC���m�")g�W5���U�M��-��^X�e���yğb��_������D��=lm}��~(����L���Q3�q�B���Ol%0�+�)c�u���+a��ھO=����#����`��e�����ǟ~�����g��KU��:CTV3������X�4�h�Q�^�>�K�1(̏�b���0��u��|�0�aC��Q�� ��Xh��ӭ�K��w S�V��
_�j�ۯ����J��og2Pm��Y��?4 7;�G!"�d�y�r^T�}i��Li6 J�(����\!�]̴����a�F� ��Q���G^*>��է��at�w���h�>e�X�����t���:v�K
Xm8�|	U5Kn	I�^Q�{�6Ο���P����b���Q��N�,BBAa])ؔ i�8X���$���O��h��q)WP|vv��������"�˹�����3�˺� r���?6ﾊ��M�IZ]��rx���K�j�Q3��-��VC����ǭ~DE���lw�Ui��ҷ =,Z/,W���J"4c.�+�i�о��Fk��gM-�C��z�ȹ�F����E$ǆ���'��To�"�*Os�ƴ��Z�GX��N�m67�fPS΂�%�3��ak�I/�=l�Ѧ?&s	�gλ��n}�,3إ)�B���t�AMeu�B4�w�,$qW��?��rj�y��+5��q�Q/���g<ۼU�]՚B����oŅEK,�P%���⣽�5�6q(h��]A�*W��}�S�O�5'���[�5�@x|�>qo�Uc�J�m�YMA���LÏ�7�b�Ǝ�1䚾۔��"��M�!E�z瓷|;�V�������$�?,ؘ&�%"P���B�B���|kc$�NA�[i�,�lЉ�m�h�q�l;��.�s�ƢO�l�M�H��T��xJ%2��x���ד<#r�=��^��^?�p�����[�ex���ܪ�n;_�jM���@S�|��朳(���Y�b�����aZ��^͔���ڣ}�6NY�m�#N߈��>)�|��Q"�ޮ��%%�u f9�3�ltホ��Es��
�x�vϟ��FH�^ci��D��|}����wc�X��^�ͷ�e��	V��g�)�$��P��u�ȗ��,h�l�Y{@����[�\�cR����j��Y;���0�vҐ����C_��3��I�[��N,���h�:|e�4�x �xt�u�����O��_&�]8~�EP9�g�c�{���V�3�k�#0d�A���zť �i��H
b\4F��+�i�+���^v����)��4��F���f�UCXb�̢��l�OДQ٣�T՗�52�s����&�W�E�'h�������W.����%i�n[���V�]�>2G5�����+�e�ic���:�?�a�t��pއPV�0�����'f���(�b�L1�W_��.�W-�n�٭=�XX�k4I(gAG�C���T�xԒ�B�ܟ�F0�Wx�۸����ܬ���Лէy�A,xv��6�����Ƈ�k���:QR�[�UqD�҂#J���~v��Λ�� �w��R7k�������G3- �����m�����
��tw��Ϲ���2�Šk<�j؃��F����UXr�D��v�����ꔕ�j
���#j����4~-c���M���#�������O�S��;$��ǥ��p�N�%o���C
�n���\�,/�*3�7Az�Q�ɟa����<�
+ӂC5O/孰�evo<>6�eY�'E�mr�(�i�jy��-?+�O*�4d�dC�z|�T���~��V�֤��uӜc��L3έ˿ҟ��)kd	Qe�S���s3�v�/����s!�dk"�LS�䞫��W�o�I͠>��֩"o$�0s�I�~&���X�C}	��*('z�Z�#t;{���G�q��]n_���mP�F�����킘���s�}�� L�ǦDw|����몢��"��#���W�M.m��Z����9s7w��z���ܻ�ERR��o ��T}_@��%�������yv�, �ט��<Z��+q��n:.}��A���F#˫/�-����_ˎ�8ɺ-ްAb:��xs��P�F��k٩�E+7_�e_�=F�3r��p�%e9�������'�O���L>K�B�2��~�6�=��Ÿ�K�JΛ�b�|��ʧ�e��h���u�F���_ ����s!:��Q������"]�	�}���`�*g
� m���KRGv~%xK �HژM}���ܽ'�?*�M��*�q����p��5�p�9����&A(��̜�<2:z��8E&H�1$ ��Oפ �����\��)��� Ρ..;���-�\��%��y��+щ]�x@�&8Nc�МhnȚ��ɐ0g+��p�c���J=3�\�%n��cmq*!��
�}�C�V�]��˓�A��x?c�E\#Ag�,6���0&����s���W{�˞���P	r��py �x��$Is����y��CK���}�{���t�_�7D�CH�Q`�S�9:� �w�n'kf�)tf���H\o�uL;K_�	^�CQ
��4�at���AQ���|�olm��� \%�+��;��Y�Ѭ��L�R��_{�hn��m>��gƼ/^v=_bC4���a<w~保?ND���6P��Q��:lĐ�V~��(M�Gm@~�᎐�l������`�w�2�SB�e�u�{�L�a��!ώ��9���
L('m�;�Ö��tHŏ4����8�
���O?�c���T�{v��v���~�nճ�?�	|�kV�l�<�"��`Mf���@E���J�L�N�B���o4�mT������� \�0�c��ДkoD�l�b���A{)7to.��;�f�	�:%�L���.���U���3[�^Z���40���QHF�b
bk���[������h���cC\�u�y�i�_��loV-�v��U�ĕsd���k��b�ot
��2�<.�GI�X�D�����M�s�!x�(���tՆ7;���׊e1�g�_��xMt���<B��Q��DoP�.��k.&�;��)"�{�Ʈӟ��6�u��&���Zg�&�;�5�M�X(�>h܁%������"����f������1!�1����t!�6�VQ�D$����B�O�?��O��^9ڏ��q^HeY[ ���\��+#ig-`��>���g��>>7�BX'�7��_����wRt� �fT�ZBj�9������BU���bR�;r�>��\c���`�Ё��~l��︁$ �kW��_��L!��	�>
��ٞtx"�z�~z�|�,^�AS
Q<3c�}�d8��g ��H|z�&ȓ���գ<��>�X�Tvx��)Xl�pd$ �s����^�2� �E���&�q%F�Z�m��D��E~m�B����4�߿�m��5��m �3� -z�����-wT͝��d��L���� /���.��V����3~\���1�z.��.�f2�k����}��D��S6� ��.�Z�	o��$2 T�*�*�%�-��40R<Ȅ_�øpJ�^wsy�C�����Y�^V����k"LR�Z]A���@�~1��8"t�X �0I�{��}]���NH�)s���1�ȼs����״R����&��H�kFo�Q6S�"�ڲ����	���D�����MV}KY9IiL:�M�K4$��@��O�lt�eۯ!0TV�����UK��afdX:�HPUy�9wo������:��S����_�!R�rY��=[eA��^:e@{º��_+ʙ	�Pϙ���!]�+}V��r]��eR�e�Is�E�p���Ggj۰��5�ry���[�Q�2�J �*��^���䒫E�j�h;jm�� �)	���IRÙ)��|erYL�Q���Ҍ���cj퇒a��
����,Y�-��j���C�:��1���F���5�>���Y�ZL�֠��P�JK<SC-'â����»-��Ie�(W1�t�ֆ`����h��We7>/��M���`�匔��{t�C��/�ǦY�>�� �`t��Ow�M)~�5J���&PL�Iu��C+�)�Ĕ����,ˡE��d����r�0��5���N�a�2��8�H�����E�M�&�ra7�y��Ηo�;���s����0���ك67@��3S�J���Y�-l��n�U4�')�J���9�+<���`���!CJ��I��)�l��Ȫ*�t�F�"tEe$y����1��g��R���֙�@H<"��Z����A�	��w�͝_�Bu��"_S��/��Q���|߃���G�kT���Ȥ�R�4t��ns�����'����<��</�[���㖑gb�[ӂ2�-D�g�L(�`V4�4T^)4�~7�B�1�t=Nx�qv�J���0�o�X��^����5��yX���I!�PO�B�K+�<�Z.�3�6�����HM� �+o>*�*�:҄>.XP+P����Vu�ڧ>맄�cWF�~���)W�aC;��Hٽ��i�u|Y�A�>3{� bj6v^�������~g�t��תu�GH�!��Mo�q:���_�{iq�NI;�V
K��
���~��^�(���K�����.擛?����:C1��
������pĕ�)���� ��W>�iR�rF�D�z
~Z���"E��kFh�Ћ��Q`�~ٲ7��bE��r�{/IS<�( �r��jK>��U7N�;�'v����~�Z�1bM��'/�/T�S�Z�Asr`י���K�����Z���Ǖ�8ZE��B��������[$��	߈ W��4�ʱ�R�|��^<ZC�V���=�Y��p���R]#^䲔��*<Ã�6]F�6�������9j9�FLpb�H{�&�@��9���x�BǙ$���v6T֏�]̖0��������R��-1�lD��PIM����C¢pk�y���w�1RgM�;��<g�4js��06��T!�z߹:�RX�m�<M�R�ۛ�
 1Ǒ"g�>�fx��FB}0��l�{���&s �6x;f�x#'�ߙ�B��#hA�]oyg�Ck�|$�@נ����OSW�@�`j�Ϗo2�_�k%���$���2�c�m5:�>V��GQ��" +�/���j�V�)�Yxk�(
��AN�?
���5~�x_�m�1���[��������@I/��G}�\��>��GBPy�a4���%Ip�h�o!�A�4����|Z��Wk�c�O85E�f���A����sM���=�.��������}�Y�j��2��U�s�ARfO4�?E��ެ����G��M;2�'�����q,'](D��EpX�w���[/�C�6jER
 �E�Y�I�~���P\'8�H������dИ��^��t0}A���L�T�'r �=�h����N�lA*�*�`7zyo]�B�5���c.߻����R�^�p���<o�3�9���=�Y7{.̼�E:������}��B�#��B}��,�}��n��AR&6YukH]#?ӳ=�q(|�^5�MF�_h2p�'�)U0�/-ïv?�(���*����m���B�#�j}�<��`�r����4��_� kmQ�����M�pe�����34���rG���Fw>b1l�?�ȳ��O����ŉH=�'9������&�a=��=��z_A�����H��H�0�P��Q�5E�kq;�]�㸢�E�Q@#W,؊�k�Ӱ9�L�_����᫔x�g���;7D�^m'TJT�����ڂ�B�0z�M��T��?/�w���eVS�Zu�4��&��M\Z�}�������\��9�P�08%$a�j`�Ǎ�'3�x�H��ܯ��-�LDæ4Sl������bֈ;�ri-$nݸ"�˗�w��;K��I��3�2+��݃���r殮�'�Q����&��l5��kQ�khK�b{�ҝb�T�� �dA��.v�7�*���f}�LỀ΄���@`�.�������{ �L\�`���i���.QҠھ��~v��j�^h��ֱ�����_�>`��;�Ѷ�p�l���� �43e�x�%��^��@te'�T�m���x^V���s�m<઀�>J`�,'|���V9B�ʯ���� '�����;_��m*ڤ���w���o5#�����aMOи�1��G(��
!#?0�>Lfs����s�wFܕ�WbF�0,�y���|h.�J< �fL�:��ϭ}r�/�͹��%_b���m<��e!@ ?����H[*�O�%S�En�{�Z�P�!�x.����U�DDf�!cQ���#hR�|��iU��3{(�㪟*�
p�Q��'�3�e̩jp,�ClH��a!����g������΋X�r]�[�V++��y�8��g��(�}��2]���SE�]s����h���/mg�P�%�5��9��v���p�>5�R��,3�J�_*���5��Zg���lF����|	ۋ��o��\�[���V�n�3l8�j��SÀrh����1��'�%	���.�:��T4��.ق,���%�8�����X���Ѻc�h�b������Ԑ�����#l,gP\s��o������ޘ��k�vkjiҟ����P�%X�pϚzm3�2t]���@,��J�tO�M��eU^����>aKT�6y}bR0�4��Kɿ����q�MJ��]��7�"��Op�o����3t*C�cB�P�����"�G����Vt�Zgk)�ȿL�T�ζ���܁?�s�]�tpq����8�8���/��`�i�Q�(v�iIQ.Tw)����R;�A�:�(����IY��?��������ɺ�.����3�06	�#r���M�(
�l�W��p킙Q����Sm�$q`(��OA��m�`��� i�Q�+�Cs_0����e/-57�����\��$ќ'�j�������M"A�2Q-���E^9�3b�B"q����kxy��w���f��f��3�֯u�x��jd��3����z��SI3Z0��V�g� ������W�ʻ��8�W��j�t�6C�L1���Ї�6�SD�b��]�9�ހ�A'v����MX^B%-�L�Pi�>�׍��ӆ�N����7G�MJ�'��jTV7&7?�
z�!��f�j�%T���S��)���h\�s���QQޚe��� �	��%Vn�d�-�.^7i2�� G^�|�YMdo���1�Av���o��03��S���^	FѬ2�[9�)���6��cj.��o,pC-�pF�2Z�+�
[��@A%�8�ݿ�v�v0���p�6�G"M�E�O�v��Y��S�0k�S�&!ĝ8s�X0�Q��w%�μ~e��� F���.��7���V?أV��H��*��Ug�*,�~��\�v́"�2��E�x,}�����Q5S,R�W�)%W��PdC2樻j&��],}�5��q�&�Q�s��KSɝ���4ȗl��5u�0�������k��ߓʛ��71Z��eJl�]�o���c����r�_�I9��^�8b/��##�o��͉W_j ���A���u�^Zf�{�ľ�Nܻ������)i20�V��3VjD�G+9
\^�E2`��h��L��5=�¯��R��n�$���̲A��&�l)�b�?Z���}k�7����w�tVM��1��K��6��xے�E�?0���K+�CQ�8k���(��"l�һ���^�������/��|����(߇n�|3|�s"�O<��jHi���̒����	��H���7ԕ����mF�?A�
�Ż���7w�1���3��&wA��V@K�`q�����_��˿�L�;/�N�Ѽ|�Aa,=����WaEsc.M�f��J�P1`;\��;/pb����X�q�o�PO�=:�@^E��B3T�f�cͭ�1a��B$jan�8���&�(	�{#�V�*#����Mи��	���tI�B8(ʱ���1 ����$Z�k�cA����O�D��#TS���bN����Z�0�<a��<u�$�Q��u���R0��v
k�b�ZQ�.�d����<�T[�6������A}����������"%*Ӣ!Տ*)�!�+�����m:�'��I�s�b��!ŗ��W��N3�\�6��qM�=-���8�,������������JR!^�A.��Dz���
ZrK΂q(-3����4��x�� 1#�b���L���b�ѧJә>]��ȯ<��-�5���-R��ݪ�%�-0�h��^�$���敮ǲ����U��6�G4�V�я�|����~�1(Ԑ
sa~��ɉ�.�+K8Ix���6�
��ݺJ1T�*�8&X��>��5({���*��6QU.Yq�t6_zxMԝ�z+Q��>�GW+�B�B߂i������܎^>Z��*���a!?�"�W�e����O�6=��ѕ}9rց���?�-�X�^;���.��t�V3p ��e�L�����:�'���|6��Ө����ҕ�s�8}�+2���Z^��Bw6��s6�D,�dC��NN��8c�]&�jb$�2cnR�?_��;�?T�ej�Tbf���(�� g�7�#܏�=(�G�9/B��4����HzRwǩh#~Iڵ���;b�;����k>�]�*�������Bt� �����a��4��p���gX=~�
�M�',Ih�Ü�$�� ��`���րހC%l����#�(��覅��o�rOq6%��pi�������W�Ȱ��QA�-1�����'�^�����{��������4�{�K��/����4�����@��  ��
�ͺٟ��W�)�%S�8��p̣%�<b����*�r5�' *��9 z �k�f�i*c�#��r�Z���_r��.wwv��P�`X �=���6Q�uQ��z�������S���GCu��_#A���7Ğ[Z�+��m�VL�Y.@<J�2��4\�R��s*�]�,�rlI"�
�^���C�3H�x��Ou��}��B]�x��z�������%��O.�<�P�Qű4��G{�u ��.|Mv�8<�jHh�5���W�ᛯn�+�TF]Y��:v�5�C����v#?�2%L�/�y[�B�m^!}G���c��T����/v�$zl��)2l`��K<|\�L�Qx�R�6l���T��<��r�y���N.~�Y�+� ��!�����r�[
*R��t�O؎�n�����K�9}JL��d|R}^E��6���1j����c�h�]�iY~���#�'����\� 1gfsX����k�8�Q��"�����[������-Z+�!����d�z࡟�@��L,��ⵇq[�=��L �˝���a\������t�ނ��Oe��:
��	V_��$#��f�Hե����6�*�}��{�(� ��\ٿHF [޶� ^/6eF�[녶;t���r���Z����
�>Sٗ�`p`?�ko�_�k��U BF���ӬD��Z�ycD�O����]@��w�c��M�p��7/� ��xA-�	a����0�P��M�I���g�n�+yB�۔�a9B�;
S�no�"_o:Gx�w�?h�������>���諫���\��a����Su�%E�jҁd4�Z�i�b��\k�xR������6Lq/$PQ��97#��=�3n��J��!V���VK<�L׳��V�ѩϐ�j7�S�%܀���_��s���IG\�e��I�u��B�(�a��/nM@9Ut���y��U<k�=������h�eyf<��IJfF���:��Nxie#�6�_-�Kw���ˌz������whM$a
^�0��4,�m�W�"b�ir/<�#�2uV��g};2�6����֫���$����)1|T�/fa�ё@3:<�H@��P`��>�A8Q�_����	tJ�,�Vn�����+7T���%���5d�^���#�mT{k|���Ԛ �����{;�$K����K�5�)�*��Q~ H�A9/UP$�� ��>��@���+[�:ԡځg �o	��a�g��/%�}��o<}`�M5�F�ؽ�����g�K��]}7��3�d��M&�h���$B<��/ݶfS��-N�ͬ�$�
妡�Y�����ƒ�ȕ�3-e����
���M<ڹ0�җ�.+ln�vxC�CոG8���X��q���JT��6��?(:�<q�X�K���<2�F�����a�EPjfxRpP~7Ǖ�vX��#�`hH���X�V�9�@0,�ҫp�s(�ھ����E<%��U㐜o݉�
�[^��)Hu\��;o'Y�-��L�+�_Dұ7���C�΁��M��+G[�G��. Pȴ��N2�|��a�=\ѿ��20������P�N�Rb��\�W'�?yX&I�ϭ�z�ә�
:�����uH6��)���W �ON���\��< ��b����S!��6�b�����%���c-�M�a����͓l��4ݢ�O)�����৘	�j�?� Ȓ@���E:���T~����o:O���X��ujn��U���&2J���?M���L��Z��w��isV�1��T���w��N�Z������.�#c��G��G�ڣ]}�Hi�`8�V�I����q�?J�V!�ɡ���������a.&>+`?�֟ ��oz��F�*�Ւ������UV8��(�=��W���i��ѹ��v�=����'�ڕ3����������hs	�̩����h��g�MLt�H��dxS;�P�����j��:R̘�m y~R=�hZ7�� �A�4vc�LkJ;��k�n����j��z�H�Ȉ6y욉ښ:7	�'P�%�͗�p��`�"��6Ϯ�a���6�T�%���7���
�X��K�7�� 6�UX�?��;��U7���φ���&��<��v�t���'ة����i�e��qҴ#�%��j5"'�4�ݞ���m�t�����w�P�&
L�z��X��j�-�%a|�~o�殌�0������k8j`�u���Q�Y��(��-��ypDQ�25�� >U�i%����)V�: W?3Z;�����^�9�Ox��+����y���*�j�|R[f�S?t��s����&c�$��`�� �!Қ(�J[`/��H�D�ireym�ǋ`}͓꾧���)���+,<`��
̡�T�O�x	�?/
�ȋ(K5��ĺo�E��*"��ģ-pp^��fP�̉Qazb)���";|+Z�L�NY�u�2c*$2.�8o1��I�him����<^�u��	݊ER�)3��g�EMG�S�D�~�I��մ����� ����{��#��q�`�o���q�����%�,b�(L�l�Å'�\O'.tj�̀��&�,�'�۱|ݦh�^�SccgX���}�ϗ�8'o�,�$׋�C۫'�r\��j(b�*��0��g<��o�Iy�n���x�Uj�Mh���5�E�p8�hz'V����èF�[��	� ���
y&� �/�|�*$}�~C��(�Xu�AZ��V�C@������=��چ�3�ȽiC��ik�}�h2C��Щ���p�8�V�Dx�p�KC�����+��h���P��>�)�����\Ԫ���T�:҅5.��	B�7j�S�ˇ�'6Z�A���"(,��71>��f��#�0G;�ɟ9�c����Ym[�I��A��s�⮫�
��$;S�����!���U:YlΠ)Q��3blb
nY�^�ލ�~��=i�,��jv�,+ԣ��vU�G��jP���v��X��A�1ίjN[;X!7�N:c
O�@����A���;K���ق��Y�%,u˯̓���n��90.��㿅x�*�C�c@��wm-N	J�N��F��h���[`|"䔪>H�Y,Z�K����`O�[���*�O�]���r;��8�3+Ǭ'ձy�=],�V>ߐ��!!ğ���
Pj�$Y�B�H�^��.�Me2�1��-���N��n]8���EM�g�ZB=cu�!dvL�����'Ř&�3�����L>'�s�nU�EE�s�'���~�㕠q�_�6hWžכ�uEN�X�K���"\��a��X��x�SD���gۻ[�-4��,��p�`L
�ފ��"ׁXBU4�W1�\�y���dR+���"��?�H$����6�;�|�]�/��6m�#�s_�$n��geg��fª��Ь��8��x
|��WCc1kW|���ōn6�`���w=x]�����B0@z����}	rI������c�úO�@#�vSZ��hw�K[���H����[ծD#�����z��d�=f��6��R�U��Jn�M�r�Ӗ�YR��X�?��|�?5��g�2�i���4���4�nh��,J%ܤ_�޵����)&ܕ0��Bx���ɕ�H3O��%6_!�~G�$l�#��*n9m���&WB�.���~)�ذ��z�qcC��wP=x�ƃ/��6҃��Rz�yܿ���ﭏ�o�&����;vF~&4B��3�k$=��1<�)���Hs#�&�}t�o�~�A�!PiϏ�,Q7�1*��f.niw�\���ɟY\�kQm"h3���w_�	�Wn�	������L�}�^������^�qƹ�ız��^�a��x�fP_y�(Z��YM��z�͞E�pӥM�nJ!_&�ߘ���ʾe��t��s���!X(����0WWE��p���M�Н��/��fl��Oˈ��5+p>�:��[ �"�jj��'�����opAʔ6��Y�]!�tQ��Y��
Z���\\�˼3Ow�ۿ���2���wQK��:W�z����OjL���*�G�)�����d�%�]���@��8�)��rqvhe�X݈�^{�(j��r��|,�>B�)���b����t���c�����8�$� kʏh#�NWI�|̧!��'��ؼ�&�7Hb����4�ZŌ�W�a�!����:�:��]ͱ�v���^hwQz��k1�H�5PN <r���~��6"����cՏn�r!8�;Td�	�Z_t9���[�G���^�HGf��
6.��+�k�[�A�\��s���s�*#�	��s}�:��j�,f@�3V,d�[>t��_}����;j��[�G���e�,��PK�Z{,١ʀ^?˓P�������~-&]��,hX"xN�"n�&�O�8�����<q�b^����kd{�i諴�v_���K��sy`D@������ݵ�|����%��MZkմS�OM��2�r������u���m�3q��}m���%��K�e���gA����71oA����H=ء+�F��!U�H8��˻���u'1�h�bLh[o�$�7�[6~�1\n��f.h�H�v8�;�ż�o���2WRc��z��\�AS�d�5O�=�:}9=��4p���mgN�O����"���I�NO����d��z����;�*����M�.���2
F$+���iN�e�v���e�Rk�숲?�).�u�6�c
�����@�[�e�)<���/��m��vyP����	'YjA�����߅�y[�N=|�,T�?B�1�����'�.��1�x.S+��]j��^v7��Qd=�]�!~
�q%�`N<T�0 ی6��t�تahр����&��Y�u>���$���C4	�y*����T���$l���4(7���C�٭�d\�=��gXt��U���_���(��rSW}�������r��\����+�P��e$pW��S�V��l�{f©(V1�">g�V�*��c��*L���(='��\�:�	v��.�Cr�e�_�8Y�� {��߽n�Sv�g������j�jw�O!(l�@8d�N��Zc����	�����<�4��VE�5��A�#�ioUsx\c����}E1 �;�-��ި'��^,��:�O>��~vXUk2� o�M]	O�OZ�a q�2v:q2�<c��jV��<��V�7.+��W�!'����»S�A3������h ��*�曽S��(�p-��ty?��{N�w P���seN��x�ټ5;f-�^���n�g���8������P�-[V��q^��6u��cH�1CݷMBa*�vg�A���mT�S�3VjZ'4h$�q< �e���9Մ�;\��`S���S7+^fϰ_��0�|��.|���P4��8Y5 `��&�JыJpT|�7OO�WŖtk���[v%��_�e�Y0����Ʈ�W�i��������~�l����M�i��R ��H�񖼯!��z��01`�-έ��kI1}�������^?���:�����|�͒�a��9r�G�q��x�7c��+	߮"�.��@5p�λ�I��~��
P�&�
g`�\Nqs��U���:���'P���*�
��c�%7:�]���r<�^W��gn�5m�I X���n��
��8��
�f�rM�b|�E���&�hK�"q_-�M���B#��k��*������(�%��3>�ڪ�n+�~��o�".�k�$�ܩd�!H�axN��F�.ݰQۤ�	��b��v��'ڍ�g�.��U�;�i4���^�E��������P�N��@㷧�4�+.�^�����[��_����/M�ૻ���&l]aW6�=���(��*��)��F�O/����d�/�!�i�����M�Q�"h�n�8��
�|�d�hf�G�E��􃯳:�L�-V�WC2�Z���,ɻ5H�_[�GQ����:(ʅ5捿���j/:P	��C>~�����Z������z�0�q��Χ�8
�e^2��"F�Ϫԍe	�W9�b�Y��~<��J���������57��rh�!3#N�1�Ԍ�a����;���O����r6�����ˬ1 F��!����=�@-M�+j:����l��MZ$��g&(��[E5Q��5!���pA�h\��!V�����\�m$�k�/NLce�\�I���z�`�Ku�r�4z����mG����	*���p���C�g��3q�q�{쮖��q�J��"�{�b$+W�C$���U�� oΗZ�����Tz��β)�L���xq��J���4܊�v�L`B߽{Ƣʩ��J��rY ���y֣s`����@#b_�	��45B�p>�����__5/�ؽa(��cC$n^���VF~��p�|9���CdZm0�i+5��.I�����!TToh��-";n֊)0HQ�Y��t�;�1��6V�"�]*�ȳ{�,~����<Ob�~n�ț���o8����;�[j�4�, �������ɫ�����^�5�XNai$к�Gާ	=�k��X�L١&~mJ@j��^hfg]�J���x�gD�kx[�w ��2��wx�~�}��x�@����F��]��&h�v���W��D�W	?�#u�C"��5n���"����B�:�8)!���������w����\��y�ZZSC�;��<�����;`��Ġ"�U��ſ�Z]JΩ�DK�ڈvi����p
����/cv��Ѱ�[;�^��v�#}7,�������c�B6(
��|�MZ��b��Ʀy}5'�AԼ^��0$l�FHn �A�V�l�T隰鱂F��d0;�^�'lน��Y�.$������8<���x.�m�=�|R��[��l��hT����ۙ+*�M�qQQ�x-�	C��w�"衭��M�=��v.�4�% F�9����aW���b� �'����"����o'[Ú��|�Z!�B8����}��I	��D���,2:�i��c�t��-����
�sI=��+&l�����h��V)���+Eg�jƠ�|ʑ��\mّv�0�K�\�����Um�lR<��,z%��������ol��e]k�ʜMSK;��d�n�6��N�+�r�Κoo�MG!��TKY꓊V�%����*t�^���|���u��9&�A���*�Pm�:�����@��8-gpߛɁ�R�,ļ��ᶼ�'hA�Ef9}n���(�ʜ1��O|$Y Jt�2��@1��]�A��G3�R�W6�p)��כ��� �:�e��ӕ������Z\�x�� G�Hj��� �P��Shލ�#+ZY0ɬ�X��Mt�WF��Ģi*���^
l?�l0�(�9iѾlɲd��ɟ��tL6D�4=�*ߐ�k	|n������V�~�6���s�~ʇ)}�
��|]'�3-F�OƋ�����U�U^'�Յ�������Z;hdQ�C�x�Z�"��������G(]i�&z}%߃מz#�*d�m`Y��p����K�C�}~*�.r:E "�U|����s������C���h)lv0�X]���x��O���T�
�0�� 7E��ø����ߵ
�.t��Cw`�-э\�bfQ�$�>�^�"�i3taV�t.��4�],��������H���ӌGa���?���'4ix�j���R5�H�e?��3�Tm�$�2_���O�u|@1{��� ��S��B�6,ɻ�8v*l�����.)5�����?
�]�6��W���Mq��h����&I� �5��=(�V[9%&k���6r���@��,+������N'U�0� �����I�l��u�1L�|�w)j�.����Ǌ��<�P�:&�օ�����1c���ˋ۴C�vC�0��
ɭ���]1�U'��r1)c!Hy{�I�u)b�rl=Fk ������#� �*S��%[%@ f�ofF1d�vzUi*��KW#�pOd��ñ�'q��#i�Ŋe������s^��h�^�K�x-�D�E��&����-r�*o0�\S�v�[cjW9s��yJJ%Rv�U�[�5ԓ�B���D�C�XA85��m;���N!��SN͔�gVyE]Ѯ������8>�dB�w�=�dXDi@��~ˊj�H��[G�0ϕ�VڬaK�t,�n����	�JݩG�ֿ�
�x��+��k@/K��5�8�_��	���N�ɔ��?��T���{����~� ?,F�1!��j�2�A]Q߼ҡ�!���Mݮ�z��;6ZbT���x��(O�~O�+����{\�I��ظ����O���|M;q
�Lrl�[�9p�Q×�8݃�C~<��B�¹X��5�N��<����P��2��N��� t��\��Fa��]L6�%sL���D�%��������;�x��BU|�Uy���;P(�S�W��u�kFFpMi��wtf�\xP��0b�r�Vq�o"Lӵl�����B~�\�������CK�6��Q�mud��a�
sYF�L���`�a�Jf���l�Se����o��/�O c7�L@Jm�!����<�I�%������/�mQ,�'�dl׫��~�cz@@��d���Z"�.fʹ
�9[�ǅ:�þ|�S�R������l��.�MH/���W�+�3���\�Tu��<e4r�i�(���&V~/�7Epr�<�y�'>��O˼�yuG0����$�yuOo�7���,3�y�s;�Uo�d`H��3uu��y�����t�^M�?���R����b�؆k��񉽭���1V��Y�٫� �����K�xFK���m��?l�����B�5��}|FUn�!�½�3D�"i5�X���6�wj����<�,G~�at����bc%7���d~�������Хx���?�˿1;;��8>�R: &n��"��^}'H�Ż�!h�j����5����٤lDR���~�
�;f�(V���<3Z��m"��W��ʣ1�pO����������x�I�E{E8�omr��Q,�;�Y�oF���-<�_DLS��\� @Eb+�E,�aDn�o���`ߎ�#���!�0�x����ro�}x�/�����Mo���'[��2��HJ6[J��I���B��(T���+���	/cP'�n]���<���A���G]7�������tX|�*��wy�aޕl8�VZ��S;�Z�]��oZE��`�a�����hI��r�|'UOCb��é��:�ׁёN��s����[���\˯��?S��MN�O:��a���G`���z �8)/�c��L�8��4� v)g�v(�8Bc��HE�䆒�1�kY���o�����ٷ�A�9��xV�oAyf�W���}r��ml��l5سhp(��Ď��{�:e��{�B��PQ!Y|�0�>�D���ٕ	�"��S��Ri�b�Kp��^�)�V�̖�j]�2kK��[�x���b���,7�F���u
D�!��cO
&0B*S:�)�SK�he2�x%0�%l]bW+)��D"|��p"�XS4��p�n3� O/:x�Zn�A���-"���.�H�K�~R�VA�����(2.�$Ɉ��g�xp`L1�vzF~T��UMf	v3�n�n=E>-v�Q ��:h����b�W�j<���=�̸$��Q����I_\�<�aܜ7�3�)���N��?��U`����#������ȇA��2Q1� 	7�O��S�6L5$L̍���Þ�
��Z �_�͉�?9�3������ޝ�W��F�R�r ñ�BwV!@��'�{��')�~C�x8�ƫ�t�2i�Q�9on���O'M��-�9��r��ɩ��n6�!��� |�h���e�<�U!0�X��J�P���2�&�-�We����&�*Q�{jA���v�B˹"Bz�&�>7H��pZ�B�D˜���=�M����EB�6'��dMhN�>�(�ء��y'�FQ�8Tu�3����*Ht#��ӕ�c� ��w\=sB�f��n$���	�a�eU(glCzYl��>�̽Sm�O|�k�R�]�z�52�t�.�F\o�p�pihJ/�_�~�U�^A�_�i�*.8�YΥݧ���O�*YK���Aw����=^�tcq(Z�F���[��t�J�΂�ǎB�	��^)�]:g]�:�7��G��Wޠh���g*��	�ŋp��'S����?p�	��Q�= G�=���	-�*p�%u38/]!hA��/!���)^�&�z
Յ ����с���!��"��/�������Mӝ{��>?9�m� �c��8auԝN&9��^"�vJÎ��TB�˘���p������7��<��=1�ƽ��KD��sC��s�Ըh���Y�5ar_�_r�G:O�)�r�A�w�����2�i3��H`�hEgTd�E��{����Ӿl&Z��E��~.\Z���[��F�$�X�����9[q<�S�ĢL�zV���R+�ٚ3{������?�9�5X�(�-З[aa;�~G�Kv���Z~"�s�ǰhL&���MOeH}"Wq�z��ᒗkw���^�0+V^#�	D�¯�7*	�"�#�w �S]c��sױ1:������_-�Rg��M��:v���]?]�x2(է0m�yP�(����h��m���Q��+B�SL��bn-�V��@���?6�]Z`�.�ƫ2��֑���u���H�d拲�P6��t��Q��e4}+��a��;�N�@_f��R��S�~�N2��|���Z�����TR�r��8h�t�7�\���o� �u��v�3��y2�:b�1���Sq��	�8(�&ط���a?�p�~���m�����^�̿���g����ׂ�w>�)F9��w$^G�Vm�|m�N�sqQ�}���H���̽�Ju����������i�ayrL��r��+>=��ɞ�ߖ��5°��Ԯu;K�S��
&����b�eB
���vc Z�n��pWQ�x�v�����#�b�]�p��Y�M�A�0�����h�d���Uhk1J�r�`4�OKd��}�I��@K)��傅�0�ǴI}���-%e�m�JP����{�,��[��bX*q2E�%���gxp1;{ŀ��0)���spۆN�<��A�
����6�>2��)�.<錿Ĝ�=OR��t��|�v������}*A3>L�ƿk�=4[�7��ՀV�֟����G��v�\e*��ѧ''V;t���lp�/�5�^��]|�#AW)�ڽ��'�:Qk0���[��iF�D��[B����Wƒ�2D�D첹�f����l�P:-[�th�X�@Ɵ{��������t��Ǔ������v��C_n��ؿ��4Y"�{7�ϊ��@��qD؈�+=�u,Ff�NB������K�;�t���⋫o[jlԘ���Pc`h���7�R~O�g��W�a7��~՘������]�HC����ց�ަ`��o3������09�g�x�j?>��Y��稡�,7��Ac",���,e> ����L?8��c�t���xj�vc��9
<�]$>R-����3����H��:ɟ�>8��e��7��>��7�J�������o�BER��Ӻ����6�!=y�?��T����$�~5����#=��DQ���(e=��Gm��ZGw���(�b-D��3�Rn7M�J�BY��]�O�S� N���&��e�WP3X����<�>�����M^-+���Bp#ÌT{�5�!w��^t��_��j�;����Ä�������i07��d���*�]|eT�o��nD�k�0�cH�q��k���X��`�{f���`Nz�ڣm�7���������y�
-�n�y�U�f�<#�r�p���ɲ�ߗn	GϤ2ĕ,!s��x�4��9�%���~�}����G5�<'0t��ߚ&��'|w`:$��|$=�$�&��K��i�(�%��=v�$���`�1����s$��Jh��U:�jjh*5�Y��<�'�
G�������Y�ĥ=��$�s֟�l`]�o�ԀR�ڿF��բ`)���
g/�m?^YN�)͕'t� (&.��
j��'?�����;��t+L��/�3�D�����Q<M��=׈w�\^�?+�O�|>-?Z���NpC��S"��l}0����d��]�����iKI+Lh�`�q�6vW�J�B®�t$��ޔ���Y�+����B?��bCW5B��
z[�$�3���K�ɂ�<\���lN8kE��i�ڇ\LB	�ɋ��G�3���Ec��Wu�1-&���F
s]���Oc����&�JcUjV�dN�;��4��=����g,��#���eN�_}�ci�0IV��H�h�/��œ����V��˙�c���X�<�1k_�D��H�;�"�<�ˇ�n��{pAyfbɰx%�Y�r���$��pAj�%%�>39ŝ A�Xm5X���J@!�t��Fn{-���� �!v�Jy��P�?g��=��Ju#}����@m�D����T�`�����K��)���h�5�,*�CE���\�y= ��Zͮ#<�Ѫ	�$�,&XM~-WY���R���*���0��j�\���mM��@�� ��5�xl��P��Zd��~����6'3�7�na��f�f��q�u:�c��b�~�e������Y��)��f���_�k��l���9�P)�a��XJk�=�sb��Z����	���=���f�Hb�R%�'�^k�j(�&Y۸�������t�z�q,�`�M���P=��x�ϊ��f>�\[�L��4Ԣ�J�dٕ��'��+N�c��=�pAn��t��:� ����/��b�Yհ�6��RZޤh
�Z;-����ڄ�랁5�I�:��9�ST�%7��L��7�l����=�;�{E���]~����+���x?ٓ��T�`L���'�f��I�k������AH���"��Y q�o��!=��lEŁ�����u��C�w��(�RT������!*$��P)5&欃��M6�V�UV��� ��f��ب�c=��#A~:z�w���3�}��D&+��?q�m@��uJ&R�4�~���'��4Cy�u�Z��D�b���n,���p��m�AZ7��ԙ� z�8T�ll�,#4�D,ɪg�$�E�.�V~���Ar���=-95*��'�|����t��3���̼`�Q�䇱v�F�}SŝP�V^>��a\Xx!�c�w�/�הq�r��xi�����-�=mt��o;mnHF��4g*�+���������� O�����Q&�j����U95ر.F͒`_t�H_���6���-P��zJf"a��%d�3�~��B<��?�_�CO�	��9!X2V]��iԟ.�����y��,Jӎ�*��B�k���R�T���Z�r��n'Y��3G�q�ɝ���ѪVGdEE ��M~���;x�GWp!��T�Id�Ⱦ#9��~�%[k�!d���(��v,zr���,������`>��L�n�vP5Tw��b��F�c�"���_�M8	l'��Kw��2�"���FB�Cf�+��@4G1���>�O�G"\�g��ai�蒷5�TK)i��R���������,���@������=��~��6}�ցR<�����`U���v�t�9���g:�L�4B����c�����|��6�j��&�w��O����i.DvHb4?�0=!����`12��v���@.�ʔ����}��HhumD��|C�a=ŇF� M�� ��ﱸT���̬�83���P
Sv���y�c�DO|�z����C���s �{5��X��ǎ_���r#����$����]�&,���=�Vk.Uu�d����\=���	�	L���r��v˘���	���}���h���D��d���N��κ�A�_3B���
�KK�r�Ʌ��&��U���]rj�4���:�b"� �s��m]����2r�Mǋ�1_�.-Y&-�c,A�T�O��� �VږV�e0_�Cd�Ķ@6���[6)8�v�����Q{�Ӑ���.��7@�:�~I>���*��	��mh7~�� �Ô=��i���Ql4_�84'���cVD�p�4f~�je���x�k����ÿ��Q�Ɉ	մf
}H�����H<�qC������C	����w�uF��|�G��C�)��]�!|KC��ǋ�qE�2�n�Ԕ4�>��=��(ٻsQ�/m��z:��7ĢS���TƵ���[N7L���.�lh�X��_�H�(^�=(��	�k:����s�4�S���S�Y��2T�
W&������?N����b�5�I�P�*N�1�X�B�Ws�sIl��䙔.:��_�����r`�ܙ�ߐ]B,��M�(!�mLN�z&s%�x�X�1'�*I���xs��Wo�qˈ5F�*���N��˅9�|���-����/2GE},e���Qc���F��De%�Ւ�bUk��Pk
���qC���u��|@�Vw��ހ�d��0D]��4Cʶ	S�G�^�l�)0-�E������E�ki�ڴ�7�]�h�4/w�[Nf��q.��b0_3@@V����B�k��K�d��ږ޻N��r�}�¿���2�V<u�<���\��Zk�~�t)b|s���{؋��kA�|�l��&��!�ܤ;vp��'����EA6uv����9�����y�ê���l�m���n4�r��Q���V����8��-�Y��$�Hv�����ڞH�9�N.wp k� ��9.<>�)���w��"<k�������98��m8a�6
ȫ妸��!PL�H˸�ض�_W~��L�>	Q�oi���{��_ći���+ؚ5A�YbM�k��O�f�p}�~�2V��:3u��Fq�J� =��Ҙ�i��z�؀���|��S_����3н�=�	7"�c�x����!,����~.�\��E�1��Hm2�a����X� [��ƕ+�n�~v�y����z�L6N[�
,�n�xS�x���d)��A/��P�|����_��(��r[��qʚ���ė �g"�f1Y���Nȕ�d�S~z3�D�8���j�G_@�:o5��2�z�M��{����'���r]�P=|*g�
c���'0=Eh/BР�!y�󻝲u&B)���i�޳ac4�ػ�yS`Y��)�k�-R�M
�1<S$�8X�����P�~E?b���]j�E���}=BM4SQ^7�p.|��4?@{	=��6_֡��I�r�9�~R�T��Me�`�Vg�k�ߎFYk��$�k%ZwI���&�È�`���_�׶��XEĿ��.��̃�%ȹm�������K7P����s��� �A�q�?ѱ�.��H@����V؍+,�-����y ��"Kj�vY��}qH1�
����6a:B����6��S	�&5��aS��1<�0�u��˥���>a1���h�4�r@i���ݪ;��Y<���ȹ���<�'�l��|-$s�;���I~TC�S��٢�j�\���i.� *�Ք+K�� <��|���B(E�9�ޱL�*I�Cn"=Q�+�x@�O�[��d�i�YԨ�]
� �½�����*��l�s������0���iXA�f��ԏx�b��^��+��B���^p�%6��vI�o���37E@Q�]��L�>��پ`��yf:E��v�a7�;*�wzDS4��:������`���I*�6,f�{�q9���!#q��G���f�L{غ�]����3r�����.`5�"r�Ы��ʠoh��tj ���_���ᒽ�nZ^r�a�z9��`�Pp fqU6��ş���D��O�;D��_�?[J�i'����[1��'�wXe��4���I0q ܱ�u�r�-��݋Z��ӣb����F��)eg�S	H�т�#��<&��$�!\�`���z��4$��}��6s^f�[
�U̞
����s�U௪�A}x���`p�1:���>��va���2�����"&����ʷT	�en��.��V@���T���c��e������ҊKַ��1C��b�!� ol/���#�o�tM��ȕ�xY���R.N޲Ȱ��-W&��m�M
b�G�	����S��[}K�G��!�<���
9��T(����;A+WX�5-]�e���>݋A�_��0E=�I��RW�4����kq��*�1m�g���Z��m�k�3��Wo���"#����s���w��$xQ{��4��2�>1o6kTںt��os����X6�{��쾛{� �(�c���'��x�I����/�~c�$�BF��a�5�ɥ^+�.��H4��-p�dA��u�➹h+
���:0k��FA}���.���1鏍��m�5�k����˞;u>�uQ�`N�J�fp���hI5"2%��~��v⼮N�tv%��~�}2�Y��S3�ī�u�zz���C��F�ӭ�:�%j6�ϼ����88����Ե㎂o �b����<@�,&�v��v��]~��\��g���&��>a�䕹zx�)ǻ9̎\ܩ� Xo�S����<�+*upR���K�uKP]
���ˆyt�o�<!�J��d����۷NMG�\�g&��_�%����}�[��AF�Z�x�D��e8/�uAܡJj��s�qt�b�K��=!�h�^L�G�w>�62�CV!�iCԘ�JR��Y�*�ABJ+��%g[�\dn��c�T��z�Ʌ1�>JOcGqI]�!e�nf"�|.�e�c�e6�`KCs-�e����;�"~V�@��t�l"P⃯|�c-��E��4_�]	+����赳��N�9�,��t|I����YW��P���n��z$PТ]u�l;=O����0	��e]��?�!2x�N����%������Q� n�&��XD�t6�����!ٖ5דG����W�Qt���5񷃕A���}��n>����E�C g��B����U�V&7i^���c5˭�l�A\�nu!,�!���
�k`�Q�H",����1f�T%���k}'j�Ԡ1C��[��s.��~�}�rQx�M#Wuk�7B�v���ꐃ�&{8�)��lNk����N����͓�!���څdKM��"4��i'��9k�f�B\�(��a�^��,mؾ93���و]ռq