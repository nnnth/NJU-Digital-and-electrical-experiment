��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���:����~׳�jB%��m2X�p�w1>�j���S��"�F�i͡���Y��q�����\�����\��Ɖ`����Ւ�2_9����ߋ�Ɣ��������l��)�#fa*+&aJ;��o� �08#y�1�A&�F�8i��Ռ]��-��R�A�|?��U�-"E�و��S���=��;^ַB��O�{u������ޜ8�"ا�,=.D� G�����L���P�6Yg��낌8�͙XI�%Le	��a�n�D�
�R��?�z怉��� �8j�~��q�Hc�P�,ŧ���.�2'V��^�q��Mv���g����fV�L����
��C���m٣�L�~�M�}�M�G2�n�<}u������-A�
q������8MV��3 Myz�7J�:S����J�9��!�T �컹��.�
���������0n�'$��f��K�U�Ͼ�.��w%�^���Xz��O�$u�l(�{C|)���L=I�q������m��i�H"+��a�ϋ�	��-��,�(���np�g-)#�?��iE*�-_�9Z-��OL�[2eEwF�1�Ķ�.�Р��P�p&q�De�>��!��HA� 7�����j��m����ϻ�K}��E0.�$�en�F��!���:�`��Dy�� ����&b��%7�#����]�r�������ETyw]Mh�#v���ܸglV��E�Vx�%��M��|N����QC9kL\���
�󾟒�Qj��j���Am ��pE��/F��#�u4�u� 2W��tq|�_B����xA�L�k����@��E7H��Ͻ�6�
����O�)d&�H�h�rѶ���<��m�H��Ǿg�lh�{<"C� �on=�÷��}�vF}b�m��If���$�rA#�X�9l��p�.�hx@�J��Jeg(���
 �k5ك�M� �=��	wg$��3߈���q����GS�Ru���>��²�|�L�.�d��r^����f���8���NtCI"M�xo�ɶ^���s�'����=J�lK��-����cR��4��p<Y�x��1+L,��f��^s��ncW���6�ޱ 3�[A�$�i.�}:+�'�؜2�H ϬP4<�,�89�K�=8*�+a��g�)������!�މbMdp�I������sS��M�N���Ox�
�I�n5��1��ue�d�����̇T�*�ݠ(�6��x������๫�$+9ӵ�+"��+�;�M�|i��V�sk͎y��hg�X��͍�8�I_���9�M�S���S���Da�ʬ� "{���S!e��_s� �S��I�ǴW?~y��+<�8�k=�Q��O�a'�����O	;,
�� ��`[���ΐ+���4Z@!����E5P�
k�q ���i5ujg���lKB(��;���BZ�`�+�\������R�Y����x�CH�b��l��Fn2�D�GnѢJs��7B�C��U��@7,o@�M��KǾ�n�;4a���H�E0H
�Of�b�s���. n�1���n�@}��,y84�8@�p����(]�"~b�ϛw�;ґ�dӽ�o��pq;r�ߟ���p<a��l��W��)��V���J�!�ls~K�m��������Ơ=��ȝb8߬�t���͇�.��4f�a6�`:4E�u{�����y��#M�~�B$�{�[:ւ�x�ō�~*w�0B}���� :7ݻ���0?�1JJCU�sƘ�NJ��1����%�@d���_u{��±ƀ��N��Ys�0�u�c��M���0�\<Vұ�����Gݙ5�4��q[�i�k�I�f��m�K�R�u�����=�x �)�Z���b��C7���	���~\��Q`��B۟_�(�Vuz�/�}�JM[���"+�ou\�1Fm]��=�.
Q �j����G�ԇT4�o��;^t�x�)����f�~
�.��r^0��� �7q�Ʃ���o�c3X&�e�*�1ʣd�f�ZI4���l��3��7�Ƕ֗Z�T���Ba��X����+rr<��I� ��@1D=t���(V�Pj����@P6�nA����ǩř�V�)�3dSP���Q��J[������l�f0:y6!@N��fŰj��rw��5�,��8��ၤ�'�֠��+�爎�����\a.�J�ºǑT�kp�z�h��S{��9�v�x���cJOUrV|����8�?���h�t��O���Y 7$?�u�o���yˮֺ�� �<�b��%��KO�G�[:�Y|)�,�����<���Z��*4���Qۼ|:�[&�#�}'v}mDX`D�+�,�מٮ�qe�wurt���r�R���+#e�m�V��Gp���;��� uQ���U��N]+���haf\�CAH�I�OIP�����̋�8Y�f��pLO ������oۃ�e��qU���;m��Yī3��7��Iu�q�-�)d J�Ba�z�L�����Z;�{<,�>,�HS���i[G��S�e0C"��BX����,�w �<���er�Y��n|fM�m��B�wJ���w�0�)�d`'�[����HYefwm0i�AJe�KM�j����#|���+L��QO�i]R�w@�P'����]\�ޏ�$�(PwT1
�lد�q��9�%���`?�B���@6+�/#���'&���z�b\�~@����U�4� X�J��cN��sy
�����dI��6!9�����40E�y�1��К8��BY�*��ncx^MӾe~�##&5��Ey�p�H�h�����P,<�/<���Ά|���|\۫^�Ih��g� �c ��FՒ���H_���bm�iH�Q^KX�	��O�+�đ�̶�C'f�5�����/?������1 �w��A
��Xǉ�}���ݮޮ�i�!�7`�uGA;�d����ZIb`7#��H�BR"�."������-k�lC&�eZ�oz���Ս�1�-���W����;v��Cя�I[4ސ0U�����?� ����4 ��7N�o���] 8e���f��/p=p�/x#�N�/TL)��k�>�yK��díxfU��ᑹ9�|�$���;��N"0����/�Uv��\���;v8����=� k���[I慘�Y��,�~��8�6��|P���ҥ�f��]Ѡ��lL���o2
�p�e���2�,�^�$���u#Y��i įid����X�C�"�z��F:V�4D�/�p")�٘�<�m�1�ԅ uf�VF��c����	���6藥�DinA.�1��Q�2�9mX�Xwࠆ�ΟO�]�����Id��"@�i�l���#��}V�99�>���$�*�/ec�%�hrs�X��:;���%N�Y�S��[J�L���}�x��g����/�M�?΀\���B�+�+i��k�	��.Ƃ-2ך�Y�.�3�J��j��(L4���W��b�ߒ/|�qI�J��*�D��2���_��)G�<~:��Uq�>>������f����n�0N���f;���޴�@l���# �{m���q�>9K�Q	�Eb戟��{Ѡ���6���䅥áI�B7[V��ƍ)����\Q��H%c���ԥ���Q���k:q�i.	L��u��W�@wN&0h1���Q�NQXdtf=���� ��T+ȄEE��5�ك���b���J�3��Ѝ��BHio 9Ed��gNך��ҭE�����{t��.̠�;l�j�ǿ�qd�\����������{��$A _i�%e\]SIx��Jb �Ns�%{`4��Nf06~:F����ջA������u����h�zrd��	��ָ�0�'�,K��E���d\������߄{��ȶ瓪,��"v�� 	+�T�,�|�u�7'�J�%=
�®���)�P�PdѬ�::'7�J^�y�	��!(������W�^@���_��Gm�Q&�@��gI-sb���D��#X6*�X�@���[Z#ҥ�ΐj;�I�	.���m���0�,1��)aХ��s���\`�qC���ipݙe6\���V�r\Hh�g"c���;��R�����|t��sݸ���y�.J����,��G���=�LY�����={IN����|�6�o�.�N�g�6:0Rì"N�E���� ��){eM�d�j���)?�������F:H�&'�n��OO�Q�~�gvr=��ڱz(%� jkS-]_�ɜ{�c��}���<�/^���}���bq�{{:`��ұ"��Cl��U�u���\���"���nsz�BJ���z����>���<�EpY������"�Q����y[�q8��UG���	�:�Ѭ�}M��XT�6)4���%��fU٠�������o��+�l����h��E�n�9b�ĉա}P-�m�r��j�M��@�R�,yoQ�����}�����E*����J�����On�����%���tyL:`s�j`�k��wO�+;	j��3@n�!���_Y�*�Q�}A^� �����n~�xZ�O&���~l8E����z�0��Szm�D�����&�I:rNXR�~�R��-��J~�ni��_@f���Q 4������Ǥ:M\,�]��A����yX]w zP�y���2xQ*��]�?����2�|�t�-ɿ3kw银z���i�s-�Z�Mi�yw�3��G��U�0��%5���%|I�-�/_A]���K2��S�<�iӛЪ�wH�SY?�b����u7
��KW��w]�*v����0����*%�taO���v�\]����M5?í��Q�p�s)�I��3�C����!���dA<"���>8�.��Mhs�n�GV��O�	�lj���,��3���p����ӣ���X{x	�L��O��p���=I��l''f����L�K� 7�f~�@dJ�YŨҌ��|o��r�m6����3 7]�
\N�>C�^��P�C}��m�Ivjh/�����-w��l\�*�1�Y��@�S.
�[���O{�T#�j׿U;mSG�OnBGzy��ɖ5R�6ji%?d��N�Ba�(��d`�!��T�y�~a �%�0�OZ�*�����\�Z_Y����
�끯ʎ�	ٌ试벇��Ź@��o�z�+����=\�CG��ĭt���n����v���3�����#��J�zl����(32����UQ� �#��V��J#����>~kt��u��	�C�N��rL�J�� �$,����]r3(A��fv�[����7���iQ�(R��®?��M�n��VD�<!љՊ�f�/��T����7��a鸵�bADB��[�.K�K�����<�o��Hn8)�ڤ-��Ճ��xk������E�@��:O�=�lI�X���nob�L�.�_̪R��%Kv6�7�忬"���;?v���O8������*��������Il����':� �2U���y�
AD���d���ε���R+�#�_]2�׳�I;�:m��Z��1�-��c��cCq��ߴ�ȳ�#Ԅ���V�[��^��fE�Ea09�1!���y���I�"�	uV�t6˘�����qfܧɡ��d�JD*�k+��^���H�3 |��]�ǂ���MJ�"Z�{xd/�^|5�����ML��l%m�o$���W�a�#�wf��:9��]��k�^/�p���~����0��Y�iȃ��V��L���I\�.n/�T����G(�6�xN������'���zq~:�7~�'|�
X��!�-���so��a6�+��݊.q����m�: $k�rk{@�����2��2d��Ɖ����M��3׼`�8�� ��;o��������]U?_��X�N��\�	m��RW7"���B����BqB��4�)-�9 5�0<n�T�_�Z���\_�����O�FW���n����;Z2�w�K&�Tf�u��B�UP��Kƭǹ�˰�����Vy��Ƨ���aF���������̹ZĠ42���&x�$�b8N�B��=a�,T�Q���?����C7qU�ҧ��)�2p�8�̭�I�����ߛ�p�����ϸ�J�����d���Tů�+i��eXwF"<���V�+��?��� �pZ$3�ب�h�%�?-/�{ >��6��f>T$�t��W�q���;���o�f����2�N��6�G�IΣE=����ڵoY�.͛v﮵3ju��xI}�4�Y�c�\j ��uۍ|o��H@�JR�4�"���
�9�9[o�)���ЫU0/����X��M�.	�?il��cy��1�����l�c<��|qh�Fh^W'ݕ��xy�􄽋uM�Ѥ^��W��(������t`�����:d���'�!�﷚g�^@Α�H�JN(�~g�$�����Ak1���Z��i5Y�o��d�DU���,�~t����&|�kwtGϹ���4�(�E��}��������y|� �C ��ޑ���>ļ���_�"G�������Ϗa��%5�ɢ�߶`��/�;�u��r� ��ǮL�:!����h>�{�����@�Vuڬ.H�/��ʵ�!P�X���4k6nms����~��
�6�� v���l��`ވˤ��W�[�"�H��'k{m�u(�(�:1��/���ZP-}�3�3+F��z�q�"����n����y����T�b2-�����ߡ�q��)�፟��
��TF0��K��]2�H$���9�X׈n�?He���_"  �h��h��I��"Q�l>q�q��*��,�^�(o� �x@�9�bP�K(�Z9V��ޮq�#��I���|?�0�ɇ��Y �1���w/�p���-;�#���C���n�!<����uS��[��\��Q�,D��T�dZ�L�$Ρ"��t��j:�U!�&��%9����^S�RJ��}^� KGa��,����.PrA�M�Vӓ�z��5�RV�*�l��~����G�3��&�/ŏ#nϔ�<�y6�H�1�o�lqi��3U_0a�̇��up/;G�_�+SŢ*��������K}��eXb}:};|�2���,�|mC&�u@�
 �Ҟ=�;�g�꜏^�AF>⮔����(�M�'��]jC�:��o���r��`yb&ɺ�U`���Δ���릏_#z�o�h1�:c�S^���p6�Ґ��ȶ)���p��0�1��NZz��E�~��i���V�ztꥧ(����ү��zw���O(�� �CN���xw^�{�`k}3K�C� ,W��I�qB�M��-ЏSL��׾� &�"A�n��A�k���3�u��w_�%6�퍱~xd���Ύ�B�C�ΜM7�H�;�������c�q��VH�f�'^��[^�A��;�%E��8Rб0~�����pi)#@!��V��\r<j��{��9xB���_�<���aT/��9{l�6��e����Oř�9�a��['yO5&i�i�N�����l��=W�/��߆��?��ۡk������؃'�b_��|��?ǖ�/���XHI�q��	�ܚH�ZČ5އ�2�����[���TE%�����Yw.̴쨙��Y���*� rʂ�$�t��w��l�
q�:��0l^&P:g�_Kk�jP��?T'�k�g?��-�r��G?|�%���8z\�`��UQ�>�zU���2���@|�x�U�=������p��+�/q�nިp��U�E\/��dVd���.����#H)�Bz�À��&�,��_��{�����Ы�� G:��ұ�A9�0X�$�iOv�޼6Q�*1�&��K��}&�W�5��Y��j7�T��Lɕ�cM�����7Jv:�{/?�5y8�����6�u�BF|��íBo�y � ��I�h1N7��������Y��`*.�vl�<{�K)��Eod^C�q	v�'aDV��Gt,�і���-����#�+�vs�����2�)z������*Ϻ��ؘE��s!
��+&�v;����>q�/�����x}|�6�K
������1�@I#v�U��H6w��Sõ�J��}�(���� ��U)���q,���pf�4�QH19����R�o��?��H����:T)�W��bn�;����D������F��J��*��`�����WO���G��:ߋ�*G��?���C��!~�/F�md�ޕ��֞�f|��K�7t�o&21轷����F��L�aI�W�X�n�[�u(g�
�ږk@#g�B(j�����EW�$���H�&jqx"�ǩ`��m���9��6��fN��J6����>���:�|�w����e�{B��h�jg�6ӗC�"Z��y�2�7��b�v�����:�e�����.4�/�X������^M|%�����P�K��t��x&0�Y�1�q	.��i���6eЈ�0z�6�\�`�.�&xRb5��2���o���4�g.a��6��#�a�,:�)��"��[K��AjW5�^x;���R� �@��츁�#�P��Gvx4�� 8�%��b^v����4��AI>��[r���?h����?.||����R�fMXJs��B�h[��;�fQu���������w8x]S9�e���=����~A\@v�nx�|�������v x/(S��R�����k�E�w4�2�dD4O?��U'�8m^۠�͡�$d!���o�b�3��>Ybv&7�U���\��1O$PT������Q(/�f&��� ��[Or�,�j�ޱ�>M���p�� r�^�ӡ	�8�9���BhFCJ��kw���Dᇐ{:m���`d�����h
�Cc���-�������E�in�=��u�~�����%��e��bkm!0��r��Ɓ�t|(��}U��ZY6^���b_�@�VӴ(���E��^���N'W�<,�����K�e�*j���~�D5��)(���:%I�;W[X�YF��o�7�[ kӁ���i���(��"�Q�>�@"�.;4���S�lM[!B������P���`�rbZ��O�M�2����7�qN��YDm��<��QΎB�n.8�o;|"kA���{��;�C�l����:�����D�A8�P�����sLvy��VG��R���1=R�u��45��rF�������Jo=�U͓q?�ǲ1t|���9�c�����\�r���ovxݶ �����y{��tƟ����o��:AN��7�B;w�h̊,g=�it�.��(@J�i���}D�y�����
��nԲ�$|YE��b!�s����
0qS�O���a��}-SA�`W9���\��:ӡ����R�%��
DeA`��0� ,Utj�j"M�� z�-����)��Ec,�Oz�H��N�7���z�w
��2R�{3Ο�����vc�θu��7�J;D��L�nU"Br&,ԝ��t,f�[��蜺t˧� ��A����a5GX�a�<]���ݳ�sI�F\���������&RM�(�Z_X�z7�?A��F��^TVƓ&E����xI�|$D=$~i�|Ѧ5�-z�ڒD�^K�:;��<��^���8�d��J
�ց�c��,��X� C��3����и�v����֖2D`7�0����e��-8�nM��Be��C|�^#�X!l�9͒;�@o3ES0U��$U.�����3wy�I�R'�C�Vx���𞵫�{m��03g�t��{��rڐ��ԝ�a�T}twF��c���?�{D���.�����{�1'Mh��ԫ���|��$F���J�XSQ�DBF��]p��I�m�" d"5��t60�(L":Q�A�i�2h��B��'xC�<۟� |o"���Uw'�?��.K+��­�"�IN`dz����2T������^�;O�X�����N����Yv#�e6����	y��S�s�����������-^��<�*_�荁T�%e�HE�LK}\��,�2'�?됷K�̶����\�ɻ����{��40�V嶳�: ��]��i�v@+���_0�e�~��Լص0|����g����{&�Zxnj�`'Z��l_Y�%���[&�E��L�^��vi�Pg%p;oj��]_"�_�'"�p�Ȉ�X4��7iQ��{!��Q�2���;kj�/�յb��)�^��Ӆ�ӌ*�G?Ѻ@�;ь��NH`8�%�~�c��e��
��Z@ h]�Ӻ�2��	�%���~�JEU]�Ӄ�3X���r��)9�k��=Aq�v�����.8�m=�+�/R�'�ʧ�v�Y{�k�|�x�Mc��?bU�f�8`�O�"E�Dh-.1)N�:rM�F�j.Fp�2[ށ�0ts.uv(�VkV �b�Tx-�}��I��{�`ԛ9����H�Pi6w���g �5�pX� [�z�6EOA,g�NR,��ύ��U��N�S��KoO��w�֚B���+�N�KЗ�� *�pD�x	p��W5E����t�p�� z�_�P0C8�5��))8k�X�<΂�����b~�<������xg]g�-Z��
�K��o��W�n�JK��l<(��b�\�T�)_�D ���{���h�E�H��cvk�\A��_�~����iCS�H5ȷY�ٰ�^AZ�l�� M7��߈�ϼ�l�9�٤�Tڵ�eB��'8aQZ|�*;ktıD���98�ʗ���4-q:����@»u���C.�65t�F[����u[��Ie4J��I���3��Q� _@{֡���T��}�aG4�T�4;d"��&1��.$�x.�ū`��;\ty�#:�S��&ґCU!g�+�\R�BZQ�'�2|�V��A��)�츠b"��#/������D�v�q��Tv�i��w�CH&4|�8'*��톂.��2�.�wn��W �Juv�g�8�+6����sex��wnS�r�Ʒ���
)Ռ}� H�c�݃��A�w�Gx$���+gQ��
DQ��r3�MS��K����m]��S㗬[��} �L��ĸPvAC��9�۝�~J',�F o�� �Cѧ�A\�G��IӦ_>�(���-���`ɒ�\�-,�&��,�K,ŗϰ�umB>�E�6M�Q�cIC�tW����+���-ǋ��/���
�j?S��t��:|��tU�G*@����@�mP%��5������W�&br�;�w�j)n�M�Ymן+3}�;�l�z$��R�2��,�=�1��p@X=Z9k&uz����]��t��﫡��8�77������g�����{]�c��v$� �!-���H�5����i�@飍�>N��,x`�����O�-A`񰢅���h۪��n�d�]���7��4���YM<B5`q�3z_88ȟA����cP*�֪�<h��r����%�s�.?�n���h�{�=�����0���I3�s��<�ӴfO��Rc	��I���Wر�A|!v�){�[b���+�m�����i�Nm>�0�S������n�l��Wit�b>b/K1��=rG�8"�B����VO������|�x�ˮf�-$@�����9:���>�3,���om��C�}�-]ܪlu�ljaL�!�m�☮B\����~EWV�*�����x�����Zڎ���u��/��~�X+��+�w9�}6W�~�6) �qA�#��v��S��If�X�I5WH�2�~f�g��r83�w��vw#f	x�p�U���^It��۶����]ɑfP�'n���`�V�T7~%����5�8�a�a$ŀT	?Ӯ!���V����[j,���vZ�X\���kq3�&� ��Z�A��ޘ�fy�XZ�s��x�]t��xSջQ��P��4�X0LM�YS��r����v�L�O�ɲ��D�b@���`���4�WF���D�Jd�
��U�Wf�~y��P��,1����U�rhdBL���5��z��TW���!�v�:������?��Pm�R�b���`�z��MեH���i!�`Ns�#�.�����&�p_=oۡغJrS��C�	�e�,X�G(�޲#x&h���5Xw1��������~��Mx[87G	z���E�׋�A����R!�gύ����~���LwF��B)�@ |�����'��1�6���
Þȱ!�NT�*��X2݇D*sK���+�pWs�"C<:ndp@�V��s��|jA�I9��p �0���&���F�8��l�K�64�k��J�І1�%iۻir?�>���a�:��W�oiV�%j�ϡ/:�H��S���n칬���r��oC��l�V�Z��;�����1���fw���0��u����:J��p)2&,��#���,� �{-=�Y��xr{�=�C����y����u�H	�x>��K��?����M�h,������%��OG��I?8��v37��s����4
���$l0������58�|�a�&�=b���&l_pҏ	��*�;���{�L���`Q�Տ��0Y3���oXOi�AN�N�͟�q�uݮ8]��VgAhϡ�7;�0p����?˼y8��]��b��!C��3�6�:���f ���W���8��ъ.�����7�L�u���F�N�<n�X��z��B��F�\�m��5H�!*�g�� ,���m�L-�:h�+,&|1bC�}0���Z�A\/�� &ˬ�~ha��^D�K���:^�;¦���g����2gy��$���u�{��1}�������i��l�JuLGrZG�L}���d��ٞ[U���M���H�M�u��8vRc�γ�%i� !äS�2�Δ�����'�y��0G\���x;V*k��wě�U�cl�Am'V(�_ͯ��o(�)d��f��O�j�k���y��e@t��N!6_�9�8P �⠜��LIP�_[���<
�� �b��'�0�뗀L#�c�����-��rz����*.-�2Rӊ���U�!�]�-A:ݎN\	��F�Q���r�]�{�� ֶ��̭�E�xa�fR�|��l�/\�_<��r��C�g��E4X�П	���| ;�b�um����n�9����r!ѝ�w��VW����������^׎���9|%j+d�E��ᴗ����9��gY��k?0�hT��h�x���&��񞸚��_;uW���=F%Uf��#9��U��"g*ê?�2�*��5X�d�+8��+�d�})�dmtfgU�2�t�m��W^(Ci�O�X0ɴ8�7I��c��4���L�{�!@���H�ۜ�@Q�7���UGˎ�%|�����=-�O�����|6e��RG�����܏�i(�l""Ě������$�ϰBW�ˣv���Q�I�h����W���g�ED���T���������v��(*E�v���s�ggT��b���X����y�AƧM&�S�no��>@�6��0�X��s�k���UW��у%3���@]{'T�J�5@���@���`�v��~%�.�cvAb ?�Tz��xI�!ЊAo.l�y>I���ま��rn��@u��y���hc�/���w���ש�3G8�F�Ft��N� ���#B��r�.������!�/�mհu�ݷ�Z�q�YM2E,a���p����%yb:wm}fw���Zm*QƑ��xK%Xh��ă	2v���%�
�r\���T�1BH�Y��=p��r��*@�Mo�X����4NTH��T��M	�|ǰUds�{��$<].7��,�O+�=� �!���f*f�Gu%����"�3bC]�=��� *����_OPJA>���K�����196zfWrW�1ô���&w�N�r\U�{��J1�2��qBC���.gH?��⡘�8r���
��V����\�H��]+4����c<�Zk����jk�cs����LXV�*�).�F��}�C����ч[�So`�n
�Q�Z���/V�zA!ؗ<��{���#�V�"
� ~I}�#��9}E�8�\�IW���a#h��K7F�����a��/B.!�l�g���1tt�(KtW֫��1�d���E
!6�'ډe�y`~69#�n���ϙ��]͡���p��E jYx��s$t���	{����瑗a1-��c�qX��{y�Nŉp���f�,0�%� <-����y�tfX�n�)�4k��N���ǡ�L�3ƻ'�z���Z�@��a��:y�6�E^���yg�Auar'�`�^<."�ΰ���4�{��?�
A���� Bx�2&6VMA� ��ըz�����7����]W� ��.�4�|�B��{�5�?��T���{;ac��l��{���{��A����92� ��NĆ'kع�'H�����[�M=�r9IW�)��ٰ��Ʌ��l��Y,�3�4��9�|��{��[t�S����Z�v�!���A��;������a��{6K��L���ԍ�O\RJ�
�+��iu�_n�_�H�Y�]j��e7��� �\ Y�Nz7��+F���c��	�EKKo�U�B�.z�%�����#�rYP�mC��w�-Q�h�6�ꩵw�δmdɕłM��{���@���4��<�F�+��:�R�3�A�5%в��V��Y�[�\H�B*�U�_S���!1�ME��Ja�ua�� �o��|�W�ӹ�r`�!���1Yq�Ɣ+r�;ߥ����)��*й���nanP��4W�8������Vy$�!����vD�㇑jv�<�H�䄚�'7��[=�y����A��G�A��zxH������h���z0M�^'ٵ��z���w2f:}0��FJ�ouQ6�w��>L���8��^L3�4�L�Rx��W��C��4 �=vd�`n���q����o�q~���X�f ��F4_�މ���Fc�V`f	
��������Ƙ���"�kwo�@��>*ͦYQ%�����f��CK���+,�z0F�eB� �=*��z��,d��5�/����]uoX�>�ӊ�N��0m�k��.����!b�L��o�g	/�UR	�aڴE�8ą����W��.H�|c�g��fÂ��TVE��A4���;Ƶ0`O0a���Vᣨ.&*���av���٤+��?+�Pb+	D�揄�����+����ErkaL�_mE��2ːra�Z��_E7����7��q2��8���߱((�]��M�gz�gPA[d��}��8�)ш$�&�����tf�Û�?FC��Y dԀg[�J0�_L�t�C��קU ��T���%���$�oX���?��+�n��y�O�N�Gs���;s�Y<����Nʑ&��1y7c�N`�$�X�e�(���)���D�.:'íT��E�ݧ��y��Wxn'j����ӝϬH�N�ayΉ��r�/�3�a�ō�A!�7b�%@�lb.�۠bC��e�WC�D�;g�� ������}��ݣ��C���L<xM���mc�̃��Z�#����FI��6�e���c��%������G����9�������x�Q�ᢡ	퇦4�x�'W\��t�W���K[l�?[=\8���0�+�q���&�YA�����!�'Ӵ�)��x+ʘ=ٓ��B���J���Q?�=���] V\G� /��_j�W R�}A���Uo�����.�l_,&.��4�{?����J�z�'踧I�]��Ƚ�lRt� ���M(F��'x��5Ǽ頍4��W\l�#
n��>��*�h`䀢�,W���6��4{�n�9Q({�,.h�>���GAt5ʄ�v����%�M�\aJl�3��[��lYd�15k�ɦ~{�>'p�z�`-���ЭT�nz���sa�'gA&7]�#�y��I�8�l��Z6�.���
�D�&�Vճ�_/F�k *�i�.��VIC� ��S ��~�j.�do�=���I�S�H�}N��JXzM�+����ߩ��%^�t7*|��:���lcQ�4�����+.���u��Pxz�mCB��	��x��@!�4��V�»����l�8��=��Ҁ+�FӒ��6b�E+ITK�z��4=�w�s9���8wT(�ݬ@�AM=�r�%�$�\�	n_���P.CF�Cѧ��ؼI�kCA��r��<�"E����H$8��w>�h�������9g:��O/�6����|/ќpk߸������-��j:@��-��.ytp\&Dnmo�0{����;�\�����.���c�ę�|��B�im��ǌR��n� >�q}� +��3�L�T��������%KX�B��Ʒ#Y9�G�r�cat���j����-o�P@�l����%�i,��&�d�4m�(�
���=7��IG�}�v&�5�'�Rw����6�у%�/�՞=����/�T�Ղ:��Q�>�
�T��Ǔ�N7�$�ϣ��  YG#zp#�?�"�f��F��_���h57�P{V]���c|ϝ�	}����.m:�'�0�z�e{����`G�\�]�Ew�P��23m\ے�~�>/t�œ!�36��0�i�NՏ*z�4����G�C}��&h�j��}u����ݱ=� �n��Z+���MF��K��ӜM��m��r�Ħ���|�gb��L��Z͌�E#�8�@�LF�n_JX־wnc�4gM`�FjX�&no��7Hh=fG:���w5�Ōo��M��o��o}�ad�K-�uQ�8y7y�k�]�kl�Y"���im�i*�]QQ��1�@�2$BRwȧ���ϳA�um�W��6&���5v�!���`���ى�g�</�خ¡��i�ѐ:���6�Y�#N��w�g�2{�(4�+��[;� R�h篼�>q�J.�5��� c��7J;�y�@Y]���m��4!F�ڷ�XV������P�D���_�}YN��5Q-�����V'�2ooI�Wl���0գZs������]>�J䖓Y5�������b�_���ڰ`�ֻ��jm	��S)�9��=���l�� 2��a�)�h�/�!~#��d����s���o���I���k�+�{�3��bö�ڒ�v����aUv.Q�ǻu7�fwPÉw��d��R��_���������ʁ�	�������yi꼩&��?��w*O�]���
��}[��0�c�e�	�]���͆�����%�{�	�s��섌>G�-8B�>b�3�\	��}B�Zw
��M��-�4k�Vw%!*-0�0���-<�Gy���r#��x%�|�R1o�;w��nu�������0����X������k�܀��La��7A��M�FQe�Ϙ�kk�IA��I���-B	a�����}��:�f����Е���k���"Wdv���Q�aj	t�U�Ո��w#>�!��c��t���n���ȧQPq-��ɔ��t��A'ԣ[F�"��ѷa�MJ��@��.��V��ޖ�!i "�G?V��1��¢F�l1�g8��I8��5�Ƹ{e*��� �/���`�WĹ���}lG�o�|
�_�S��Y���n�}���0�{��&T�a� Q�<y�3���b:6�B�	4c�7V�d�|�=�6��	�\���VGdd
��;�Ԑk��fx�u��bxZ�E54��pP�q`0(�O�"#�����v�rС�e*Z�wZ�C�>7'YB}s��^ɥ$�$��� >�t
�t~Kσ��������y�B������Y#�������`Դ!�����L��a�M�b�uR���7)�]��*Ia����.�ޅq0R�� �֞mE*��ͤ͢�u=ɺ��f�>�[����!�S.�{�B�`��O�u�>k��r�{*�cH���:G*���<!��Br:��d�̎��ވ�jcb�*<��T�8s:n�I����'�A;���f�;�'�����q> z=��>P�A z� :{�w�����I��B���>��5dSn��6ș��4E�,U�ݝ�'�J�B�>�B{�)�ͼ_�f�0≴͐��蛔��}�Ѥ��r'��G���1d.�������_����֞"�@���щ��s��Pj�TJ�ր�j�lq֫�h�jW�%g� �Bܯ��/K�,#
��-�͔@�:��#��#���%&���[yHYD�^J���J҈��g){�6��n�[��"$��`� �$��⥏��K?� �ς���G��Ew�qy�u~�7�E� ����g�j�Ej��`g�S~����KC�yȧ&}���y��e�r�c����Q~pM|F{�04�;�IT�>L|�k��4�ơ�~���nϳ�U�����AEϵĴ=}��t��n�덊��f��Q֩�me�j��7��Wb�nY��8]���=v�A:߽��KVSK��Z����xZt�KH���_3�k��_�b�(P��[�7w��(�5�\�y+A�
�G877)9Z��eI�C���GV��e�cvAD�|;��S��!�(6K���z�r�V㠑9�bCp��-#L֭L�C�)S%��Ub�Lw�pD�c�W2wi�P0l=:���'�3C}��mW{ F([�t����=� I\��Bץ�%�r$����~���qk4��)Mm����2C��:������[�8Q�C��e�S\��ʃd�6���w�����ei<4?ؼj=��G�0	-÷���)�
�1���v^�Oꆎp�r$0l���CT�����0��h�i̠6��ɑ�_8�?.��(7(uJ�.Lp��D <�Z]KLQa,U����&�#덄Q���Fflct�
 ��uLŖu1⾸棨g�`y��? �4� (=QH��4Z��Z��2[�4	����(ů }���	`�+��Ť�l��xq���{�X�8��+�)���=����L	�
�����h���K ��c�.��'�����(��!�n,��_[<��8�'>�i4���CBSZ��Yk+���A2̫�}�P�g�*�9���a�����e��`ŗ�[^"�XwN~k�cR�C=Hb@sG�]ώ��y��J,��d%4��+�S����]6�e�;�X�����Yg�ǿ%`�6���%���d$�ŏѡ��g�KE93Wl�Һ��^��~[r�H_;�ΔM؋��y�n�h �;�"�q8����ۗ��"����)|�lo��`�e��8adQ�S,���Ь}�9Ć�˓2��vY��<(D����q@�/�g���������<���*{zM�p����ҵc�{e[ �Vh��
Ľ�f��d��`V���`���l����ǁ|.���p�X��B�Ҕ.��mˉ�G]�~�˗ή��������lv;:ݏ�{�69/��	���}Q��KF�И���'�5������tG�uyͬڰ!�QN g���/��TB�����l�%�ch�aB�r��M��E�G��<5�S ��5kU"�u|�9+�&�[�#�S���a�(C§��P���MJҸ`��8d�D��� ?�(�AX������h��l�Ʊ�m=4��[R+�6^o�32�X7 '�í������u`;C�����35��󵼵Ҍ5j8Ӷj$1.���$e�˸[_Z�bH�� �nF��K,���W�+�M|�u� � #&<g{�Ĳ��H�6�
 ^j��V	�[":�(�`9�=%��x�	��adHxMl�V���� �� F@���6�NV1{Y�7�u�{��m�h.� �a��&$ؔ�`DUO��;+���.ED,.D��DD��֕x�+���^e�� r\�
Y������5<|�ل����D��=�4tY��_��ۘ���L0Ȅ����t����/�Y�I�����nO��O)�pֆ�&D梔zP0	��d}�a��(q�V?����(F*�.Y������4�0�S?��$�������V�ks�v����e�f�A�=�¸ӈ�X�3,��,;)#�P���ˠHds�p���'��Y�S�`~��PBt��3X�m>@��e��w,x�o��^�m�1��M��>j[H{V:����=�~�#�:yw���,�6��*�
�[!}�]Em��$���,�'R��i]��(���ݡ���h�&v�d�V5�޷Aa���{LI}cP�� �%�$�=Vk�DMP뙈	���j��?�Ѐ���S{|/�*i���V�����}�t<Z���\E�oV����Pe��<���Q(ޠ&|�0��� H�5C�Ҿ�
.AI���v�B�_��|X��H��ُ�>9����)n-6g@.fv&	۱g	�i��^�����D��m��YP������І�D��|�Z��{�'�F�c�D��5�=��U�fIC���z�clp�FN %��+��uQذP��6��^�������.uns�p;T_�,�y{#�렒�Ӵ5��n�逑Ss��7}����#��{����!���a۾G�9�����\��o�o���L6oFB�(��{p�X�F2��/-�B�qX뒤:,�Emd�y)���4Җ7�E9}�*j!vMp&|R'Y��;!؁����φ�����<�v���	��֒e��A�����hT�p���]a��w�vq�Gݿ���7 �������҈*u.HI#�7!=�E�1Gb���p_���ߧ`-�����Q�8�	�o-8��d�^,��Q�r>����a�,8FI:��<�k?Tu�v��Q,ɪJ��4SI��Pw�r�K�DH��Ía�+5��
�lD,xtw���_>b�Q���Kn݅[�T�����"�S���m�3ڰ�(�
\C�ȧt�OG�"��(�t�qnll���/7(T����Fat_�0��v�M|-Y=w�=�X����6�Mb1���Auy&�E�q�e��*Lg��]���[�S�ς��0X�	�x&�WM�>�0�H�w���-�=�ʜF��ҹ�]T�0`z����qs m���j�,;��)<b�^u2r�'l����y8�޿b;u
��MU	���p�w�o�EWX�8[�rs�Rh�h Qr���*�v}�=�����c7H��I����0RyS赠	��	P���Ǘ\_<�� `n6��
Wֺ?�C�:՟y�E�wx�!m��<y�/(3!+WE�:���T0M��Z��u#U쵂1v1ƍ���V��{����y�^��Z��(7��F��|�� �X�(W(�$Jh�WPz��C��Z��2@D�����K� �0�O�����Uo�yD�L��Љ��Y����q+�L�=k`�vRؾ�n�z�a@	�~�68�3��۸,{T��8��e���=����ߧ �qa��s��Y��6�9��ڞ�5��U@�3=.?}�m�l�^��EB�T%��o;(����� 95N��>0D��f=��{ �"��!3>:h�)��&r`���T���=���ռ�ms5݁�M	��tOdog�<T���#+Y��M�`���8zA4��!�Xj��i��E��(�ghu���J��w�;�wJ`H^�<�>NW_\��"D@��f�����1;�Ǝ~�>�PI���1thz��x,���Mv�̴��b(O�d�`���LkL(�Y��X���͋忺.����8T���&���խ/]!=h��B �x��4�� e��l�E5���uN�+��J�N��iV�ɨŝKI[3� ���iڬ ~y���ˆ�U8�)j�ܝ��֟3RQ?iL}	dC��2W9f=����|_��/��U;�	��-��w�cd�s���)C�_X�L1FGB�n^���4��;��-\R�vƿ�4�g؉��Pv(��N��i*���A`��pOD߬����	����jwEQu��S;��(�~V��m�Xw��ű�bzѶ��� _(TF��t���⎘v��M�!
62�P/)���_Y�C-�!���i0�C'����0�^�����3^6g�6���� ����?�j0�a3�4߃�3@����A�XI��y!����']9�..h���gV�8GO����T�=�o����ۺ�������)��ƢJ��W'������*>���_e�Qn�v����X@81� �*��0k�4�813(��3�"�1O��W�;:b!��m�b$�C��;�S#��v�x9�];$��:eI�S����8)9S� �Q	��Z�?���LUؽ�a^���X�>��fB{�p�����]VĐ� %����?L8_�ꚼc�*+�]b�(6
t� �F�tX�$b��/�(���]f�ז,� (.�35X^���e[਺��:���J,�v�rDAf)S��[��!�2�粎��0�H��]�x�'�
LX� ����^�jk���d�=0�DJ��������/}a#}a�ի¬@�1H�J�ݝ�C�3ef9U�fs���tIPd���ٕGZ��w���2ssơ���  �|ӳ���θ������4���|}fP̞�j�	(-4��|Q@7V��+���WF<��ꮫ\�X>ת���	�Q²�]hj	Ց�k�@���K�t�)3�~���
��G	��l`��ƪ	�G�д�E%�1VEP�fZ[�bT�|r�x���.�e(�Q��lf㌚���Ț��n�·<sN+�����6Fr�87�p��iG!t��
-l�{I�"9���z]z�(�eG#�P*��·��I�ϕ��<2�<2Mfǂ��p}����jaѢN��[9`��w����/�<�*��S8�mSu�pR���*g���{n�U�s����V���V�Ag|x[~�t%Z��Q��n\F�`�L`!T�{A������w2}2����{�t%qU�.��n+��0���uXb,k��N���.���e �V[pC����H�:�;ډ9����p�C�_�+ּ$%k8�T0C�M�U�d�#]њ紺I�b�J���"/.�B�x�@�u�?��SFHJ��lQy�m.(4����}ހF��/�E�Y��?��y#��(����)l�(�����ayԁ�Y�tE\����"cf�	��i�`�A�����5[XWآ/�a�F{�=[�Fʩ�����V�C֟�"��(7.�Z��N�Q��CE��E=��1Tזkċa�"��E�U���o>�S�'�9���X�r������P�`�L����g�#�ܨ�C����ş�����&� ��p�y�$ȋ�<���� ��-Pl�۲�(t3`6?ĸ�E�@L5�z�'��lM	9H-L9ADZ� �C�r5�F뙶�"&�Skt��s�_3�ӝ�C��g��L�&�� h����ң����O"�����.mu�'D_�r�=s��R�b��-��ޢ�Y@7�u!�5�=��*���m)�Y�
�;dk�����XM�熌;�H@Ԥ�`��GUrTw�7�J���S��_ݜ���f��"̿1[��%Zb�|��D"`�����n5w�r�<��_x ��i{�1����������ئEu� +K�[��4so�'�@��))̖���gyn�O��	�Qc�	�p��rB�����㨵d%�n�b����>�{��V�}��2]�kՎԁ�c�M�g���bH��{:u4��}C� ]�?4��ŷ��i��Oε#}O1KDq������!���t7���ǔ�I	���m�ܐ���h�6�����1*Վ5-�	��is	����,BoR�P}N|"�7}n�;�\�Y�����yG5�)�ha�
�,�[9���H]\�P�1����ɜ	�р?v���^?@�g^�\�͑u��9 ���'����6��=l�Ȃ��s]�Q*�<��Z�f���#uS{����d�¬�)��gI��ܽ��w��Q�A��_.�d��#	��}襭��f���i'2�t�X׶�<ᰐ<��²�]ւe+���aOX��3�l�s�4��8��)Gl�d鎯��̓#>�^���<z"�Xq�
K6
*
�P��# 8X\LZ�]��kX�̵jO��V���C@��<���瑽A�^� EW�G5�L�xc�)o�i���½S���N�2D�|D_B���(oHD��4�d�&8�,����8�
*.K6 ��
��x-��Fɺu���6�Z=���D�bQ1^�o�UO��5T�Úݠ���j��
���7��"�:JN�6� ��ЦJ�o��w�OϾ�`u�l\�C4G	�>��wFS��Ř�?X�)�֑d�0@ګ�$J�.��)?g��<(_�Sg��p��=���a0G�O�!]8�/?x�IV�Y�����bnK���������9.s�.��N���@&�1��ޞa����jA٧BcӲ�l��2��qك�ew��,/���]�����ּ�8!pC7�,�y�x��ߣ���&���-yޑ����VƗ/���@З�}ޑ+IS�V�R=�ahEf9�Lق1TB�B��|(N�b�`XW�G�z�An�O�$�_��DN�bB- ��1�ʱgɘ��.����B(2jmRga# ݩ���~�3�ƭ��f��������ta��=}7f�� <�1=��������	QP:���١n9HO`�4�xr�������� ��S��
z���-���Z�CE�?0�U��9L�u|5`�?�:�Le�4�yK����rޏp���>�s���E�	Y�=� H�	���Uh�(''>f�PD:�]e�8>#a�Xª���n6E��~�RH;������/�֫GJ��e3�**��T_�/��f�c4��pr���!���*��j��
�Jv6� ʯ�L�-�E��s�ڎ�Z���������jyA���q1Ԣ�ԣޗ���~B�Ri��F6� �[������>��7���6�"(���rH�p+S;��,5M?������}����nf]Y;�l���y�V�}� g��=�!����~{��4M�k�~ٙݓȦ#�7�m�j���.̨+��= �N61��ʏ���3�u��@6����J�zb�$~��$)9�1g�=
��R�)�| `Ѝ�ʩ�)l�d�B��w��N��1�c�\O6��͏��&Q�E�ٵ��mA��,�1&�$Ra�`rh�6k+��3/yus��
?��Jְ���!�!��E���b�Io+�]�����)�����e&�k�s��V#�"4ѧ�!���zW^~:��Т�=����+��;�׷��J���̀wT��C)�p�/_6� |F �/��Xk��p
�pr�L�B9uP���!����3�.d&�FE�2q������u����q�9S#�}���	����{D
�-׀�r� �ޫ��Ru��O?%��Y�<� k¦&#��^?7J��9gx���~Yk�@�BP�G��7l�ׯ�0����]q�YZ�����*�Z#����25�B%j����P�l3,*�Xu2 ��:�����n	,3�vY^L<��1��J�m��訡�n��V�z�1��qz�pN0����E��H��d���~L0­>�f'2��q����D��WAkd��׎p]�2��Oy޻KB-�E� w��y�Ֆia�H��>����s����*���h?�k�VZ}6�6R���A2�~<=�t?�[)�A-�Ů�\%;Ȏ�_)���0Ϡ|ޞ6�����6p�''W(�"�#�	�7�5l�����RH�|�� a��ᝨ'�E�������#��}e�~i�P�E�Rܶ��`m|ikBwM�6�Ҙ��#�̑���m#�7ɶ6\Ԭ;�r��Uq�+oI�V&d(?�5S]�5˦�jޟ|a��\<~�Knt�}�ݪr��Bi��+'�� ��2�~�ދC���ns�9㌝!!(Nn�b�dƍ��l��cRW_��wՉUwa0"&�\Z�'5s`�����J�#V"�;������INac�jc���L_�vB?�����ŋ\v.w���C���ѐ �	x��TRd 1[~/�>+�
(�s�gaܘ��.9Ƽ�I��|@�B�v�*���U�	e�Qa°��N��ۆ��%0�C��$+�L�H�Ѓ�� �b@Ő7��.��M��Tā�nW2�4�ru�^ VX̒�٠�BL�o�$dj��n$����LU��2�����=�&�5�� �$�sh��\�Nx
TB��G��X��$���$H;V��A����~�y4D�:��o��>�3
Ѕ�VY7Ȳzٵ����~p�<��spB!<�t�_^U%�pԦ�!B�ܚ�`X�����u}1�y�2=�7��h5a&�h�G7k4�+:*�k�����:�ȗ�/s�6\Z���M�K���3N"�C��jjN `N���`u��+ '��d%��$v�����H�a�E�{��mY5� )��D��sQ�#���p�+�#� ��䣹�]<�j+A�5�_�[D� ����B�scx�P�Q�Ąv>�D���k�
.[݅+>��(S�������:�byE�.�hV�kL�aP���)���Xh٫,�[.}@��eO ��b�T��tn�	;ǋE�����A0j�8V��7���einr�К��ԧw�J��������{R��kү����<�t��Uk�F��,�AML�iAS�Q��+TV��;hd��x�cE��_9~��C��#�B��WAEaGȄo=qi���u� �Ԣ`
\lD�J��K̯Qn͆�~�0Jx��m�&���\��JGu��&A�go��0�
>�la.P�ڐ�w`���c|ϗ"��.q���p! ������9����ď�Q6a���Vғ�.�����H��(���c��m� �F?���*t�)�x�Ǳ�ՊR驕D��>e��׉}S�c�p�|�I/��'|6o<��Fm�!J��A ~S.�\���Xk���ƛ�O�7���T�x�2O��^O���
M_m�jc`�����]e;���7���y�kڑ��ŋ])��2�	M���|��ݶ���I��d�@�rd�J�V�^<V���#�J���#���x^���k��5�i��Ur^'C� e>��|�l�>#�Nw��>�X�|�d��g�<����ش72&c':���vD9*�Ad��c?ڰezPh��y�T���&�¤�����9�S�9��Je���g%V��kh�n�9��сS�%�/�Ur|M�W/��+��h�������'�d�|�7@�R�A5��_�!��5�-s%FgiŢ�!I�p&" g=J�K�;_]o �,�8-�(0;y��7��|�5���8KZ?�YZ���������WH��Z�|R�2��=u/�6��B�{��u��WS���(-�m�*���j�g��k������!�.�؏>/��Q2�������Go0Ⱦ6�o�흥�F|�y��C��,�8����qKHibwIYE=�g����k������F�/ ��G����j];��TW3�Df�D�bX��kL���LN�f@�|�kT�����G��h_fd[c
��˰�A��~�1$���,�����Ǉ0����$�<"v7[�y�`pb�^�2^s�I��k���'�f�`Q�L���_��l�<|Y��.���6H�So�"�#]?ѥ�����/�Zل�������1�ɋ�����̻��C����<���NB jt"ܣ��%��e�V�܉��2l�kL&�{�ڛ<�u ��#�#Ȗ�V��p���[6W����n���
��^�!���Ń��h�I�����p�7�z� ���kr�+�p��+J
�<���c���>T�˷���^;n�����7����\\E{�~ٿz�U�5j�ό|y���>��E�A���z)h�O&H�����ݛp!�n��{���������p k������#dOA����<(�'��e�hO��04�_���!?������u��XQh7�ZZ;*_R��L��!d
L���W�2'��J��OW�!�(ހF�f�w�p��Tg�q*m/��&މn�Y@@����Tκe~�0����j����$B�:�Q.�%�����Bkg,���t�����9
�m�M���߬ȉ�5J"^�gG̨t�!h��S�ih��#�a�<��oRF�r�|�N$�A��JX���@h�}�Ɛ/��b"}s�:lOd�6���V2������<? ��h��5�2� ��dD���$\`���b�X�7�t�+��Ϯ��R8���l����T�k�����Y\��Q��ñ8-�oYa� ���o�5���3���2�Fͩ_������^�uw�X�f��ʅ�����Wb����V[�Y<!��F/BgeBM&�h�����2�l�[p&�qV�X 8~����3j ��M����[���� ��-�-�M��(,������HC ���z�I��H�ᚰ+���{Ox2rX��\a�,t���RF�	��F�.����)ض��l'�^"�h
��_���q����}�a�u�̈9l�`  =d�g�$MosM��֛=�E[�B��1�>p,g�J�{��t�I.���Z{���민ʡ�0P����=b�LF>�¯\���p Pv�Dy����}�w2=�Q��=K�Ǵ�lh�7��k�Y��~�'7�ɿ78z�~t�?^1��f��qjѮq�w8��O�S��AC�ő�l܄�oM�˻.�G����J�3�l�ZH���� "#�FKԺwa>��n�ϻ��k���n۳-E���å�A"E�H;��e6)�����FW��k*�g���I�Ё���ZJb��!��m��F{��z*�eX����@
y�'�7ܻߖ/�s�Y[�ϏI��ud����9�7h�FWo�$Ro�Ew��h[iV��%E��-�t�o,�����}g��WR�1OI���ʹ+Li*h;��W��c��d���EO��kL�wv��zX����uw*��@��
?�W&e>/3�_Y0��� ��l�X��}l18�ȴ��~�.6�+�\p0p���C����p��-���;]iveR�v��	�98x����(��T�-G�=��nM����?��ؼ������0}b	2�r�������M�"��9	a�	�A��RX�}ő<�u��Yt~MU�
�m�\��2|��rT'�Թ�G�P�rc�}��j)��n����:*^^?p���L�u^`9�̣*�G��Z��W����"�Σx����`�gلIYB�F�^cқ`�ɡ��
����"/[E�&�n\H�$��)�Ph�#G�����:�~&h�E��-F�4�E�����i��bp1�cY�@�e� F��^Qw���{���=%�{De���=�����H���K��g>�u�-����95^��� ]�bxn?Q��W�k�|%��r	���9r	��L>��O۽Y^r������)��s7�V����{%���zڲ.nJ&��G��H[��n����+�߆�0%`{s� �����W��a���&#�U����Y����*n�jSU�d�B�Tz2¸'������طǈ1�E=��$�䁨�>�M�'[ya"h��u��s�<�>g�Bu��l���z��&���碼-�s%j���c��"#I�|qM%9/ע�������e��Waf�$)C_%v�����6H`K�lz)*t�tg�=�}MYQ�[�SH;�b�@�*���Q�Y��.�8�hԤ/�G��{>��ju���g�ڰ�G6*D{��'a`��U��\����x�%�+�����>E¨�ρ(�kE��o1qדP�'�"�]Ӧ��׾
�=%cR!O��G��
o	߯��V_ ��r|�����S��Oj��j�0�v�D��[�Q���Ұ�.?n�Mbt���+�6�q���L&��x�����IO���I=�P�� ��=�|���H~}7b��&5���\�~����ŌB�v�{� b߻�"6��~�Ԏ6a{nXrb���E�S3�Ojnl�ӧ�:�	ے��kvy��Ww���7�bp�ɉ���k�f,_����9��?��LaWD�ii `�%�m]��]&���"�U�=�j��B������c��c𵍨�jd��j�m�Bݗ_��;�J�@�8!��)�*$QΛU����Ǭ�
iyݭt)�R,h%�@"��I�r�Y)
��eڅH�p�}�����3��V��(��x��c��>�ԏl�:�̹ᷲ%Y������w�v�����h��n�,gF�����^.���a�PXN���G9g���h ����O!2����ۀ9�껄� �m@ l�o:gđ������0X^���ْ�B
@iz+T�ȡq�� �pys��n;�l7k��)�
����*��1������)�o���q�kk��f�L �����i�(��CK�Yl��~���ߡ�
���⇐Q��l�7�[a�� ���y.�lR�����P�V��r$n�\����&��t@��w�v���:ZJ���Ԁ!�>�`�Ht
�e�&X��A�z�"F(��zC,��q�K�(\T#��;T���x@�o�ŋP�l����mO�ϑ'��{���l'�__��܊H���Y5�����3�\񃡂,�%T�!	g��┍�������F�Ҕ����)�����bQ5b�d|C�5���R^h~_�i�^�e���*@��eRN�ke�M�2g��N�gߵ��ɬO��&AlB^}W=�\Ɨ��߬鿑��;rv�yq��|���,���10g�1oy�7lW�RWY>��Ȼ���T��NE�᥄4�P��=�.9Gx{�X�)�"�h޻���~�r77�+�w��O�i9x�Ch�����P�b��cih�
����AuTL�c���n'G?@e|�t��D���L��`���̤Td�(>�� *<��#19v�����dg��ӁT������C-�B�77L��O��5�=H� ����<��ŀn��U�YD�@,���3�������t�,�"�w8�F����k·��L{�7�(�o����6S�AZ3�ۢO2Y�.V*ɹ�xXYkQvF[3Jm���Q9{���N�~�Va1d�cs�pКp�1�7�� 5)jV�e�j����T��o�A:���XDj���8u^G�� �HE���j��F��>;U������%��@<�(�)&�	��#�D�t��A?�ӧ,����q^�"�1��/�q�Kl�I�r���*��@��n��O��(��d��"��Rm�����5���R�z{���m}?�D=�J����=wE��-V%�'�l�v@�d>4ܜfe����J�+�:Q��j��rE���� (�t��
�ca�yƼHy��/Ԝ1�H] N��}��bէdsC��&���j��6��Y�;�;�dbb���EP�{S4F���65Ux� o�Z��6.+.��y�z�Va��6r�m4v 	����/1�c@�1=�e[�RТeW�hV�(� ӄ��t��S�;��eI.`㿙�p�zK.YE��f���IE7XHʘm��K~X�h����:�� U]�4BLp� ,��cePM*��+_�|�e~�����D�"T�r�������:��g#���i�7��~s����g ���ZA��%2"�q�Gsa�b�z5��+el7�hGӄ~ߝ񄔺�_�3YM@���\�`�G#4'����	P�<bED�������	)WP�@�tBu�%����%��f���ń�C:� )b"�A�{B6���Qf-ݫ���K�h��Τ`��)=7M���㡿?"��%�1�C��	[��Js9���#'*d��<���q?`��C^4�@}]Zm�h�w�=��6����$��A�����

��m}���F5��,�l�N�Y�
�����ف]|�+�*��U�.
l}�AkI>_����?��Cs��\Hx{�m���3���q�`rS�>�7r�B� <�zW�a/@���󤳜�{-����3~)(��5o�B����ֻO�=4�rny�PgE ,�|ES���_ִ��t�����)�3K&��"�+=R��+�W"0��p6h3�F(0������c^ mJ�=u�Aϥ�/��V);:D9:�J��@@�.��W�7E��w���j�kՂ��-�ld{ڎ��\/��W��E!n����zuT��˭�m���J��]�;�m�)S<<���è�:g<ԭ���G_d��ȓ&�o
%T?c+8jc8�����5��v�Z�5s��A�1>!�KX��$%����X{PB���"��8�6��Ҕ8���4�$K�R�d��.�"$�:����$�����ϦXZꮣ�Ա��Te����44�a��0!4����G�8�;F�{�1�924��ɱy�C ��\1��ª�R�����	�>+�`�?%S���IM���e}�5:�'O2�F��X���=v�-���T�+Ξ�����m�� id$@��wM@��1�����1�zg�lS&�[�$2�	VuO��uw��D�r�ّ�Q��1e�چ��ì�E$�zR��0̼Ҵ{F��!�����
Y{�N�z�H�9@�TøJĚ�ķm�͈���,���y�Ӧ����lQ����%B*4B
W���`j�CDa∺��;2J�o,1����\Z��^���_b�1�қ��tҟsUEB��E�饏���q�jό~bI�ݗ[��e����g�7c�Ƕ��׃B�C���Z����z�:3�퉒iT`�0	Co�x�W�`0�ڂ�ײ��I�R e.�3���&���0�IGz&�JT�Ox���� �P;R�d���6��3V�[��S h%�?KľB_g||�� C�������kE�1�jl雚g���v9�JE�6��z�.�6A��#Pd�T�o�V4�]_���ż��(�Q����8�� ��vkAKO[O���I.c����Xp:,N�4T���	Pa���� �vI�L:�����<�^�����\�H�w�x��vW~U���n,������B����|ps�y��*�B�'$iַo�5"c�ZۯgJJ��Ed��t*����.�nT�~L��+�N�w�~���B�N�������U����7�\e�ƃw�$ko>��#ah�-5^����J�\���"��g<��mD���He�����D)�cʟ��_g�J?�J�R01�!����l�.W��=�s��t���nI�$�IM�"��[p��+�y����l����F'��9�����O�a����뢇�d���2M��2�9KBޟ8Q<T��<5����#�"\LgjD��,���&���L�oU[�i��r.��}�kh|>���|�L�F�/������͘�à3YEnAߖE�̹�*�
f�r �\���c[����&�?�P�_v@��D��HO�������WD�&��F~�dq<*�)�Ƈ��su	s-�}����d	�&E����3�/G�ۍ��V����ҽ�6x/9��p@�D���kKI�^�v'�a��h�����=�IET��4�`p�uJ)槗Ul-�U�X/��+�����5X;�\�����~�P�qhw�Q�%���!�H[;Zj5(��֓��(�{[oD����v������&����UX�����u(��QH[%L�[�/�iS��c�?K��g-+�&�Uc�i���6+j	�,8�ʴ�����3�g����7l��7�o��$	v�́�z��AB	aDq��?�����:9�w�����?��u3_EO��ē��Z@^(�$:v�	zR5�N C�Z���_�М1�]����8�4�/�i�Kdՠ����w^J�zt�LJ��r�{4�����&O�v� �vǇ>[���sW����	�XJ�D���	�����D�w�<y&�"���3�mP�}� 筣�ͺ3L�<�O�l<'k	�]jsX�͔�y57䪣m7��\����c�7�?,a`FPW=�y�<�˩sׯ��ۘS_,�����8Ui����6�!���8g����� �a2�6��v�P����[����\�:�t��(qJ �9�������Ӵ�X�ܿA���`'�=����!����'ѻ��]/}������9��������D\C�ȅ]/�z�OB$�j;��WVp`Z��o�vy��A�MiT��۲�(`'��!�}[(���XUo�,ʡe���}�b#~�Y��E9��-I����h�Su�jl� ���Ӡ�7�#�b�Ă�s�]/ie:����p��*��}Ja��R���]��M;9dʸ��?���4�΃�U��St"�9�y_����R ��M3��#>\bJ7�Eّ�u��ʢ
O�|^�� �/���whRP6����>��#s����G`��;KJxXc�ef�7�pF�Kr����ŷpm��+�~z<��Կ�^lI�`<�z�1�l1$�]��{c�,��J��H��epZ��iT�n�7����{5\��(���Qy����Ü���d���;�J��p ���ޅg�m?ę�� ���)8�"��Y\��Gg7eT�9�$�2�c*�HPc��X�`�+�o �6v&�Ħe��Y�7���@�|���t:�r5�u k]��֒ی$c��tp
2��XJ�ʓ��Syw� ���� j�4G+������kƩ�Y၏���̏#ղG5���asN�W�K� ��ԩF�ːoI�$���'� �v���	n�EvʟC_����{��y��dO�9�B��J���b���E�8�)?V�����ޟ��p�Q#[uHX�u�6�"����N��Fx�%���ސ��~�[�4��EB�q�vsf:��5-�#��c��}���)��uA�!-� B�i�Jzx��50b]���O� �2��l�Is(�p�MZ�±�[�n-.��O8���i��? +E[?n���3�ZS�	f���t͢s����Σ����Ѐ�j�ϷWOY�!�~����~1;[��h*��-��9��D�����y+�9M[�F`��f�4`��wk鸗�}�w�u��_!���xi�����rzG�i5�{�>h�i��Y�;p�^�{.h��pI M��%NJ�L�@Ϊ��^x�cv��,_i<%](������Z4�a,{�I9č[���yUi��&�J`ye��J�\���(���*�n����ΟV�]�n�`�1V2"8o�1���H�95ҋ��������F��m~Z��K���P�Q#�nTю�QVo�Q�L��� �rvG��bl�c�"c��6?;T�`��+9tt�wC]V��O�[,|���Dn��s}[K�����Y��*l��g�!эA��Ҧ�/lk�=ƪ�뷧�߄����B�@vg�I��)��> J�ߺ
�!��Ej���+�u��fu�;��6^W�B��sI�d\�ZL�t��N>U~�	vP�d
��V	�Iӛ��F^��`�wWf�}@�+j���r�1y��Wg{z;L�KQ��7�6��?�*%�k��S{S0J>U�q����/L�}��ԯoCb�C�#jP*l����NhC�&�&�o&��t�yA�wc���͎�/�蓖\k�Е�`���	ׇg�q�|��b^7��+F+u�_"�t�����;�3�qJ�� ����3?lL;������ʦ�p�� ~����܆�?���	��<���ҫ��@�A&�[P�*O�|�q㦥@�+]�~R��Ӽ LF����_"6I�����E����3����o�D}����.}Q�9�Zp���7���]FII����Y�A�uĉ�l1`�00�[UYQ�4]���ڋ��<�38�+d(l��IsuJ��26��q%�hI5��m�h/��g��F:+>�o8�w��ƚ(�ؽ]F[-�T�7�	 g�5>V�Y�lTf'P�����؟9��e�R¼Ռ��8�EZ��o�=/�)&*�g-�-������,u~$\C�x�<N�8g���Wߐ��@ oY0&١i>tT�0�sw�	��ᴖ� �+��!�X�3��aP�q���RLL���t�c�\?bE����D���4�]�ױ��%Ciռ\i��\�Bq��R��"m$��@%�4bD~�9H�Ɵ�� �:������Y�IcLuz�I9K��|G�<D�>�}⏜�SF9�%^b�%�,0W����l�%K���
���X�����L�Y�@���Q��I��K�C�����l�P�5K���gE���q��  ���~�D�8��)�̚ڐ��j���"���S�'L�D�r+�f��$3��S�$�:�.[�$�:T$�i3�
Uu.m��OK���T�������;֨X� ������
�RӏK���O;�r��胣�Nh9%`�Qe<�����g[��Sv"��Fq��["�t_���	��W��W4/�W�p=�rۤ��%"�F�Og��G�`+��Ek�@�����6i���[֋�7i�4O|�����c1[�V�h9�u.|"��
W_d|��јb��i� S� ��B�X��b�ȸ�|��]����f��0[�G�6�hbŮ:�5c�gP�f�gU[���Z9�7���Ԍ��%PQL��P,�3��J~��� ��zjR����M�ba�l�j�i��^zL�L��J���ӏ�e]R�$����U"]AyI�}�n٘
�/ҹa:V�v>���p~�t ��L�q�,M��?�b�|�G0�ob����l3��"�AZ]�3�LQ� Κ�����CȎ��]BQX�o�C����!]����Q�r�0؈�4Ӊ��ώF�C�Z�o�m[��dAe=&��E��L+n� Q��"�\�d�zm-h1J���VK?��iv�s�^#De�J9��d�8��KNxY�0O�D�(h�����)�QRi7 ����|n�`�{���1OY<��m�V;Y!���'̤�17���N��.#�'��T�<S�Va~����X�&6���t�������nEc�)(�	��X�wЍ``T��`V�x�$/�]��ӈ�V��V��2d�=�+D�z��H�h�`�j�`|�N,^�fr�oiV�Ŗ�%5����T�'X��7���g�����M��s8�]-�G�)n��~u�=��KӮr&�-V,q��D3��AU�d��H{����`��=AX����=W��R��(V��;� &uuG��:N�&kܴ�sH `�A�
��-��}z[��BrQyOvFߐf�p��0aDľ�ſ�ɣ��$�`�!:�Á6�Ьz�7U���(G�D��i�G��;y�P��8X	��W�!-��Q��G��y��i�Yd)��l_��U�@5��M
�̢�{z�T`J���D����d�]P�L�.'e8ӏ��S,T�y�(;r�r�����}S�03��%�c� �\z�|��I��Y�XN������H��Ӥr�+2[�����H������C�������\d��(��.zb���vB���h����j�7���XMк�y���h��7�Baɮz����G���fһ�<�(�&�z	 �o�@bm	����׍����g�k0�|\ʀ~���U��o�{�䨁�p�5+k��K�3��c�o�eb8�خ/����,���l�Ʀ����{Q���衧b�>Åi4' &���(�-z��a�VЁ��|���lT�A�^=�]�(��H�(m���XEz�.�YG��_>d���Zk$����q<�hko����[UN�<j�V�SK������yUܢ*��+����$V�҆�Jy��|Y��� H-��*�#��XKOwt�9�e�W�G�NfÌ/J�6�=��O�Į������l\�"�bi����E����Cm����	!�^T�D����e�b��ٺ;����><R>�!�Y�Zx���|n��r$<�µ�����E��?hyO��E-��$㓵3܄%�~�V�9<�����!�)�ՎĔ��v��LҔ.����_��l�,�^���F�R'"��ݰ�W��j{p���ݢ�'q��0���#����"���VӀ3��gdۦTc8j�o�fx;q�&�����)��gOj���
�9�/���L���X��}�j~�mU���Ml{���Ő��_[�|��_RJ���N�.���V��T}"�M�i^��8낐��ߙ���IE�=s)�0H��/��~tnE�K�G�����}�G��-�D�|��g��h�
 | ��'Z���3�������@��%,�bU�F��3�6�:V�9O�3x�v'���#����N>WHA���7g���[^����9PB[.of��*��$���%^F_�y%b9��oh���ڝ��Tz�c0���7� _���j��0����Į�go�Ǭ�G�\�B����������W�
���Ub����r�S�!��e{hW X���$x�9*bD� ����l9#T�wڙ4Y�����Z����Hwh Om�_[�F�\r�҃�X�Uy�H���R��aO����9�^lf�1nFn����q����B��������)�R[��T�����F���ySIl��?��}w�I�p�#���#%�/�%��YE��{�Q��}w�̦�Kx1<�6�@y�������k)wH�C�j�ޏ��Dh��.�֓�;+�I4VO�	���w|N�=|��>O�F�bu����#��p�n1l��i��Nd;��V?q��+1X�Cz�j����&�W͵���1��x�]b��r*�6�	��"�?��~��gK�q%�x9igG}��7�7D�4�1��	���8��hy�r����57�H�Mc7��� `/�T�Y����`o��|{Z�}��R!�j�glŏ��I�n=�*P�6��F�T� �Ԍu���g�����Aؼ� ��8[�Q
�% �i"�-t�ؠ��b�TUr��!�8ܤ/=;��ʌ<��~����f2�I�'A��-w8p����s "��Ic&Z�oT���:U��;��㈂u4�$[��:��D�k�<S�)UAθy���^ �m���i~�5���$�.�ٌ#~��va܋\�}�˸c-6�Ux�[�1�a������Z:S<��nh%A�j���~t�?*�]�2�Xw�9����d��P�Ow)k��K��}߄Jm^Rg7�2�c���Yf�"����`� _g�
5�(�{�����$�W�HV���;���2g&pL����7�A�ˉ��w����J�x�]K%e��p�0�%����~;, `��^&�Q{����7�uBߋ.�Hq�#����~����e޵��JS��6���cyD0Ȏ��sG��B�:�i�A��S(8h�p;�uU�+u��|���Π�luD�+���3���aS����*����"�����)�����2Nf�۵c�3Ӡ��o�t�����
"�۰ѵ���������߶zޏW+�d�i�y,�V����I�W�{Mɦ��STd.�k�5��f���Z��.��H�:�&�)[S��iams��	P}�Aӹs�q�#KEவ�Sn��Du���]4욈��9^�u�:��J�t�������Z���-eq�I�B�	q q �+K�hڲ�9e��-_�-,	 M�Г��O8fp̓B��q�TNd޹W����d��Cl�M���V`�ﾜ��]������Z�H߲��˧��ت����0���5q��01�Rխ:&?l���D�6yƓ�y�V�"vxv���%��HC2�,Ș�7��gh}q�5{2�$)��}M	�-5�Ș�@���h��&��2��_��A�_1qiw��0�aVq�� ��"���/�I!��%�r��	yZi:A���Iuie�U��<W�0L����%+1!�?9��B�Ώ�ɮ�����W���D�ǅ��c�^���^�|V!d/v��B+����F�������f�:/��!��@�Să%ě��%]!���`��&�/�&Z 5��kS�U ����(�c�[�;�S&Ca(x��Z�(T��Fb������u�Ţ9*���\�4��2!�'B�p$3�� >�8�_�qT\&��o���{o�����}�L�^rGEn��ƪ�NU����l�c]�kv q�(�Qa�T��ybS�V\�0h�����x0W�4K�5'/��Y�=�&�9�Z@��5��� Q�z�5c.~�=�-�0�~�e8����>w�Y�4��\�&9�@�ph���PitS���-'�����hF��}���H�{������˄�43i�&�ͥhʝf;�性�2��T�F��X��d��I�p����^;�����@��z�ݹ��O��\O ���ֻ�1;��!��e�a6��f�>��m�~�q�@뛔i	K�v��衇�mXT�֧�h�aP�#�dEP'����k}^�n��XR��,����MH���Γ�1e?;�EE �n4T�'��_0�~�oR�������Na����K�P���B��<ħ1	������"��NeS��9&s�h�F�\,����wJti[f ;h�
��W�����������>�K�����N��Ԋ���A����:F:�i��F�Y���1�砨x��$S��֞�t����p��I�=|۾�ԒL�ir�6��[�b݊����Ğ_���!(;l�^o�~J��+֣�§+J�k�G�Uuw��,C�� �Hз��*1�L��f���Xh���)B�����Q�����j��,S��<�*���,l��Z�(����H}�������Z��,�W��큣.���h��'��چD��pa�����+9ñ�&�!lͩևEߛ��&�X�[|��y*�Q�ɒ��ڪs��%��l�&����u�k��k�,%�I�5�kx�\��R�}�#���7���ŵ�b x�?Y�TyT"�қ3���W���\�u`��MyzB���O�>Xk�ا�Ri�̨|sB� M��짪�����JS����=sK��,Q��C���W��Y�a|:Yt���UA���5���*�֖L��>>�n�A���A>��<�m�Y�T�	,I8� �A��R��:����������G�(���8��e�'�xmsA{�N�6�������`)�]�F��=/Ah(M�������:%����'���h˯�Qp�8�i���51��~��^i�4#�����l;�ߚ���uUߤ#��������v5:?i��ML�e\��O�����L|�j��L���{?F�¼�"�3�8�3Q�))>��Į�$�/lFvES���=��'�Њ��%;�L4חf�� ��6?b7=�c,L���2���
�¢wb�����K(>oP��{Cl;M��8�K�r8�W;}�aZ�`f3�\���s�Ʒuʳ��U��:<�Xhv>ؐ��TF^AT��"����_9���-�1iw�qk-U7��nć��J��6)9$�Br���9�S�1����==�~)��b]����.x��V�c�/��Ios-Ʀ�^"�F��6�-n�a���Y����x@��:�7��O��g���oo/��z�J*������嬊JNn��(��{�ǁ���K���@>����D�p�2�Ζ+&Z�X�L(� i��u�U]��ϻ]=^L���=;�z?��X$�����p,:���F?;�����q�÷�C&쏞�v=���8�ܛ�?s|bq�h�=����s+z~��^���a������:��=�[siJ*W��YԟWt�@'XL�^�,�	x�4��;a�+lwNY�?�a̯�!BvP����ꀼ]�#-	�-+	��aa��< E���a���,�3v�@��[��Y�3�Y}`j��_�O.>Z��f~�����A\o����n���<���b�f���O,*"�r��>:=�F�n���9�!D�)v�bQ/�%�Z~Wl7k��c��Op��s���^}|�b9�7��q���+MJU�`<զ����O����1���jx�痞/3�M������@W��k�e[����7n4MfƤNH򥔉c�k���D�A�^��r��UQ��X�O��wO`3��d��gv��p�8t�m�bͿ�HqN<;ɝ&IU*�[�U˗M`���TN3g��r��o ��T퀼;	��ThN�O*�Æ� �<�)օg���&6�9Vw�99;��4�f�2ո�D�5:�:���<Ԅ2fUυ�[�*�
J�ӳ��q��3��I��a��z�'23[>u�W�ޚi˰2�5Q:�p�1��=ս|�l��k')���ĕe��b �����m(���V�VM���;�� 	��i�^Fk��"���z�!A��0��h�Ni`q��"��+<��yUL��Y�_�9�`ES�y��oO�#��'�[����>��߂c!cC����o�
:�x>q�=419k�_#�W�pQ��WA�����UAZ"�t���"@��o#X����up���x;a����P�,�����M:��/���i�- ��퐓M'��9eql6�����x�$��V0�r�!��S=���T��+��c'D�wR����������\G�>��y���S�z�EF�,5떬��h��Ԡ��� �=��&�e�_�to�����o -ة��,T��C���������/G:T�17���|�	���G�ea#b�FX*��m�&=� ���6�k=h��-0�˜CkL3/��x��@��1n�&M�C<ί6ߋ8����o:��FC{�1;��ѥ�5	�� Xigz��K�A ;Ю'��	�����`~�m�>�F�������~��Y?�g�O)4}�"���<oI�P�zNí�!{8D�jQƧe%ܪ핳b�Koz�VG}�Q(w�XĚ��=�ݷݟϼpE�8NRPH{�H�/l�(-mO�o���hB!�l�Z��Q=a�n�V<jyА�Fw�"`6/`�(q"�k }��m��m����i����?��͢�]�m�HS���\�A�^P�͹�禐�?4���;�9��^�.b~&-wT�O��!(I\e)��˄/W�i~rC�n}��w�iQ�M��8�IVsr�I�!X"!1��{�(oA����ZE˿L�4u\Qht��2�!��	�P�0g���SRl�҈,/_�,�c��Sǩr��;�)t1������xE��6���;6"�ÇCʾ�wp�ڎ�6�3�U��������;l,<�Ɵ�thH����2�A:�	��@�+� RP$�ι l�����z�ľ/��z�uR 7�����`pM|�}\(�U�b�.�\5����U"dZ#g�t��U�F�p�ۜ�#���cr�;Lu@%���K�ZZr�1��:߄��b��X�|>�����`!����L/�e��E��;�s�U]n1��U�^p��U����(���iX��&���(�I�
�u��&�K�c�>@��Vh�s��=
Z�����ҋ$�����+۴���:3Q\%��&��X�z
��@Au����N��Y"j�b�xO�Bj��`0� �.ƭq�W(;x"Cɮ�Fq�Nd��i����rR/oD�J��u�$��ANQ���T}X_�J	=��&�j� Z60AΌH�K���T��L�q����$,��p?���L&����m-XE�t�*[=�Etѻ#Q>���$��}���i�9��:�eN/�h�\��"~E.-G�*MJC����f�=@��]R�5[Ԃ�D��]�t��*4�屾����P"��!�h��k��������yM��=����rӕ�x��ln]�v��Ĵ3ssox�,��1>�;	��mV����K7�Lu�FAg��IuZ������1��Y�4��H5u�*ZM�m�YV �X5[���  ��~ Ѵ/ ��'���);�z��=��9 ������B�w���������/%%�0KtV$���7��5�h���\:.�*������g�ꋀ�~�  �����闈�9���?֖��Q�D�ةF�&�f	t�����\7�~��؁��ٜ+k�Q,��T.��ٶ}�7k>���C�Cݼ�e ����'D�}Pw�B;�Υ�w{�-xJ�kM �M����{ΒJ��s}yݝ� �n>�O}+.tl0��z�"{E�/b���{�1�+/��2w�d�&�Gh:����g��˨��/+6h1�Ka�lD_�3�Qi^�u��	R�B��2?��%Q�����F��>�f�ʬ
��H���~��ȗ]�i���5�q�KM}/:�5B�{�#�*�i�5ɻױ��V��tԡ�[���YYxo$n0��5�V@�	��꿆��ݓq�וּI�����d���]��^�\��2&�� G�S�y���U���i��決�>�x왺Ndy�S���nr���⾌����K�E��-^��b��"��^���Π�ʦT��r������|H�O^�)5[5sM]��AEE��>4���m?(�@Ũ�p[�	�b�T�Rv�K��4�a}�"؞㤬˭����A��ʿ!�0�_�{];��`��� 6�=NHJƵ�xs�R{��AO�#fj�����:�*GfǸ&����T����e>3i?ul�O�U��q�_}f-'�:��ts;=�k��sqԷ�ʧ~�������}�YHW˕�(�]�b_Ň�9 ��M�WO>�����o0��Zg��G�6Ap�����ͩ7,&O���y��?�J�mt��#��QBh��-_0�#�H�ھ�3O"i�5+�.���C�a�GV�Vѝ^��`�vUHɾ�0=�\х[�wF�t�Я��M&����=픫���O�aN�J����V��ZsL�o_KD'�[�� ��O�� �N,�'AM�Zủ��G�O�C�0�;T���+�sC4�Co��z���8�v�`&�7���6h������R8�b���K5lJ�N��ͩ�b�q��)ʷmIb�ɻ�G��[��y�&)p����>���5	���ְ�)D	4�����.�&+i����ĩn�@���L�?�F�a�/�ND��:�LE���L��j?'��e���"���}{_h�A=~9=�MM� IyT��;}s�Q?�3TdD��^|';KH��(Z��*C�d�$�i� Dق�P^@�@&ݟJ7a	���~���ڐs���qU�mn8��X���g��D�rm��.��.^Ȥ"�d�$���u�"��:i�R�X�Ϥ���2�ԍ��n��:�ȟm���Ɵy�%ХE�q�FTc֩쯝O�Pm;9k���Y$�����k�#GM������;��y]����>ΰ�?U<�ɞ+����ϡ���~�]��<����]#^��[?\K[HۻvXN�P�c��ѫ�ΟcGo�/H�(��HڬV9$�Ep�"ܯ���ÿ�GE�b["S[���"T���ҙ�:VmH�Q�`�p�j9�am�e
�QX�`�^?O��Q�
���(�q0��ۻ�u���|JJ? j����@�S5 %UZ�5Q�#�M������|r^���7~Ϲ�ֈ�u���ṥn?sW�n��9��r��[��8��Fw;�t>�Jv�7/���߽���,%�Ѝ����?�ˌ�${xl<\2���߆4gU�q��!�
�>`Ai��f�����'F@{ѵ��m�i����I�pg��?#>'��y�0�0F���I@�j��̣.5r���;T��^#�`s��.�nw��M�`@�g�gD"�Q��r�HH�/��m,,iA0@j�kϖ�z��,<q^~��>��=�Gq^�"יb᫨ϳ�b������	��AeL�Eㆼ��&�y�_͆�_�(#�rݩ������<���E�pf�6EV|����Ϳ����~ ��i&��>����ma�!�|�F�^��<R��V^L��2I.x)U(
��"���:�lt�<���+���4ҊḂA�_G>c��9#K.-�ɋkջ�ݩX�R~�hض�ĎHy^� ���{��\�&T�v�ԗ� 3��+�˟!���|B�-��w���?G�_�@f�2�N@��~��ļ�^N���f0����P�DZrˑ�"NIS��aӢ���VJ�����q��d�uՍ˺��r.qbn����P�s�>"x*����Ye���A�lD��k«7](
]��$��}�OWWr	�����oز&5f>�Aa���J/��u��L��v&�RYf�9��\ֶ���fN!�C�^���|�f�USDv�P�y�ٖ�eW������襆"�>љ*�W�j7Nt!�XR�أO��D����3�@�8��~q=��z����MT#l�_M��
��m	����:��A��1�9X����O�~${�)���Y��%�ૹ��S�\��80��5���%���g���}��b<{�7�2�$FNE|.�a�I�k���IXU��j�&}8��s!^�q.9O�6���o�P|M�tP���׷�^����hj��9=y���>�O�%�����BR��֥���Њ��	p�.d`,��"��7'N��xJ�Q�r�����hO�o�q4aؽ^��s������i/+��Nmu˴c<:H|��DxO��B�YTtK�t��J��ukqkl�:�����5���HQ��(��^6v����ii.������'�dI>쌗����4�_�NYL>��Ӻ_m��%"��i!�G5|M�bWAi��D��(s'Mdzef��Hl�[�B���fm����)�Mf��j�F�LtuÁe:c��n�
�!�c��'�~��~�s���Vd�8����l�,� ��6�F�����|�0 
+ЭO�`��FX׬^�%�w9��2��UhT5^_QN{���8N�>���8%(}&L��j:ㅧ�n>�E2�Zw{���p�^���� ��m=S�x3咟�N�Q!2���+P��%{���l*ʏ��*>�!�L�7['jĬ���[ֳ\���#)YC�z��.�T����D�F���.��H@�i���2\�`�^-���^�*��9)bR