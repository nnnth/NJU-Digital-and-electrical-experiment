��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�8�&����b�B�
���:w���w'y�GO���w=���Ȫ)K��S��.�5��Qo�.v����I��D'��El����4�@���P�RG�ERC������(��_���Iv�{���E�.wc�����x=a���v-Wv2zo���	��)B��|�P-���ɺC@B�'#iU�Rx�k&��A����T�-����@ه:ɳ�@� (���#����?�ڎ���y@�`t�f�KzV��Q3�@��ʒA�f�ĳ��Gz�uؤ�!��2�j���\�$QF�18��!w�-��o&X�]����\͒���%�]���I�4�w7ٽ�k$�?	(o���M�U���"Sj��3 d�w/ ���pu;�sA�t��p�0]�.���ʷj�(��z�����Fo'�R�y=O�������A�!OR��=���&��H3�$٠�PU16�[h�c�ꉲ)�F!��_x��|�+Γ;�$:���%���R�)&��~)@��u A�?�'S�C]��o��Z��>�x^��!M����?X��2Et(C�<�Ys�?�(�4�5օ� ��H���&�p��J�'siRp�kTzY%�o%e��Σ��ښ�"p������e�w��2#_5Ua`��7�1��������*}�cJ5K�˯����&x���4��k�<���3w��_�Ѷ߼/Q�����4`�Z����Y�U'͞("��nU�������f��?2��0?ӛ�H!b݆��_=,�K���$�:����=��4��s���c��0��#?9��wB��.QPxVu�mD G����,w'�$�	�������p����"��2ܻ2s�A�H��;�mw;�?���tH��u�!��ώm�uc�
��a7!P"a�Xn����o�h<%}O���n����%��TH1���x�t�(э�x�頢V�:�ݽ?�&�L�T�0��R��J�� �\��/pա�e	���T���	����)	��|y�2,�a{�j��B ή�N'�`�!�l���Q�݊�U���RȺ�'�-"�kh'�j��?N�T٬e��>�}�S��p��,�8pQ��}�9�2�ȩؕ{��K?�A�������\���m�0y�����n��bX(M�=�x��� 4xB3_�].f$� �=��[����)o��6ĭ�B_
����op�DB���Þ}a�`0&���ɛ���Eu���V�0��uY�Lۯ]K$B�xr̭"���"f��MĽ6Y1��ʉ��7�Yc���fq�������1`������^
'��I,R�^N���ͭ�S���f�u���$��I�s������1.j]I0��D�5�������iΠ�4�7[3�O����u��8�^s��	}!�p�������N�lD���̈n��ԕ[q�r� GZ�T	B��1Z�#2e!ǟ`_'.������CpHy|�j@w����X��Q欏�cO���E?�=lH��zOl�f���Fs)0�q*��@"���\FŃ�,�	�倷�n�V�/�/E�h�V�:=���r+V�L�)(YܙYv���gSm6��6���s����n�mO�'O�;���G-�ɇ6
Y^>sA�f3��S����j��V��H�G/tJ/Y��c�S����c�I=Y��`K�"��֣���
6�.&�w�e��'W�1�A�#��+O��5Z)<1���
ե������}����V(����R=v�A`�Ozh�[(y����YR�'�C�K0dxS{��H���I��N�T�!��=cV�=� �B^PK
&��*�٥�)O�!��RXA�P������GKS�E"�j��� ���@� ���S}�s��F6n�J[�	:�=(8���+�����ܪѵ	
n�F���8S���XUC�5u8E�-�iZs��ue�JyEp�&�����"ɏ��²�<Y���i�Z�[ԅ;��	k��A
��#�{�5�7��!��k��|��M��E8�2�I+Lb�t�W݁��!ɏ/�;��_^!�~��ᓏ�
*u���"&{J5�v؋�0E���;X~��O�R�2�(I?as�[�m~�b�!<+�ۆ��I�9Z�<�w����(l���/�~?�ÁȈ�R(I���n]	N�>y� ��_�sn�v�,���?�_��c��B�1p��R°!P�ց߻R���_9����Q��������s�S<U*�6������t��%��Q��!իŽcA{y'zOr�Wx���;���[�fr`e�jHN�&h�[\T|�BlG�e�C���΃����̍SH��F�����ݽ[+�_��>�R� �x,�4�4C����:<���Yc���bJ��G�)�w�����PB���VQ�)��� yY�G���0�V%�9m���Qr���� ��	N�Q�uj�{!]�4���(��bg���J�p�p��_BjqAA�pL�qo��Φ���8�f!~w^Bt�]0����ߗ]Ζ��{۹�BojM1��r\O*�]��{�OY#�8�.�t��Tܝ�壛m
�e�L�%�(��J�;nh-�e���ӈbn�ǣgY�J�%^�<o��e��2�4��=H(��M�V
&X��W�!��9�5�'��ٟǬ5�\CTeu�x���s�TlF�j���"�;�!]��f����c�;Ѯ:8��M|9_�M9J�Q)3{\�H�|o��\�� ﺭA�{:�-᭥����).&�1�,~�����_�^����l��~���6Sy�@��lA�̬e��Ո�.&F-�'0��l���/��u��G9�n�!�4K��h�9�1SR��	�m,ￏD�PO0GzoF���^��_���i�X@؛�Ɋ�{v�+X*��#L	g�@D���\���E����1mC��#�*{�Π���,8A�U��aؿl"�L0�ش�iI��J�9�]f[���ktB�Eh,]Q���*��M�P���xk�����튌�d}�)!���:o�<�*� 4%Np@u������~�7��|�n�ӻ
E��_�!�L��[@�wx�Lo�?�;wx�k�YB��H3B�A�8_`Eep�D��s��$wz��z:r�*c?�4����{]�+}�밎���u��D�*��k%�<��ad1-}ŊI����I��2Ä."ӆ�j(�[��]�8o:���Ɵ�Wkwr���J��.ӊ�s�m��*��d�"uaI��D�mGPw[�M�H����S�����4���MfoK�Αc"���|��:��b,R?�r�����0��'svw�8.�R�©��%���F׺r��Pc~��a3R����'zI9�Keh���t�&�F��a`Ua�����d���Xl8�
��c�J8H*��2���,ļD?n=�:����E��R�zZ!��A���f����g4��<�!"� ���KΘ��&|v�9�OB������id�hs.��m$?���2tP�|-� vcvX%�q���[��L�~x��c )Ok�Y&D"y����:`k�6��`�;m�̭�	�N�U��酜u�n�q"��ֈ�iYD�uD3H���A�)1|C�R�ð���Z'�3Q}�Xq�^"�6՞�4�r3�c�E����]�8C�����Sm���l
�48v7�k�[#qEh�KD�b�o9����h'�*s�AggF��@��,mqƈ�3wz��+.�N����8�~�R��R-Uʸ��� �g�@��\�T(�;��ה'�Ɠ����}I�bv�
I/�*T���-���o$��������B���F/{c�5u+�����3�b�'��L�����Օ �����
�Ҵ{���Zvk�fST�,˚�F�݈�'�Ώ�J�K���:�xv��z?Ι���_:?�@��m�>�K���'í=�'��-�����&+��/��9�1p�vb����D���-��:�S-��RHrp�7��ieU]���}����`g�#���@��n4�ϵW0u|��!Q)�G���\��� �0�R�y���M����q�n�%���g=�٫��4'%�j�D��tm�@E�)nc�Q+��7�#M,	r����i+������o�����������|�܁g��S�v0�5�'^��Ml�\��7�۷
[0���`���<c��D�OҰ+/g�RPB3l���B$������ ������o�9X��O�ε��Ӆ�� ��朽�U�N>>�Q�������t��v���d���6"���=
P�/</K;�G�A_�� �v*�d��Y�Q[�b]"�����3�8!l
�?��F��Ж�	��zQ�$e#
"̗�یG`]�g�E����v&$-�s3��Uc����z-n�&㇟D�5�ɞ����3�Ο\O?�! ��Ȣ
��8��l���)�D��o� 1���_�I�J�,P�7��bx帿�W�"��S�ɌOz�%�I>����X��BOM��^� 
�C��-ق�sq[=B�l�aꓱ����$�.�'�*�`�4��(�3��%�aO0�S�l���&@��l��(�p��za&��EI�|;��x�vY(��i�y�>o�lSA����X���g� r� ��<���R�O� ���\�׍M��ח�p�����SGYi�^�tmbP�F	h�Tx�&_{Y ܸ����3�2�<8(Q�x>����R��KX��N��\q=�)���Y��Ѡ�^�h��^�	;2�m�}�H�,�屛h�\R� �S�M7�����tu�ږj� �p4����T����c#p�]�]�#�����n�����K+;���X)����W��6���3>���,h�����=����`Dwb��A\q뇘Rc�dI�:>_J�k9�a�jF�I�{��D����{=ĳ��Á�qN�h!|��SQ-�-�i��u�JC�e�"�H�Y$r>�����њ�Sy�^ڛ��#sw�iiA�8�8#�D�%U��D^�:i,2��`�`9]A��go�~�U2���cv	�I�� /���RS��16uؔ�5�B1@:ϸ�5�D%c�'KT��$���A�ψ��>6���uںm|ۼ𐙶 �P���>Y[�0�7���U��[��
7�O�~3���! e��}]{EYn)�⺓�Y,s��5� l}'}hٟT〪D�>{c��|�8�ᙀ�u��eR���;��#lU���cI5��bַ����,�=��)�>�̅e�EH�KC�<�������2�Ս,F=�K*	���p���^�Q�pe.� zڕ���
F���k�m��#O\2&P���sG�?i�&`�7v��A������/�Ι�(�J�ٙ����$p �������'�w�~%��,��K_`��f<�,���.����Npw-��\���n�S�I�o��NU2J�LH���b�5�4O�W9ʜ2���f���b��ܛd�	ɧ�?�� �	8���j�WI�KU�hɅ9����6%�������Q�؊x� �{�b���h����S�ܵ�>Su�����;k�zԽ�D�&�0���PJ�J$}s�8H���Sʑ�B������f?5$Ək�-͞��s��~%�o�0~9�ڸΛ7$�sƩ=�y`{�i3�Pϱ6[���RQ:� Zz����&PX[^r��-t�p�:\ZѮ�DX�%�D?V�;�I�+��F.S5�b�B�_����Fg�*�"3(���cl7�a=�m�S�,����4s��9��>�Č�='�!��^��oL���.��5�(�S��`ţ=i����ټ�"��&׀�Б�-��E��bAx��V����7-�x�}RV&�q>L���4o�"y�A��[�y�H�U�r�`sŧFU�9R��W椩���ypP�52�����>��c1EiqA)C7\o�F�n��^������qǲNFI��6%G�mۍ�֠v��C��k�Ƃ�zp����$��^f*�E�i^$�*���Q9�t��5ɠ�ˑ��ٙV�lm�L�/CK�Y	�I���/��J�����J<��������:�� ��J-F"��DiDjE��ə���I/�JK�0�0l�$�tH�k����щQ�eqo�ُ��s/;p���&�ޕ�� �"�A�˾ҽ1�����REZ��
���q):�'E�hm#T��e]C�#�	��@�|�ٚ��ЀRPN$����|��M�z�dr��E��N���T[�����cf� �j��E�ґ�2I���\��LP^�����Fb�|�/��$���`�ހM�a�P�Lʗz�ym�sB��s�rdG�z�1xh)!l��L_Tj�"Ic]�}_��]�Af?�4
n��ɤ;�Ls�/��o
��-5�%�0x��7;ޞt��ځ�Zq�4��>�����9��7�5��R�t:PY��r����p^@�D��![��9��QFQ�^#}t�����_G1qҵ(�4ɦ���7��;�T�
�����_\�Ge�(�ja�,��S��ֶ-��>Մ0޾�+�i��)a"�6�U�"r���cc���%˟�q ��܊�m�]P!6��$���>Ut��Y��8�O��D-&����=gmv���E۶�Ӹ����'M��7;�J��Q����#����>�B|. �E?������|˖�>}��뱌V�M�(J���J*�嚚$���$p�|��`oL�y'�1��G<�[Z+��'o���C����L��T����Q�Mp����Ғ�[{�C�j(�|�����eU0�/Wl�i䥴���(�T)�k"�e��z��
Î�҅;4*��v~r��%zp'������ZD1h9/1}|��K��!�;v������Ϟ,"�~����[�i�������a���:���QәR/%[VG��1���I�<��P����I���+�+8'i������Â��իzʧ�
~��q�S�����oM�ʟ�w$�r��%
�9��ᢲR{&v%8��v_�g4�.��j���w�>�x~'�n �Lj�K���t�q+kL�������Û���ֲ[]�K+��� i���~��7)ɍ���}��	sc�a!�|KD�?[��:,u~���33�UYQ��+W�ӟt��&-��Mۆ�o��q�Cv�WvG���j�.���<0�r�6���;#��C{��Ǎ���L���t<��d��U��9�A}w�� x)��eY���ur��܆Q�w���[���;�׃���g�:��/�> )��1�;Q7���!GT5���5W2!���=$��9�M��\�/��Mw뀋���D�B��s-(�I�<g���=�G<��N�?�69Z�Ϫ7Fs�Kݤ�-�~}F� ����C��� ���6�� �Z�C8Ip�9#��so��;*xř����4�Dk�7�J��}ep��L�$ߠ����8��&����@�ɢ��?��7�Z�/t�6�o�1)ЫEP�o���6�>.6�XV]� �'a1zN�R�VS`>Ѻ�CQ�t5]��[^͞�s�eE�M�16m�o�	��`]�}��)1Ӷ��Y�:�[��
T���P�!M��[^�4<����8Sa$k<g��'���1��U������P�����s
��RóAy��
��|@�A}����M|q	�S�5��}�Q>�K�A�PֆjLp4�mp�V�j�P��+a�$�7,f#hx��.%�3x�w���o�-�OC`sY���Iy^͙C��/������������.���7z0����I<f��F���