��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t؍�^��F��X�9�i�uV�$3���
�F��ɡ�	zU�
u��oJ��e��K1.h���K��O+�+J���,o�(w/,�͈w�	>@��O�,�� =Nڊs�FR�o�?Х��I�˻P3?��bd�V9֭>�u�<G��;Ey���I�B���b>-[�����W,�h��yMH��6�p\�)�t=��E�.�	��/�8�����_�x���c}�wo������ό>e���5KH�~�z��OW�A�o]��3��\�*��U�Et=3���p�Ұز�~�q޾R��nI��^����2~��Do�����ѐu���K	�����^}�Zj��>���ܹ�Z�
Yr�fR�<%)Cr�h��=�j=z*�v�p2���ܣ��))�tl��!G+'ʍ�oH��
C�*�{A*�a��R��97%S�ٮ������\����U��#��c�w�:���F@؟�u�yנ����n�n"wJ�3)D��pD@��w	/<i��o0�z���5PPY�4碁�W�Aj���7��t6����h�nSrsX�Kk�]1�j��E+Y����+ʃ�lO�F10ɒ�.�)ge�x�A�lW����8.�0���\u�G� .�E���wZ��L�_:x��&-�@R��`�t�Q���?'���,C8����~3fn��v��ۄ�^�s؍p�?��u�d�B��t0a�ڐ�kP�[� �ȭ�����f06��ϔ9�(�$�k)3ҟ��m�^2���N�0�_��V����Ƨ	݇~@N>1�^9��Z��n��s�O�>_��l'w�5Wk�M|k`A�����؈!�bs�U�f��WxU��E�¥P����D�)B<|g��r��s�n��(ܷj���IM ���sJ���+S�>K�sX=?��y���3�SaHv��b!���ih��6̈į0��w�,�=�W2/O�g�7���������~E�w�]Q�γ�қ�`��is(1/��p�6��	�ʤTL�B��EA#C�>�� ���w��wj�8�!��Q�DcF˅��h�#W�N:�l����Z����YN����E�vm@L�TNdn�DP��-^ze���͟\ܦB���hH�mQU=Z��/ �)7ѿ��#ʯ�Hʬ�>���u��­f3c��Y���K2��i�N)�mli�q���{a.L�R�8����f���Z ܟ�-E��-��)6+�3�#�!�$C3"��{�l}�J°��͇K���mP��9W�ЛTbs>�1����S����#�Ru�^�a����ѣ@�T���g�yE4 {�����VRL�<�^�}�#��<:"���>�܏K�ǜ@�� � C��G�U�:���	6܍��3+�eFE�|_���YaդP]��㊪aÐY�Z([`|��$���G�x�Y�qN{���{K_��he�Ώc?i�3���� n2J��2-�Ȓ���5s��~ی�&w�_�JY),��X�w�%��>��%9)�:�(W�����e�3@\�X5�!	���Q�ٟ2�e� ���ne(>��	�#E��Dv:��w7
��T�[p�L�_XKjV_]���ص�S�_��}�M%e?*��J��+`���Vq[�k��Kc���w11��A��F�kmފ9���������Ӊk���l��
��y���R`�Yhn�5�J�F�.�p��w߷Uo�.��ϋ:�F���4�e9#$<e�3�b���~���e-���f�oT�ٓ�����6�?)w��w��C����|e?���䵰�#��-9��F��6��S����3�}x鯭�
:(�,ʌ�+��*(OB�9>5̭U}��Y���wD/��N�����{�\*lǰ<7�A�(���ӗ.#��K�;�[�&���l��C���Ed�cҀ�{���GF�jG���%����q5��p�qE�vᰃ�����&8��V�ߚ��M	�Z�	��~��0�L�.����RM�}����v�K��iQ40��s9m��;OJ� ]b�� �Z��Y(�Fn��W�2T-jp�)=K�	o�y�-`:�-�J������������?u`���#��L�\r�_�3���C��+6�U�:t[v���1�%��wFO��S��̷�G�6�tʗ�*I�0IN�~=�� ����u�	K�EY5�%<]��{��nS��?WhM!����7��cEa�?P>���Gu������a9�l��xմq��ⴁ��0K�'��"�ڐ^�4Ό��Ple�	��>g�6u(Fl�����f��<��ND-t�d��=�c�_�H�2ų/@��-�A��2"SG�d"Hb�dI|�B\��HF/4�b5�
􅮯���a_���6�6"'��/����a��䨻�.Փ9ퟱd����q�J֋`1C��mO�6�E�|I���B7�̋
�H.ٹ���(=&C(?�~z{�p���^�2,�D���+�/%E?kKk��FkIa�W٘u���T��c�Ͳ�~[=�
6�ҳv�0۳�jGdU