��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��#ls�թ ����2��Y	����+L3���7@�=)��H�Ʈ2B r�2i�&VB����f�%8p��6���)�X��!_�����	|�=%��B��<�p�:O��TL�;=���ܸ��o0�a runh`�xasy��rO���C�ݏ��#��opي�]�<g�����D.�C���Z��a��Dl�<X�"5���T����5�;1�})jE�\,YM%���EYR��)a��"�3a;�U��g~��|��/@PJ�^��#��o~�����_�1`L�����O��'�~���'Z���nm���i�T��(<�X*�Sb�*���G����S�nL	�����~���Ħ���� ���yb)���o	x�Q����p���g�3-R]L	����}�X����)��f�?'���U�K�R�,���:6Bހ��?�w+�	���iF|��p���%%���\��ʗRkZܴY�e����c���߾�n������d������I�$�&D�J������q���ޡI"lH* 
��3;���P���R�گ������0�w1�O���R��%���hɕj��K�pJ�����̀nJ�t{N$��Ĉ����Hp���*E�0cU,�5�D 7���Ҁn�mW�G2�K
ic��w!"'��y}65Y�T8�JxP�j��{0[)�X�:%�S�Y7xDH�8��̌S�0��&���Lb�3��� d'��g����A~㚭K�Z�X�b�(A�t�yV�@nly#N���W�M��(�Nt��]�]�ud��Ed�|�ٌF��[g=�w�dO�O4��L8�'�y3�\8�ǧ����/:�k��8*��g��E�8�Kf9�Det�6�ǭk�f�l,�^l;��f-l~���V���}|+i��?�/����ѹ�㦡��k?��.~��C�l�?��Tޕ&)��yZ�	�1��7h���Q�9'@�o�N�)�y��l?�6%�6��<��PLVE���ӄbI��]�A+U��7�>]
�MKo�H@%�k����.FNQ�*���G����d<s������]�%=����Gˬ��J0*x�ڗ �l.wÚ\�]*��)U5�0����N��^M},i<��
W��<0����V�;ꭲ�lv�q\0��\1�V�ʼ��U7��#�-omj�(�x��߾��F2�H���>��g����y-v��ߘ�O��q-�{�\1�N#�}Q���y
��K	�̉e���Xg�e�N�ȗX��E���%�óiM�U��Ѝ4
tJ�G�O��sF���l��2��Fn�h�	0�C��_�U:�*|�?�R�2�3LC�s��<�S�&oܮ��4��(����Fz�8<�`��|�i�Hsֹ17b��?Dx�P�����q-�Y��M%�g�E9�$�����8i�`�_in(4j���E><�.ʌ\�ɲN��+Э�p�Ǎb������!t/�P�I�7��uz�`DZQ�3�M�jٹ{'������u������݆y�a/���{]q�v܏��#�#��n6��?V��,�@�A.���\n�s����������^"��1օ���v�^e
�G%	��z(Iߜ�`���D%��c���}�.rɨ�a>?�aO�`Ĭ�aD?� �2�?�'⾿�0 ��b��6�aǫ1ȓ=�� %F�q�)|���V}2��׋CB;�s�N��"{���pR?�e	j�>��y�}�L��ȇ
iAv�v�yu9�FY�d	�!*��2�F|8�}j}�p������5~�~�5���V���$��2�?<�@Um�2]�'2X�f��4W'צ�ew)g��<��r0��@H��dy�b��G���L[�gU6a���;���l�. [��"%�x�zך�O4��)F|�� ���f�|���oL|p/�$�}1�n�/���d�����8�"�N-`5�"X�9���)+2	�a�(W�7y�WC�j��r�0���o�����cE����C�9�q��l Ǵªŧ��_-��Xr�z�X)r��������6��RN#�?���G��o��]�zǛ�鋓M.�w��f��wu7V��%Qn�|W�D��SE������}�u�MQ�^�0א��b�bϐ��k�8��^�w[2p�q�Ʀ���<	�H��N@0��?�t���!j&��#i%��N�A�iF��l��>� �.�8r�3�-4��)�z��0��jպ�~Vܼ�w�q���	?y������
�8�uo�\mݫmS�0�Dc�c/k��lQ����!��Vou����jļ�<�<�i�x�L���m`v��\l��ҧ@\@���0�A�1��ua)�͆�(D;��0�����~��"�Xc�7��b��H�cu�_�z@�e��Kxm!׫�JB\��Ռ��s���T�����ę@`���
ƜN"Q����*���X�Ls4NB,tz�q�_����������.��ot���B�h���>n�N���2.�J߭���x����\hvd5x��=l�_N�g_ktR��!á�� ���B��b�HT��Ws1m���Պh/����K/=SY�v���3!ёu��^'-�[XkFR��B�����e��>gʲ�ѯ���13�4�:�}�������n_���7+/�-C���d��ׯ(��v��;��FKtc	$���I��[b(�mF$)�Z]s;�s��jl��j 7F!}>&��&Z/b� ��S#������A�m��$�~��P��+}�+��Z�}b<�_L,��;Dr��I��[�������b�xLq@+z[2p���2[ޔŋ�j��3y|��Ѯ��J�&]?�no7Z�H� ���E��rB�]�'佃\��Ĉ1\�d}n�sB��l�f��N�t��$,sؓ�V,�=~$t�Ȃ[mH�a�ܾ�̣
�ݫ��(E�4=uT�&#~���+�cN����0���ח�Ni������rf�Dlam�:���&nm�SíS���8�C��d/�������+)Y��GV.�1�jfǃ]V�+bhd�vp�.����N�����=�5�� F��vt����~~_�ux���񼇯ޕ�8�n,# 78.+�!����2�� n�]���=���C�#��_���Uy{��|���wc����}�c�eIβy�H��b���� �6"H��U���W���A-��rϵ7�y�$|�p>��b�*���Q��(p~����A��rT�@?G	H�t�kY�7��~p���Be���ح�bҴ�Y���*��3����#��{|���K<rp���CjLu���׫���X]��5)=��_tbo����IXU���`�w'���RG`�2��n�ɩ�t@�R�ш(�,hP⢒?'d�U���6�{�^��|�u���c1�i�v=<�s� k��B�Y���ǿ��=F���y�c]��ƙτ6��4/s���SQQ�\��JőP���`V��3���e��1�x����U)�6k����2E�R��&%�
~ѵ�lLN�[�$?����j�[��X�����U���<޽��F(�<Y����yFl=.�-p�&.�G�C:���:u!Ǥ '���W��:k��X�������u��\�2��妁��T寨^s���'r�g�5��"����l}�k��X�h��s�RW�����#��%�����6��9���ZJx5���`�W]\ϯ�3xF�o<N=O�����K.]s?{o4V�֋����x�Bz�2푱)S����~���h��f/�_}G��������i�y���6��+��kud���7�|��`P9{�=�G��9�m�D��~&���JSA.j,���z�c1i��v���*�����h����%F*!��<�U��Nw���5rj5D��j�'�K
(hF�%��F�VS�\5�$Z�a�����"�qq��G�
��x�R�ͽ��:V�+�NS"�?�c/x�~��Ў�rŗ�_ ��@���Au-]<�HJ�ʺu�kŜ ��R�z+ϣ;�NqN�`��3����kf��[M!t-)z��M�m��T�O�3U�E5'd`�Pl���5��� v������(�T������:����|�Q��%>Zr@\��lQS� 
7�\�[�U�}}��ex��2t
�~3��Qm1������*����^� 	�˜��f�Xb�:�z:f�L�P4���E��s�7�&�A\=<�F{�c����f�(����:B���6a��?��`�j�`{��J�S$~���Af�k&B��6la@W�gx%�TZ�1���|�>0qd�S���ڵ1�;�0auG�wHj�Hn�>��J������7b]��Um,n٧���B�Q��`!~9Z6ቌ�" а@�I��|~pME�n�W�?M��c�w����|K*T�Q@�1Q�2�O��(�쭬,���[\��EoY�i,�U�q]��ҵ>�J���(���3��e7��y�E�X����y�7A֕gü�[�-�l�C�Qz|��]��z���3��7 _U���BR@XjjF��=YQp��8��"������W�\ϖ��UD��m�X�i/�[k�ӻfWc���@ x�Ӭj�9X��6*�kC˔S5�6�o/ο�g
¨�M:�uù�h���\M��R��%]z�g�+2�r|�x[���}��q�v7��Q��lM���@�2ͺ�@QmѾ˳�[Ĺ.��0!����&�
kf� u�WrNi*��x"/���`�"�s���=[�V��å��y� �kF�F}��2�bօϹR�5j��4���L��S��WN��]���`{C�Zn�����V��ɏx|�6RN�a?�{��-�2E&���	���44����Sbhiܙ25�c���
�|�V���2���h�l?���z*ysy��A��w����e��2��I;M�����1��/�T��}qڹ�Dߤ$e'⡂�If�M���4�3��7�A�����~MYqBǗ�@E�SYa�0�Tf�b�*��T�m���3��c�l�/W��xߥ��7N�Y/A����W�����5n��洛䔒�ȩ.(�=L�`j����@j���k �ce|�xց�O��PR���W�����~Þ�m!����M/��~,{���{6z  vp����r��H�5b0s�c�k��k�4��B:r�����fOb�4���*�I���(T�QM��k�[T�|:�,8p'�S28%��^�[��2�^��N�F���H�2���?�����˳����,L&���j�_�5Y&�sJH1º��ƛ+FO��/�Ur� �F$�
�,2Z��sHO����_w��z�Y�{�����iAȭ:�-�^���2;�Q�e�b>���R�*���ǜ�K4����҄�#�~�_�;ڥ�Lfo*jF�� ������`�aw�+$V���k���B�u$�зu�����'M��V��X�������n����g+�M�tNt(�3�d�}��K��Q?��y�c�Lj�&���X�,;�o�K�nCG����2��N��zM}Ilq��(��Z����y��;��u��c�Z%�ct��6z� �
������&���y��^�����TiD�	/�|��}y�f*�\_���Vo�a5�n_�+*X��Zc9�\�4��T��wjv��YY��h���2�ʨ� 
m�x�FU$�����B�֬�)��7��$q�b�M�U"��;�3��a�҅�?`�����/��ER��;��J�����%�u��Ǭ�� e@�����G���S	�*��5�\�ݓ����f� �AP(ϯ���_k��)p���=����Lئ�)�����[����|�9�Yl�,�������S���kD�����L	Z�~-2���m����7_�۟ӳλf���;(�-yD��3u[>�*����ztg~^-z��$�� !}��weL����ʆr$,����G�&���z�}�F����a�z�`�v�~-�]��H��z����8�z�8�G<�S^����J�Ͼ�RӼ?�䗝�����ދ���,b�/��+�߇i��՟0:�X<zz��{���O)���œQbV�c�ڱKb�3/{n0�K��A��j���[��ј�QF)��D�?/�dc�_�8�f�vPB��
�Ч^K��	�p���s����u^G���8|���'���؟�q���1b�@��5�dpw(Y+0���G��z/��l���oxӋ�<��箃u8�9eخ����Y� 6���>��c�m���f�)P��_R|�ªk渴k B��P��2m�������k�P��<'�g�@�V4/��Do�7k�p���u���p��r;og��v�Y���k���Xea6��=�����K��mWʹ�ݨ�A��� ZF;)���Ǒ9�t|��.����%u��Mtϡ6��V�5����W��0:�f����b-	�O$�>?&���ʺ3���Ly��6���k�$�&7�ԩ��q���EBT��w��/奤���U���ο�?�2ã���k]�Zi�!�"��/���(�U'�����\H�+O�ѰApyl$�xe6���j�PkC^&� �HK4�S�i�$���!߂�w��F$�EmAV'�c?y�8�U=������3/����LVx`�A\]�J'�f��u{
�ԡ崇J���� �V�B7��d�Y��p:�am#���������հ,T,0��l������/|�R~�W�<�������m:&�2cp���BȒ������+Xs�i�� 1��;�?VaMVN0+��@�ˇ۴!<��'ʤ��w�6x������C��JF�}KB)?�;$T�^*^����Ñ����c��53��5�c�Z�ܔ3��K���$��y=}�N�ro�W� �.��V��ͭ �
YsJ �ܞ�	�E�]7Rw�/��-b���cT�r*��Y��ޓ�����H�E�No�ˢ�t2�
�kwp���w�DE�N_X�O.�I�K���?�� ��By�ct);k��\d�;ޔ�lWǯ���Yž�_�G.C�BpY^MV�.{�wl�jrs�	�Q�D�)�o1�YP!�����+X���3�O��ₔ#:Î��ય�V鷙xK|���"b|	j;���D�6ݸbطX�R�C���y���D������"�,�['
LD:iU�=s���׆��懺�"+0�S%L��j�����]h6��3/Ik�����Ze#S���='��q/i��s�'�����.���.�v�R�qx��}�\\��0�ـs�����BySG˖����v�L����Kb=���_3«���b�\�\�f���Lg�o�Z�j�Gi�Д�a�G�U���&�p$*#,!}��u)z��w%{P	T�A�K�[�i+9S"0Sc³�ǎ�/�K������4	��#AU��Tu�x������w-���^���}CՀ=
9L���� m +�I��l;�q��{Zc��	)PT{J��#�������{ɑ�sI� ;�Ӭ]'y��D`�"�Y���u��c��?°a�2glntk.d�;�����gs�;��<nx�Z���ʷluF}�QWg'tf��C�%Q�����;�֙e ��J0xY�c���Ъ�z��%33)� L���6�a%�����O�/B9���{Y�%{H�����NV��e$~f�my��z�k�nuc����Gt�� a����x�y|���%�f�4�)ϰXt�\����K �M�����ܮ����X�s���Af���32��?�W��ױ*O�L�dS�m�sl2(k�������Hj�陌1�7T�����E�Kƨ�d`t(g�z��ǚ|���F��,q�eqW-�+��uT�n꾕ڠʹ#F�^��扎�3��6/&W~ �ђdƲ��	;��{F<OQ����1��(��3�*�ͧW�~ڜ9ub%��������##rM֯��r���r�I9��jڱ��Ge["�وi9t��}����@��E1��n����:oT�M�YO�2�^H\�{�r��z)��q]}v��o���ܾ�TWM}�o٥z7g�W�6�]���qSwu��a����PTu���T\R�5����|�J�t�<[w-°k+��ʇ��!h|tKk�F�e���������,��[[��I_��c�>c���3��mb7��W�5P�E� ����AE�l�a��H!�"0(�	荍��~6{���@�������25�+jσ9�6_�u��a ��ĭ����k�UF�'H���r	3��&\��ؔ����ͭ�����!b�/�Vf��n��Y~Nbm�����ozd*Ey�e��O&`�9g�q����.ޘ����xH��ǽS��AZ�����졡C0Wa/�<�z�gL��.	���,05����y�VR�y�zؿi+��m�+���6�aZ+���.[�@)��*7����P�.�U/ �,��Me��nB����{=�"� K+�6<���x�-U�D��fq]�
࿝�x�"S�ڑ: <:�M��z����`��ș��{�+���C~���y�U$�_!W[3o6�� P^�Հ��߮�`������Z��ڢ���<��9U<��
c�䅭:2'��23E�	�3zUj	�f_:�'�+N
3S�
��_��h��p�fՅ�`�noh`(��M��FE=9�b݅�mY�S�I�ŻJF�<)z���'�[cߐ`����͎��'b~Rȕ����t�A����E�G�Æ9�E��ڵr��[�T�qSD�Zg�yQ]�#�yB�M�a�_�h���(�����*nx�s��vB�[j���<�7pFm�DXs�$�e���ǰ���"A��D�	�E�!�����f������
�[�l� �m}�R���M�J�$sB��!ZB|֎=��8�ʋ��/�ߩ���ED�H�Q��cݝְ+�s�v�g.jS�6"2��89�6�Q��#��e�,��v�>l���=�E0�.��A�� gp}Õ[\O-�w�ҡ<�r�X�1�Gˤb%��/�u�9�<4�J�=��#�ey��v�"L&0�?v/đ��6Ɠ�?��[����+�_ê�3H""��[bך6`y�#;̞���w��Q�}����'7&�{�sH��Z��:�0W����v��g �9���m��c��|T���O�(;��XM�M�����y?��P���}�1t5n�F��\h�����4�s��c4�k�Se�� ��y��J�C�<��KZA�+���
�nC26Z��Jk��޽�(�Q �/��Е�"���χ@�1"�ꖐ������&j�%�}[h�hJ�l��lV�'3;�ax�S1��/�� �)�Z�?��������_)P~���ﬞ�y�u��Mr2���A;����J��A�'/ݟ�!�E�8��%�U-��י�$e���ȡ2�/e	�F��P�� �q�|ػ�»����
�4g�\�4��{`G����	ԟ?IK� M�$�(��s���|&�$�s�N��S�#u+���d��T#f鼹d�A�-U�Ur��p��ً���9]�f=3	H:�3Gv�	��Bq�	qcq�f�s+
E[;t��ޝ������%��8Mr�q���g�0H��΋O��Q��a����.Y�{��s�6�h.쯻���0*�m �r5`s�~�E�������;�&��:���$,������p�0���T�ʵ=��ݤ��8�[�j��Ϧh�����Y}�X!�m��::98T��+��_���X�ŽְE�B8�=��H���?�Hۣ������9�}Ƌ��m�l��$�Zp��׏I!^t��"�2�7a���y(���O�G�WX����VB��%��]7$a�(.u����[�����a�nEv6�j��:=�Ny Ů��7w��=F�{�k�lN� J�#d���=$8�!k��;e��9v~��p��� i:�Ϻ϶>�ϊٯ�sh;�ɫ�A�~d�4���4a����Ղ��c��.�{�ς�Z�Q��Z�7f��SץW��5{���%����׶ `&��q�wL��վZ�(�-i��IhS�b*�y|� �L��nŎ�\zZ���G��`g<5,X�����.G�I��O�;(�3&�:�������t�,+��G�O�����T�p��<!��HY��	�6©���*+Y�͔ʽ�������6��P�֘m�L#���dc����5� T�#_E R��)���3D�W�wk�ɞ����:���T+M���6�� >t$����zPj8���ρ��>
�	�zK>J���w/����j]�e�>N7E���+װ��R��{���c{9ɇ>�R Y����2L�TLqІ�ÂI|Ȇ)�iA���\4<�����¶=tn�?��W�K�4���H�����*��\�ӱ��zA v��*&f~=��SV/��`�:��	5}� �g�5^�f��hIj��0dU�e��٫_ D~��9��+�L���ABǋљ/5�~�q?fc/�����_���*:��t��^�s)��%�zǶ����	31���#ڢ�x�7̨���qH@��=dD�"�D|�������5��̸1�)x|R'x�[�6�t<��?{bƁ�`��"@�	���R��bn�N�%���,�NK��Jc%j:���L"ڇ�0
�����m �s'	�,|�Y�j���y�� ������,�yss�4Tn��T�� -��Z3�� #����>�a�]��P����g��F���g��'�����E�橁uC0�l|���M`�]�F��.��D5j:���vr�ɢÖ�ߨ�%��2����6t�#o:��Nh��$�W�5^Ι2�=�������H�
���X�����Յn�T�h{f�	�˴�_�*�NJr��%�E�7<���[
ȉwv�J�8H������{f�%���܇f���x2ĕ�� �1�l�À�F�-�W;�V�B�����	f�K=���t��Q�mE'��%��M�^�FhӋ�ͷ�y��	�h+�c���|Qe]#ح9ڣ.�,GY=��T$	z���tDr�ݎ�v�U>G�bӢ��7'0"���|_�+�8FI� / i�T֡��1x��]8�E����7���gh��H��]j+2)��_Iω�9Y�%��,�dk�nѕ�\�(��)5;8� }9X���VO����?�j�j�����?.\�p����)����E~����rg�v�H�N����P��>�5+���5n�:�+���k5�GlJ��tt����a(��|���uj�����^D/�Ω�D�o�k��M%X5�L����P�`:�ԍah�%"�d�@���ޓ޵���t�� �
=�"�xS�������N8����K�T��T�= �s��*�`Ll�_h������K���Q0f!�j-�m�ŗ���{�U�����K�K���p0����W� rB}UT=��#&���l�"2R"�X��eH�b�	#ݜ�|I
�D,X3A͝�}���O�.!w�9�P7��}����%K-<$}����7�"���_��<����v����iYg�;�6���?@��Y���3�ו.�׿{��M{s�4�[b'����I�Ʀ�-G�>{�vx��?L&�P�&1C���񭚸�h1����GmQ�A>�b/�Q��L,�Ë-_$���4ҭ��7C\����K�4�C���C��H��ˊJb�o�*�r&_/�s5|�e�p��>�.d�(�%�b)rh����<d��Z88h+M1;�gE����U%A=(����7��G�*��L���Q��
�̾:��1�iJ(���$���:0#�Oa��>�g���=؏��x����V�s9%
��]u��RL�`����E�Gw]zce�L�@�U� f"�i̓�xJ�~��Sw�'&��}Sm��Z1P'&m�Dr�5A����q����" A���
�hֶ�Y^0�e��]�&܊3��hV�.N��k��PVU�k��'8��b`Hu��R_N�e,O��̠�J��t���Z3� �c�� �<��bax�Ȣk*>L2yI3��`��I��xiC��eʘ'g�uV���]e���pL�c�[#�P��d��*課ݛK�Q���ysb�|Hf7[�S���Y��v܏�C���#V����I`���6R�-&j[�#H��v�7��ރ�i�	�G��z�c�{[�v}a�NQ��G��)�w��鋚�>�G`��D�H%@`[��P�T����]�X
�R��+z��T�QĴ���P�0>�A`7��=m��\�+��j�$��"a������b=�E#���<�)�a�El�U����{����:RZ_��r�֢�����v���̬�8G�2��1��t$uZU����KhH?����<�'�gN1�a!��89��?�~�A��GB3aÚ��Q~���5Ѳ�O2K��X�,�O�|��ҵF=2l��j��P9pj8�1�;�XT��֥��{��k����C�0��Um��]k�c�Ԧ5ب�E�!��u���cمl�3�	�,�U��ȃy��oű6����s����>���EG����P��sתC�D�_�<�[�p'�T����������r��gn^ÙM_�n��$���삗28Ι���wk���\��H�2��J+"O��� 'Z����|�KI�	��<�&�o��)i7�7c'�g�ݻ�i����7@Ya��-F�O�x�'�e�?�+���G���?�%���[l#�UH`٘|V�5�.���a���B �~~���7Q�����)�phl Eٝ�����?�B��ZI��0��cT�����%{�%R�BOH�.*���|��juǽKga����|���bK}~����&?��N�[I��O�V��x\�4�=af<��v��?�Wz�܇����(�� ���� H��K����w��ސS6�E�u���p8�.���.S��S� .���
?X���D�k9}���@�?-�k���K�n�Fl%���9��[��*/K�ȸ����U��}'�4�e+�gV�|��=�A�U�S��B��wv�fY~F����r�ɜd��	�0��2�B�19_�+|��Ah���s~o�`k\2��Z6H��|�P��}p�����Uߊ���u4Ў��ۈ�>wԽ�� �Mw��{{ؕ�93o<z9��<�	��Q���G�G�2-�e\2���������Ў���$�8@�z��\|` �8�ut�?���t��.�EY	�����,��)����=��r�G��P��չ}�=s���H��"�}d����y��ΟCiE#�o�C8
nW��.g�{��$ad���;��jH1<r�퐿#S0ڝ�\�>+3�
��`�l1>�n���;B&K�J�6$̛�<K�T��P�M;2���rl����@��,��Ӎ�O��.���쟊eyY����I����^���L��^�D�O9V��s���Y�N�9U`���9��r�aA�r�$n*}�߼Z�\޼En~���%��'�2dj�*H�f��_M�B��?VP����1����T��d�!hk]�ZY$6���6:�} �5N��������n	���qK��m-�q%
����� b�&��RRۿ�3N��4+�.�9���HBSV�I�Q)(��.�H��$j�?f�U�gwT��d� G�ݵ�(�=L����D��.�ҕ�R�񶳶&�k�X����d �6�3E��Uo&�/�ۚR��嶀v�2K6r��m5X%8�V �i>�}�t�C��_a�Y,�J�L��e��,
��/�E�ZL�?�u�WňU�	�� *м둪ɦV�����#��~��!����S�}m�����憠W����bW�*_k���岼�URN*R����%�����w)�)����$3$u��綜����:��e�ҶFaX!'��-?��:���2.��xT'��`k�,ޅ*3{"j4i'��̿b�ky��~�_��vN{�TK�Ϣ����t��U���.!#�$i�����g��[<md;p��û�6[�4D�䂢���#r�YMݞ/�=��a-��9=�+�o�Zh4��c��Z��*vxJRZ挼�&�˟���>g����B��l �@�HV�FQtIv���qH�d���m&��9oO2�|�$:˽�7[��r;���n�������E=J��q� ��P?�e�_����b�m�jƦrl�C�$~O����grT�}�5����c�g����̲1X��?�=���h���#q`�כ0�L<�?�,�z$b��)�������6�t������-a�z�%t��������:>���X(���|7{���+�5��,Ȍ��[���6��{w�~J2\�������4$g��Q,�C���IG�� �����nݚ;X�z�	�cU=�@f�  B����D�@�nO�Ol.Wr�[ʴ?���7�~���mCv,��Ր*X�B}]���n֡/��g��xy4��r�;���"�O�����zq&��Nb�נ���O���B*���D���H�3w�0[B� a����R0:�(<����#���%q�l�D�$F?��
��Ƙ&CP�B~��l�f�o��Vפ~[nF�s���V�� Q�ߤ�J�����W���|�ݕn/Bce1��1�JI�љq�Ի�W�'�~�r����r<G���?�+�b��>��E�C�lr$��� DN�Ď��b�ȃ�ՙ���C,�8�tcJ��Q����|b������T���x^��2~���k��()��#+г���@]1���3��f��� �������^�*�䗚C�T��x|���Ն�>��s�7��;��2��
�~�u	���~Yy����7���6�������P�>�~@�?SY*0�����A"��X�h��v���=c��_��r��Y�겈�d�wp���گXb��@Y�ӏ��n��$Hm�'�������%��Y0ϟPs���%ŀ(GB5l���R��J���[�(����1.���􉎖�%��0��Q�e��C���
s���V�z��Z�u�WR',!)a)@�
�X|���=�X�t�5+�RcyX}v@oj)�)
��'r���N���h~nė�e_?��т�1
���7	��@k��&N�P̹.B�Ʈ�O��j:k[k$w~#l�<�S�Sq�z���s}���m6��IVح�/�`�#'ܠާ�"*s8�q1>zְT1D�_���Ԁ�=�������W1@.��9jg*�>V �<�A�6��O޿�����̓?���}3��h�Y�ܳ��-�WF��5RS?t�R�
�=K�,�3#[I�Z�:�xbu3�u#|���V� �᜾�7(ɍ���������������Q�)|�U��[�BٓE2)KFaln��M����O�}�#�>pX���Tb����P�
�X��U}ϲ^��
��~�^}�%v��&�#��]�����d��ҥ<�n#�S��ఴ��l�N����?E)Ljy������W^���\� ���゙�˔x�h��ǳ�t
����&�?@�@���d�����j�Y��ʆb�$[/S��BJ��NE���<26����U��rb��h�=fl�ђ��p��#����]bg��u�+�2��J�,�,��ǽ�O��{6�@�q�5CV�i�+�_��i�b�I*�;f\(ʌ�/ؔ�7�uG�n���𔕥�8�')
�D:�8N���J���vJ*�U�X��
-�7��� �k9�!RV�lx�������t���;�f��tZ,(��+����v�RG����"�):�22�%�GănG��h� � ���{�|�n�e�����3�k=�UC"l�ClPl��--���!,��s�Z�S�;����o��]�Kxԇ�'����҆/)�s3���|VM�0��)��"�=�B�P�Un�G�^"'9����wwgI�t׈phU��&QS{T��{�tCS�9��Ox�U����� ���_-��jT���N�r��Č�I�JO���[,�Я:-A�pHq�����7[��1�jC�>�nl
���O?�'Oо\C�n�:o�>��ҍRf{�`��m'VH������P�B)f����oN��s�r�����tGfQ��K����4c0����_�xI��`4s����L/>��S�&�A�r�pA�+^	�Q�6�C�ߎ�a�J�H��dޛ��yӽ��	�O^�B�96�;���WF��;�}?�����>J�$�"�؛��!�u��īM�fr��a��^�Uy#}z�X]�lW¸t���U����ϲé���XSc�8F R��O�C"�Ə�^�^�h�K�bW����2S�s}�FT�.4�4���eSc־\�����q�j�4���dqo�0C�O�)X	��5��Q��$4K�
u?��i�����﾿tߢ�$U�	U�a�x<W�'�a.����s*;R�@�3L�A�uD�̧$��B�r�(h8�h߸�?�������؀����a�w휎��.���d��_��qp�G�=����>kg�y]�?»���̠�b��/y9F�B��WG��Z��Zd�P���l �+w[ۑ�o���""5B.$���5��KXu�C×|�t�+�Q~b��W�ݥ�w!t�l���I�&�R���z�>�8��P���D�L����k�Gi��<9�m�������$�%U|z��ꒀ.4��y�X�P�O(�s��KV��s��-t�[��j[�K�O�_�MO⩙r�͒�b���첈��ǝk|�Q�hP[�s�bg�E���>1s�F�
>\R"%i#{�!�Y�P�w�b����Ft�NRٲGs�8^�@�֗�$F�KR�ǖO��"�n�z��	X̙]�j)���^����� vM��*Oo����xu&H���"��4�e�'&����t�zorz�z��{p�ٜb�?mD��������Rl� ʵ38��o�5�b��������#�Tn��4��nOy�1�i=�󎶜����d&��ma�Q�sS��4�T	$��3Lq�!��E��B\݇� +�R}���)!����*8�	P��X*>b�Y�4����g}��-b��I~{�QE�"e=�ˣ��A�
���8�<E�W��6�s��գJw[�{�� �����%����ؗ�i�տ
b��\/;��?_wN�NR�����s�
Ѐ�N��dfI���]�TWnIV�Ҋ����R��I��d,��EҸL
=d��D����F/ �W�<6���P/#�n�և��$�G�.&�r�o�J�_��L��l����$1أ'���R,ʼ��k����� ��Մ��1�{O�����L"|�C�3'���A*�>��n��O�G�T88M3��W��*A�Y�9�%�FmO���V��d�<Ih�F� Tq���D��tc�1p�d�Pĥ��V�����B"}�n��*c𰉻#a��19ŭ^��ԷNJ~�u����y.��x$�ơ)�t����!$� �o�s��ȧ���Wo/���L�ș~�$(�KM��h��Y{������_e$Y��緕��郉z�z>��c.$��r�W(����n�1^j�4��(�vg&�T�(��E�h7=eX=wbp��C�@붊��ӆ=�n\%��&�l\D�C��h1�冂���ko��OT��a�6�]���l*9�z�E�@���r�!��0�喸�M�@0�/ ]��B�C��-�c�Ձ�)���.�4ѴNӫ)��6��O��.x�s1����~ ��$Hը�O�<ש#
������5"Y��L��7�P��'�6��\3Ӕa���Д��,�`�U�l��ݜk����(rM5���$��Ndf��]B�۳'+)��x�B`?H�'��pN�ڝ�Vc�=xa�@<y���ڿ8�jD/���чtͺ�[�Hجs(�X�M�.�#�	�h��]k�J�sϸIŐF�6�ׁ�9�雖����5��×�����	�����ͣdLu-�%��5D��3���y�8���!����1'��a+
���Ny�o�� �wDf (�O�E��8Bq�e-Y���$�
��QR�ru��a�����~8�5u�pokMc������c��!a�E�m��3~\d�KD �t#�V���Et�IpZ���^�[�������Tn�J!}�FJ��z�e.l�HP�ί�(��}�	�j�n��OYfoeg+�i��A����b\�	vx8EJ���_��{3F=;�$f�w�(��8O���Q����v��M�A��
F�ʹe�B�ED� ��@ f��>��gMM���t���4ٚ��?��z�m��m�	�(����>�D]����p���F��?�^��@��8
�Z��̈�p���	6Ç9�O�B�N�.�Q_��VG��ن(��3V�����+�Ӟ�����z��"�d�r:۰�1���?�<�t,
�SCgp�U�z_� �}�GD&�"]�! ^�U��D�?	0(`���pfja_z��f�Ԍ�Tṑk�rb4��[j�i�{8�gE��>�B�Y�U"N�y����AY��~~�1�I���О(�kZF��sc������9�T(���7}����0K7��W���W7B�K�"�b�`̄}������WMELƥe����ԑ�ž�~��*�����(8S�b큮����$~�Hq 0l������U�uyȯ��#�@�]t��D6���Y�	��<�������Y�:rp�(����� �Y?.l�?�,p���Խ����L]0!W^*9t�L�a�����y*_���sB�x�RM�1�WH0�?�\��(3����Y��5fn>�H,.�3M��۽��ɱ��Qu�W<�hI����D;��l5��{}10����5'ٕ"���b2�Mw3m.TT;�7�^�찻4�M��b�}���o�t�6��mրU�fw*x5R[��(�"�xm��.œ���%��ٸ���*����Ֆ�yһd�"WVi��նx�q�-`m9�x��fu��۴>��?�T;�̸���[�/��%���|E�$K�G1�Tij��}�����t�N[MewrnU��@��X��5�<kU�QPuז ͚��>SA.������l��>4�`��Kz,q���-�'q&�)�S�y��=�Ք��4��^ 1�F�����[��9��҉�6	y�r��22Z�'�67��D����I���k7?j�aD��&�8� �I��[��{��M�xw��ͷ�#�C]Ƙ�K����VV8�~kms���ަ~���rUA"hT����,�*��R}7�����?%�/�R�rV�i8'��ؙU`h��ּ�[�铕8��W0?M��Ta7o��S�]��{("�֩r`�G)�Pf-��.*��t�#L��%����{�c!p��OO���a��w���[���V2%R������ƢB*�O�Y���(t�-�/����E�1ɤ�eҖ�k2��W֥e�+�C(�h�@͔N��v�[�9��ej��-���ly��j_$�D�[l�Yf,[�+�U�X��E�?j?���¯�Xc�y�q�wȰLʰ�� �����3�DSu'}!n��Ŗ!8�BY��N����U0����ӑ�z���m���53��h�30#tcoF%L�� ��N�TGT����@��=ȫ���$l�Wn��,��o����Qą�)�]���C��Wzb��JQ��&�luy7��_�<V>��Y�8���cD���݊4�)f���Z�|�1�Gy�v-t+����BwA鑂d"kEA�,����vQ\��������ݾ�S��,�y�Jhи?�t�?���u��	#L�$%���`"�li0G�b�'�*�E4B��Ҕ؁89�U��z� �a�6T�5��(��Z�;��bb�6��X�����+���;�5�8��ԥ�]�ѐ�Rn�/1�WZ�e_�E�m���)�$�!X��<��ޡ�����?/3�����v��?T�^�-��z[x������d4N���rq�u�h܄���Y�,�8��[z� ����s���kR�N��Ű�}֢vK^�,\?��R�@��e�/dO���'�@���q����n��G�Ս �ē�?���E��l�u/�>+�Ձ���^ij��Y�5^2�v	)�(aV���U�( ���i�c'Kj�w�&�k�K��%�=8� |&� �oD�W��U
q ��A9��wCͣ�/��i�m��Z2��4�l�Ǘ���̖��c;�+���zl�*j��u�'�N� ���O\s���ȗ����HD8�� �D.+u�_�6w��k�����B_������z .�A!,)�?3I���9a.AW[-wFh'
�=�Qe�-cq�]C�)��8ހ�c�Ֆx�����%�� �O9�����{�Ǡ�˝��ǐ���*s۝-)�A����n�_ub��[�sN
m�� ���I��(�\k��f�@z�(ǥ�����I��=�Dķ���
<�RL�㟿w�$��:/l�45��`E>��"���`���<�:)oU�oH�Pz�Zp������4�IC!�Gȗ���Q<ۑ��]\k��+�)6'Ɠb)�bcG��`�v��B&������S}�j�&3��<�B L�la���ѵN{҃��3喋�x��]-�ayN���ד?�
������22�j7�h�Vt5���q��E��Ic�6S#��+���f��|>������B>N���7^���t���&�_[!Sf���d����˜�_��z1�f�ȑW��m $�
���F?;�q��逧6 H��tZ`��R�rF1oT�OÃx$�
�Ƿ�Bp�ׄ�����'�|@��č�*�!h�j�#�ὦ1�����N^[���{;��fM�����Dr�~ :��))w�!�pKH�@D�8���}S@� �u)Q��`�@A��Lt����X.����+�ۉ�L�ݐt���e�<�Y[����6�Q�ǔ�K�¦����F�6~|Q�ߍ@���uÃ�B#��L.���]n�S��v������dp�7�����H@oB�J(I�U�ػ8a15n����	B^jX��'��Mo�@ �}}�����.$H6i�4�,n7@�0_h�N����c�b�!�C�@����F�z�^|�-i����k���AUIZ�vӈ�IJ�c>���+Gu�lĢѥ�'2^to��Kpo��w(�����\�DM�V˜%l������̊5I�����
ȅ�bс�!��5���A�E�U��^�	ca�q�a��5B���	m%vBE�3�;K:��Ro����Rhat
����~Xk�y�d���L	]ޖ��äԊ��kxZ�Ն64�E�+&��*=�H�E.�r3+. �#��{�rB��\����P��n�p&.E>J���Ч�8��c�'����Inp0f���d�����6�ⴊ��� L���Eo�y�Z-�'3�V��\g9�B���z���KF�!3���	Q)3fa2�Ϛ�IW YG��]��P$�aDN4ro����Ԫ�ڨ��Iɲ�Ѱ�M��;���Y�0]�դX�{JK������j7��V���J��6?U��Cq��91�
�؃6l6^��g���/ߪ3��F�(hX�7�
���4�f��c%;��x1��uK�y�Լqr��wލ0#�o��i�(��j<祕��4�+*��Mh�;���3�OѧB>��H���e.�r�#{,:�9�9��7�DΩ����ה�x�K��X�3̽꫟�{՟S�\+T�R�z3��k���@*��ǃ��(�`��2�]���UiTg���*dL�h�k��l���m��AVdS\G��1�D��	{9D4���U����5�Qՙ.���!�N��n�?^�����Dl�>qNG�co���J]s$��pW���N� \W\Bf�@L3u��*��Ȟҭ�e\�M}�;�W���v9�g��?��V�;�ŵݞ��4�H��p4'�#���������D�^�ܧEY�w}W5f� �I�dC�c~�R<�UM��Y ��")b���yC����+��V��@���_�P�Li*]GRѓ��͟��aN�O�%�r��\�t�6G���
j�����6�m�y>���-�ó��f~�8����1�u髫L��<�w�tfz��F�1h��-˟ܒ���-�;0������ �#�հ|9l��M�Y� qs�묦�K�>�/���TL (Y��ފ�E��'�ġF`�o��R#h�w��A�Ϭ�r�{y����N�_Ɲ��1����B�����hNT�C;��Т���e�H�R��\�?�$�qk�YƉY��@+7߲-{�ܕі@�_3�r��MϽ���3[��0Pj
��j�މ=HP��B'Z �l��qY�߉�F���+�����C5�7��uN�fE5��7�L�ؗ�;b���՝,�����YT���u�;�VFG�Rs�nMyu^�Yv��,t�4�<�$�=O���1��bk�pr�����h�������A��#��i!��,�� *�haJNW������Ȣ�l��
��t�����2x���x#�^���&dm�4 �0�q1e�����M�lϨ���(˒5�#�^Y�S���	G25���Œ͈��a��F|DT�C-N�I�#q���M
�[LguW\I':����f��0�(ⶸ�ȿ-^�PĒ��{v*���t���cX�x�ilݱp���R��b�k)OY��ܮdR����� ;��xˏ��u������)����c<Ҟ@A4�۬����:w��f�$�:䭴�e1�GD�(6�!W�����><M���v�͙�H9%����6�Gx*E�	{��E�M��7����H)�f7ʬ
�vV*٣�b�^< �ٖ�K�C�	G[��&�3a��덇�,jZ/�:"d��u�bQ�TA���5~��kD�D۴k�#@{�M�~4����ze62H��#�xx����u%WY���3��R����3ؠ<�˼h�����-q�4�֜A���sC�1����(�Oa�����}v��zk#N�J��(����XD�L�4,^��}k'�Zȱ$bQlݖ��@8?���Z����X��7qsY\� eWv7� ���e����n�@�(=����2{�$`�t��5´ $p��WLH��a{����iuu/��$$ \#C��������Gp|��3��Yrq2��Ac m� �A!�ȏ!�	�U�5�@�Y�v�Yg>̴��LaD]��Q��g���^G�պ���#�:��-�+����X�X��=�+�O~��cL7��g����8y�ܫj]��O��X�B��wZ]���/��I��YʗQ=0�p�>�H���?�T�$t7*�`MZ�fi']��N�B��g�j��&zǝ��,x��lJf�MK�O#y�r]��rp|���M�֗0�U��F��LL'�­EΏ��Hz�������w�*/�=��gĮ�B&����0�{�؃�Z��!�L>��o��Tn���<��V��U��.�D�^�h>\�@t����^ЁX�ZV�3�?�"��@���K7�R�I�����F�l��%,�����O��y2|�)���-R>,�ٷ����w5e?�>��ɗoޥcx)���'�o��{�V�P�$s��� k�����_���Q������|���{H��� ��m/�fm���]�Ac�4�k���̱�b�]y���QY��aK��������b	�<����f�a�"�Na����@s{� ":��i�]�Z�ziVީ+Q߃������V3b���0����1(�<
������jA�mq���������܅g����$�#m.<��hp�?u^a���r?o�*��#U���a%�o�ӛY��̸m��l$aC���"Yg�V]�ji�?2��3��Ł��ǒa�N�-W�26�#��p��25�H^�`���^��b�D&wx� 8���4"�1�⠂"����ĩp/Ћ�7��&z�F�� N %�i��e�����,#X���{�����)��`<�t�ww���?�̊���V3(;�r��9����7NaJ a�q#N�تG}V�c�q��o;W��
���p�`�
ķ�#G��%.)_���
'x?@�o��>Jo��ٻ}�6��S��)��"-@/	�}R��D	lM2 , �h�G�[��~�ѥ��y�����$��t#󽻜� �l��F�UD���?�F�id؞��Po�?5�_�5�����2���H��'O\q[��ht�J���N�^���y�m�^�t������yf\����(V��Ĭ�|iR�+^�c��mR�^�3����_z�n�d�%�9+z��yO��V�����?��8u=�8 (�"YHU�/���K�����{s|`��̧٤9.հ%�{�F�C���U�FDe��9?�G���X2�!H)�ޑ�C4O�.�f
�K���=bѝ�x �����I%�QM=%�1������L��f9o���0�6�:?���`����.��ʐ�������6?P��yw�v	�dk��S �U�"\v'�M'��=�\��@�(�x��ciF�˻/5��w�HA&��/�}���z���s�s��e�P�� #Kw���b�V�
�w�{����$���`=��
՟(2�m���
���y��GVq���ԅ���։�f����z��V�����(�u���.F_S�a���T�w/V^∅�{��Hi ����ǵi�27�e�n�VPc~�O��$kL[JJpy���]�:O�A(����ßO(���P��'5�	�C�o����bb��s9�����DDߧ���eIL1�/I�/,w]��&F�v�)O��bk��L�l
��빓�v��1!�;p�?�
��/��zA�qnX��)fdl}�����6?�M\�|4��ܖ���@�>%o�D��U�\~�� uR���נxt��K՞-��� Z��l�����p�n�_�X�"��pmN{l����	V�Ɨ!s��]�eX��Z��z�`�ie����-O�:'3O����,y�^
�=����k�z?S��5��hk	Mp�(en��&5[Oj�J�_N���wڵ�4��p90�X�Dy����$͏Ȳ��Hځ�KkS�(�³d�C �jU�	��=>���']&e��kג�PW���Vhi'��2X9�������g��<0�uڽ�?b����:L�E��.�Wq��b*�Hk��nK`�*l�4�KԜ	G��>p[�eU�N�ȱ���/�|$��o����]�8�*�K�[}^�ܽř�?���8�yk�n��dfnſq��S�C���'�<���-q�#�������?G��'�l��&�����)0Q�/��nD�OL�:ú�*^�����'��a�ۇ1�j�e?�S3�Y�Qޮ���n�Ere�]��Y����[�]Et�Ջ����O`�H� }T�\}��]�-�N/�k�\�C�H�%g��I��?��� �<8>ܲ��T�˱Z��-`KI?��('gD=1%1Y�G�� � ^�
�����Bʃ}������g�n��HP�j��.�� ���K��(��ɂ=�s�Ș:��^��^��%�^��o��L�	]���!_�2amݠ����Di:���`Ӥ"�����u`�D��=w1Kk_;����$��d����+�6�z�%pV�h5�J K�w���!�Γ�i^����~cm���@Ysc�9�������Xo�v�S��A�^$����Yg`u��fF��"岄ÛwF�ʦ��ڗ�uu�f`Ԃ���)j��C�Kp���V���T/�M��x��
&E{�t&�>2pmS�e�LVt��a?%�6Tț����]*[�"���� ��fQ(��R��>W�T-�_�%$=��Ҿ�D��>߰�G��Q�cwx|:��q؍rmF��ۓё6�]@��4�@��jn�ئ��B�/�!j�<쥠�����ౡۀ�jb�l�).�5�k^~�M:�QMe��!�4"0-:�?E�A[�0��YfVhDo�.W����5��`C6+L��$�B~g��:pM�W�h�B�T���3*3�Q9Jc��G������?m�a#���^<�0¦b�Zf^t�N�-�x��ݹg�P�&�xy�x���!����괻m<>�QYs�Kk�E�ʍ��0���yi�P�$�$3Z�c�=/����t(��Q��t^*h��P9$��4m��0^/��--�#�����̹�� ���*��|�(P^�+8��ki�u�G{�v����XzD{�d�49�ρ���YN�?��5��ü6�{���J�e̴0�mVcV<N1�r2�gio�R�����[��\�/^�(�^���n�?:&,{���6��6�J�9��nr㦥F%���ќ�pl�N �,�$���l�_QC�R��5-�5Y�9F���s���:���kh?A�����h���FCX�
��zR��/t�Jjq�
�Ӊ��N~�ѥ��	�{'َm��+�+��W�E��p��CI���LYr���+s�	���p���R �~����>b�LY�Y�I��Ec��`�[�ΑTy��c�V5{�$���2����.�rj?�9�bIsY�]�������pv�KE���@#���Ԩ�r'(�����?�{�}{sf�`x��vc\�W���/�>�X������N�-�����ĺ:ݟ�"�}�t܁Y�����W�! �P��_��h�Gŗ<��`��v�M�❑����8��c2���ԁOR�	�x�����;DyF��Zt��8�ԕ��t?{�j�$�VD�b�*H?(���ʌm&�:�p$Y�u��	��<�c����Iǣ`P��q$zrT{�8% ��蔋��]'y�\���Ր��[�;��Y�.�;Ǎ��@	[�\� H퇴�	�H� �G�U(UZ�|%p�{��f�:��!��y����rPvT���Tp%�jQɿ�S���/�ˊq�0Zp�xt����\��A��)5���`��X�����@Uf��6��P�L�ʿ��Ժ&ϲ���By��5�}U�^jq׭+	��`_�}
T���9�vt���������{f�I�T)�C+��(����ǊR�ɲH���L*�^h���y� ���Xp1rɼ!��14G��f����g8:�!�1�b9|#�f�
^��4�XRu-vde/	x�y��<��bڻ�gh|�Y:�1�u�Hq����;v~;<pJ,����C��&��f�JqrP;��YK>��w����偛�X������y4�BH�Puj���HX��gH�팍(h�W��$�&��;rX�O��:YJ._�si'�-�B9L��tնB�^^o���|�y� C[�z?�c%�A
��@�=I�?zV�(n�X�̚�aZ4E�H�~eǨ4�x�{mU���� \R���zS
�u�`�n8K�ahR��`�Ck����6>��1ߒ5��L���P��J}�}ur��3�XlKKݍ�8�g��@�6ʱij��������;�,�c���ա�ݦ ��?�0-��L&1��	�F����M[�d<kg9g����c��l�v��d�t>G�ڊ�0l�?�c�Q��&��Lz�r=��4�Q��� /��WᢅT�]�[��t\/�?r�{#�����h8����o�,���T�|�O�"�#W�?���v��:*#UFt� �[T�>;��5�xA����v/��8�Xd��&��AFO���~k����Qh�g̉�a��荼��m|��������1&[��׸07����?�� �ԑ��K�� =�O�T�:|��4L:B40"RSZ�/�Q�tiP��,Vz��=hի=Z-&(j�Z�=a!�ʊ�����8�m+~2ht�JJ�4rϴ�=[i�1&�RM΋�����!�*)��?H/�5\�c�_�g:S��9DJ��6�Cf􄣹=��c�k���UDB���8mi:,�(Sw��] �����5�r��>!�^�v;ͅ�z�����zT
���<�'ZzJ���X���;��
^ω�}�M����h ?&!�*Пi���VT��PW���f���x_�ca��~�TX�&z���Gbk�0ڭw��+�Q�)�GL=e���l�d�&�^��],\о{H�L�ɝ<p�.�@���f�"����T�^���K�(�U?�S$̈I��H�<�>���B�ѽ��}�!4F7y8��I��C*Z�ʊ��Ji%�R��~Q/�P��}W��!~�#U2��츓����R�Ϋ�[ny�o� �p�(�;�2�iƹ�4�� d`YB��J/ߎi(-�y8��Y���T0��ܘq.�-���*��O�g0��'��M�E=�)�uX�*yur;*�;��c<
m
\�og�}����?z��L�� g�8h��q�[~��ńb�.K��T�ZӢ��"�b����\+B�Β�� �:�AQh�E�I����E�`��p`?'��Ԅy^Ww@W�CX�lH9?h=���/���ce�>`,�!�k��)�f����*�3O�Dl��ԓA6Q<�=E4�d*y<�����׈T�am�jii�ɣ�	xr7���-�8'���G��bp���jT��%u`/G�R�.��a�����$=���È\"Ӕ�2Q�*(��h�f�|,g��zŸI�!\����	�ܺz�䦉��2�L�R��_M_���ن��	�
�He�䈒y�����B��1�s�)��`6�FN�����pqB�5�kj�r�Ϩ��#�5܎�8J�N�i��+!�T�e�#��f����Z���������������P� ��q��G��V��i����*����qXd�b��: ���jxG�f��I��x�~���G�>�S[ܤ1����U;45�{Bz8����;(8M�����!)�G�D�B��@����y��~��S�z��&oCnRt�G����'.�q PК���4!(��?m_ ����H��:>n���P���j=ł�j|�$cB�x�I�2���-���ݰS���%��vNgc[ZGj���2� +.Cw//��.*�! �ic@���E�}�΁����&��x�	���E�<��A����5�T�,<��j� ����z펁F�D��An��Ls�?��� Hb��|\](�"�Crd����)e+Jp�����ߝ�f�V'�%)~55�ߵ�������l���>�G��ck^���G���Rs*T�$�Ck��7��^��>�r�`#cO	���+�2��h�>]����iH)N��aɝ�YM�B��K����2�d�Э82�$�툭d�aY��ȿsq������@��Q��u��R��]� ��'/�heHA�X@�#���E�R�]�7��WZt�V�E@�_F��Bc�W�I�S�!�L���}ן��u�I6�U�����Q}�y�?�B��J�Lɛ��5 Vr�;�-��-x��?��~qNe~�_�YR��KP>μ��%�U��`_x�������d5�1�|�>�7T�Ό��/���� �})XT��^����t�A����x��l�G��>o���b� ��ꌙ/ǳA��z��̏Te>���2a�轆��Q�Iz}�*oza�54���o
����O"��������tv��)%��n>pIB��a��)Nr��{=D����PZ���d�P��p[�o�QFBڍ�tЉ��}����q��$�2g5=Sx�|V��	��DuOa�Pe�:�E��.�1�iU'=����;����r�S��H������_�BX��u��{X�[��#|����*��]�^�C����P >����J� ��Z̦�ʈ4B���/�T��O�#9�8���'�7ۺTl7�o)[Iȴ��;SϫxD���J�����h�-z�.|�Y�]3�ڊKʦQDVۍ����e��M�ƺ-�7T�a�Sc��z|�*�XB����]�A��r��ʋD|10�/J� ��{�����A5��r�o��,�{��8]�z{9�n�����,�fփ�A�I��,�W/�8����g�4�r�Ά��y��0"�3�(��Ow�I�ֳ�����KƖ�/����!>,-����gy��A�"���ki�#v�Xr8�N�X���CZ���iШ����$i]�x��/=����:�$�D=++'���*�� ͧ{Ɖ|幩1�rSp��Q��3�oJpb��mI"�,��q�³ĥ������h6P�VRګrxgA���l����O$�[-�]�1Ju��L7_���r����I�YK�V�����@K�{�K#���Z��pf''��Cze��传�O�-�q��N6?��@��}�J6qRT��C��y��d�}�*y�j�yG�j�b(:01���f�?@���^gROt��� �+� /�� D���	Y�ԅI��~���w��}6�����u�1G�l���TQ_3L,��5�J�5�}�Mn�[%Zjp�\QL��k(��!^��%Jq�{�km��_!@�G��sԙ߉׆#�v狶m;a����@nu��35��3@�Y���r��>����RM�Ǧ�D�-��b3���K�T�+'�����¢�O1o���}��"���׃���a2J���>�h���I(���=53����]�f��U&v �f$��"(�H��&gqo/Z�t��sa�Do��K���.�ĈI�i7#����k��9d"�B<u�J¶~/O&�̋��T3��:�͟��Mzخ��i�n$2V��',���S�@���?Ȓ`�,9�!�h6�pI)K���=ʁ���A��2��sPI��@�E]L��+n�{ �1�+0ۦv��ǹ��j����_pp�B� 8d�U���l����,���m��n���P�t��
8��} 
�R�٬���x�]��S�[�����`�@�P3�Ed{�l�Jr�5y�s;P_"���v9"��ZH�h��@�Rl����=��K"]y��>�W�zn]u0�����e�g�_�R�\&�t�#������Y%���)oԠEޘW�v�G�ͳ��iG�/��H�[��Y,��]�!����&^_7НQ7��=�d���C�����G�QM4)F�h���rrDz�l���Jo���+�/"b��*b��On �q�Vǧ����%�U�G�;��X�h�<g���'�z��Ŕ$Z���7����	<j�{���Vc�Y>�Щ5����u��ID!H���X1w@ϓa��՜���X<.Jr��}�@��N�A����00�h�)&v68�O�mӽx�?�7�#܇��3*~��P3�c�%v� �!����Qn�#�}H��L_{Ę��1�^��<�e�b��WR�h-7Sw��2Z,��v����܂U:!��eڡCp9�h�����N�\g�w���:�B�C�Zb^ i���v��9,�5�l/��k���Ӆ��mK M{���d���{%���|�}�7O@�k<ki"k�$k2)*�"}�{���t�/�/�"s��\+�5����hd乚y��$s0l�^?�B�8&L��f���s�z�B���z_���Q��ׄ��ֽ�ѵqS9�f���>���3�D{��K�J��}p��ظ�O*������k[{�8�dDiه-����3g��z;�c�.?�Z���i��F��?�X�}g������+t$氏���''e��6���nG���;i5�uQ�'�ڤk뷅��
M���4���H�/34��{�\(�3�PV�4ґg['�F�N3��X)d��9�;W�R�$W�Ö�!`�@
22��"droE߾g'<1.&uPƎ�|.ߒ��БI�U9�i`l���C�
؅���@��s�;>�s��1Ai)��ط��y�mPEN�A�lf'/�S�����ų~�fSH���#X��Ƽ��R� _����>�d���t�c�a���C�e5ds��\ňD��ڸ{y�Ow�I�d�e0�>@?ǰ��WiF����!��p8��e� ���<oȲ,�����:�U*<?!g��c�]E��lƘ8�
�e�4�S�OH�$w: �6> �n�L�G�Y	?O5\��0���'P2�0{�N
��-�"�@Dh�D��/�s[�S#�u���m��n"���~��]�"�}n��Z�i�"��ߝ	x+��-Rt|�&�ܘ�
ֹ�`�Vis�|�o�����3	��.q���l �?t�Z��C���ٝ���q��/\׳s�uq�a��g�
�2�ʯp�c�O��7iN	wwܨ���$K.9�!�ͮ��݊��c���c���x?e�dN��4"�47N��))0X�6����[FX_��;�&�:�.���-Q1A!|?Z����v��	f�HP�.Vd�g�UkL�܏���/wQ���뽗h�ǕMjR)���Q��K�R+e��bzʬ�Gw���׶��]3�	��������R���t힬W6ֺ���7b*����I��a;Uq#����*x�����ź�M`�Ul�D��J�-=�x����8�P�)o�)��!�Ό���G��A�U5�V�lϠ��G��W��[�������=T/��QkJ�Yl��j��i~a�cZė�δ�)�T CKݑd�MB��U'��s��� ��y�7MN�Z&����=�V�R�%n$f�����9G�T��'�x2�K���[�F|~����x��7��C�Ǳ�G��s�Y��/�NVLt��ca��jN�y�a<�/5�y49�x�2�U49��5�V�P������R<}�L���}�W�'����j���c-�_���~'U��<z�c���+�|��/\k�`�U�HҳA*�N/w��T��=�ނ<.�9�}KA��k�(q��ʟz����H�W\��+?}^�`#�ߕI8�em��W'%T1G!���}����qc���qJ�.���u7e�3���,4Ck��gc�����������n�������<�Zc�b�57�c�cC[m�-����Y���Ƭ��!/u3°Zg���\uLS\c�w�h�HQ��)G���{�C�:SZ��Fr��3l�*�"�3L[���g^��l�c����W�Ј�e��=ګ�$&_1�*XІ��"�{>zǎ�$�����L=|(���8RI�����2�J�a��`j��{�[D���@��(O�b��y@&{�vKr5k6�A�#E��b�eM�Mm���&���G�3�u1q��{����FXCr�B����O��t&\�Ϝ��K�ޛ��q�$˴��i�w��tM6@؂�Ud��NZ.�h�|���l���	 �^S��M�f����7�l�,Ȉ�|�� ���X�ꔾT{L��������F��s��@$m	�g{� ���ㄡxºsr~'Vg������#b��� y<]�.	�zv��G����>�nγm�� �>iM�Syd��t��T�c{���ru�[{��c28�!>7"�r���t��)#z��X�� '����ÿC{�zq��\�V�Nk��]���G�t����\����o��L��xS���C�f�U�x�ҿ�+��ul4"�:�ܲ)k����v拠�;<���R�T���=0;�:��$8�a��J �JwE�2���l�Je�a&J�K��͔�]'�a�S)�"o�5o��Fg��ZcF��W4&M$������}��_$y`�ۃ�t͸���x���m�b�Ա�U��c���Y��-ze<�4j�)��d�mՕ�<����<��4�I~��V��V{x'��n�~��*�����S�$�M���:�O3�T�k����9���]�)�b7���F
Q ��µ��x��N����"4 Y���R{�'�d���d���8/���{@��M���غ9���%������{���{�^V��k�{�7�i�*�%��M�vP�P2��饛��
vO�I�1�P��Ya.u���}�H72�ԕF���Ex	�����_?jX�NJ��cj��|���T�O.���V	7b�DW��:nR/Lۈ��9�B#�r�
��%τ���Q��dN'jɬ��P�	kا�����}�zL>ܴ�FP��Fzp����A�l*6�Ee�:�_� ��n����tj:��},U�.�F��Y��TA�����(��iB
�T)�~��q>���w���~�z����%A���~��I<7l�ֻ��-���mB����|���G�|vpb�s�я~��`@QJ�^��+�۹�	CQ#`J��R_�եh�`<�� ?�4���U��y�b��@�Nmp��d��%��O�ټ��۲�ٌ�f��t�f��ң���n�i����0�i{��1UY�mi������0���x �C��ְľD5(H���D�tY��p:x�W�O_Y	_��w�mN�%���^��hǤ5�r�_��1D^X�}G�/v�F���ؓni��v�#���V���)z6o@B�u[����!�"��X%��([A�͹���{�3�Ϊ�\�u5<��d�0��Z�-�����%�5�*���#~?��`5�M�qh�^F��`���#T�W�?���5��L���#��3�K��� v ��kQ�9Y h[�B�.�b7���(��w!�(�F�bO�l;�t�����]�?��Pc4����Q�L��){�|����0g�=+_�I����y��_3���{���o^�#Il]q�T��Zwof��>���z	���a�cW�o�耋�LPщlC|N���e[����|����K{�D��+� �u�\�V���y��f�"F<au<� �;5�F:�s��}��e�`?Q�9p5L�aGx�#���`�T�W��pq���4�"���D�d}�g�E�G�Q%P�-�4�KOs�/�
~���� 3F���#�h{��jOEo��X���@Sx�I��'{�����T�y�!�^�s�lѹ�㤉\q��N��E�І�Y�r'X��[�Nw�3��E�gkS�/%1D]J�G{ͅ@'z�	1�����-A���g �|(K��4?nB�d<$̞��]��:4	l\&ֱ���mpsy���1��AX�uc���6:;>:��@-z�NKe=��0��U���}���X�^tRKb���IC(-�3z3gDhO�����k�-Ϧ��W,�&�o�O>�(���M���k����� ��(5�u������N�������{�f���@2Ma�w���kg���תW˹�>���Hc�5擱cF8� ?8Xj5%	��Iw�/���s;4��?��a���-��0b��e4����5����9��b,\�]1�Bc�)��/��ܜ��z9�0��5K�GN$@%þ�(~�{_#��������j�i\��VÃ �~�c����e+��W%hB�ޭH��W�A/TL�	�3�/$�ۤ��*Z���D.I�8q�>�(�;3��Z����-硅�eKwo����2����}��T=���,�H|�?Y
gio�9(�+dq�n��s��c��P�e�5?��U��tot��'��ʎ�T�q]j�/�r9��"lDD�T���%�ᣥ�	=_�9�O9���`�s�?�"�1�M���h��M�EO��N�8��Z�Q���S��!�W�����ǹ��c��N�A9�|�c��K\�,�5�ү���X��{J��>-�W�	�
�צ��\�{���\�\� �����Н���<��fv�Ly�N��Xf��kX�c��¦�@��/;�<�;�P�V�3����=ق1�	��f����������j�n�-�g���ׯ��A�AE8w��_�u�F��D�ww�������pqR����A��^��5�D�<{��_�h�vv�@��L�״)�:����p��Z�"o�iT���,�}O�F��薎����2�Ds�iwA�X�4qV/�u�.�2��l([b��F����y:sa�������e�EU8���6f}u�vہ�����]�����)�W7�}�#2@��vS��\��� �r���6Ċ��+�_�&4��/4,��|�eQc!Ui�B�3���5ݱ�Us�b�q$YG�dR��l�}�>ٞ��ԾƋN�6�(���5WLt�Y�媞���d�W�$�2��{���aJ78Ɵ�:��F�>(MC��f7)�9h���.��k��i�f݈Δr<,p��Lz�2�0ixeCO��37x�q4ŀV��ӭ)�^�&-�b^E-vR���N�������^��g`��[\t�#L�f6���k�L�,d�y2/�t��ȡ��{u	#}�7S3�\
�kHZ�r"�r3|�Zm�G!|�9�r�`��N���q������X�1߀T����Ss}��D��,/��b�f�1hY{ n���'����.�D��Α���b��ʗA��n��.�����3M!���f����΂f��b�ǻ�V�,15I�������IV@N���n�HF'�����J�#I��Ƚ�������Z�J]��I?sBꌩJ�P�vsZ~��-�W�'�k&'�x$F�gj4m�t��P�a�;�k�g�/���i�������)K�]y�U���>wcyI�֙4Q�߾��Pnqe�x���w8�c$�^��%B���E2?��{���ty��ZbUY��ed=H���J�'j�A�����7�A�?�;ۺ�ԉt��;OK��@c]�ϫ�['ĩ�T,�F/��*%,q9|��:���q�ᒺ�d0�
��������ŕ���t��I��N+.kO|lh�<מ�E�S0��6��S'����ݠg���c��<�t�eu'�{�|���v��c���zx,�b�=�ʗ�	,�j��Ĥ�{�#9~�3�j�M��3�!�J� ҞP�"�d��d��t:2n*H��D �7�j��N>�h�l�M��}�Ü>�����u�,���0yzo�x_� ��vj��W$����{�b;t�ɔ`BT@�r���=���ZkV���Z��=�Y8�P��&{t=��uw��(����4�t��&�R5c`�,�8�H]�6F���T���&��8���pv���^N�b��rHc�߱Pj��|*8�oF��8��Vͮ3�V��F�u���%�];�NZιj1�s#�jx�Kz5&��n� �:��[�A�T�R�L��T?H�}-}�b�����qs?�]��DG9K�;<2A�7\�Z9�,]i&� IA��Y~i��pO��X�eJW�K������$�,@S�)�8��`$�T�K,�ٚ���v�FF�.�e��*��;{�Q���ê�J��k�  4[}W��Xw%���x^xj�u{sʍ� >'V�T�*�F^��s;�aP�if�: p;acw�Q$�T�!���v��/�σS�^��Z�٧�4�u�e@*%.|����q�����W��a}���OP��P����լ�!��C¥_��u:>5��Q{�!���B�u4.=ޤZ<������#��ՐG8���\ � IsȬ�����@�q:�h5�Ͻƭa�76��v��!���9��oU���/�w=�"�﷫�:��@��bh�<�{��(W�`�B�RYD��DI�?	�b��8����܎B3�ϫk�mȴh���<�]�7�����H���B#�k�R�f�.|N!�ըe��w�*R)�#p����S�
ؗ�'��d����iG���?��Y�����R��U�~$�*������k#Pt	�!�1�:��@ Ւ��P�A{^~	��f(�/�ڣ���m9
�\��u��n �놽��)�������a�Aj��Țբ�4���%��M�w!͂��j
e�[����á }?�T`}�/�29���c����zW���<DK��G,5�C���]�k|;C��j 5�)l��q��B�M���Ý��������˘�<��S�$�5�C�x_[�!x
���R��*:�w7H`�#�]����������Fr#�N�u�S%���fCtJ<��E`�YnȽ�Oa֤^ܶy~Pb�����y��k�,�e���rJ��d�͞�gj"FE�7��@�������yF\�)fu�����c~
���{�O0u�Ϯ?��Ae����d�)^�z���r/��$��O�̀3$x/{R���0�l��\@h�u[�D�*��j���r��T�l���*U�jR�kʻÁ�����.��������4��է�z
��d6l�Y�0�T�1�Կ����IW�2D�M:�ӥ9�%f-J�" ER:��T��N:�V�0�"��;����8t���_�͗�R���)�&e=�ArOJ�a�4���ٚNp�r��y�J@�X#r�JZ�K%���)���|�ZQ��Eb�/�d�$��D]�>��;�͇,��*�����4}&��;����x�v��QY�;�����m�:�Tĩl�o�~��� ��2�n����o<9�N@qVh-�rC��2�T�	򀂗
h ��I��E���H�Q�cN&�������Y@QX]��Nc-q�
g Di���s\t�B��Y��p:s����G��jx���B.~1��}^�y.�#�ϟŇ��
�*ڈ��:�P�u;��EU��ޠ�޸��9z��o����G��'��t_�����	f�w6G�e�o h��I���{L�VS�lOL�B!޺l/nT��*�Y�7Ny�Oť����g\	niY�0^�K��_Տ?4Ke/dl��?蛳�&����#�P����p�d�)kA=����վ~�0r��g��2x�/�*8�ݘ�)��6 ��o�ɣ����o+��6�M�ɩȓF2�J�T��A�D����k����U�3ߪY�Q��}�R�m@Y�X�E��l�����3��o�� ;�$7Aqz�r�,Dd$��=�"/ݸ���,.GC���is�wN�ߊxKBRP�<��p�5���'J���Fސ��A4����Se�.l,}�H��	�HǁC 7�C��!��d���˷$8m�|�3D��	�/�&a������p"���ܔ�|8�0ij��-˙|��ﱰCaD��a*��ڗ(�I�q�Ϻ�����9HÕ���Nķ�p$�����Qo��_�o��Wߧi#_W"�ڞn6J����x"�xz���a�ցP�OXƱ�$�K�!1�&q�B��S
p1L�\(p@o����bm#&`�uG>�yA�k�igk!��H������Z��5�x�ͬJ�:p<4�:X��K�X�d��OC�����Ĥ�`$uQ�}��SB�[��=S]�4�uP�A6�r�~��haWq5A���E:�B�?;#�kgA�RMj�byY1�������@��'�SM6�
n��/���,�ƞ_Ԗ<�>���l'X�>k_-lʤqH��|��:�n��z�)�+x�G)�d�.@a�9JEa�,�&!&��?k��YB����|�����5����-P#P��l#��`��=�@��e������\?��(��W� �o������f���I:��0Х��47���x��Mw����M����&y���y�١;訸ע~2Z582�����PD%��KI��:+���W��[�/�g�E�@*ɢ���6<:4Z����CdۭP`@%Bu.�7]3W�;Ʀ���CyA}��^3���;�?��ؒpSA�����|����!��� ��<T�c�՞e��9+�Zx��_�L��u.m��+k��+��q�M����IZ5E.py�/�QI����F���v�FXXFh���w��[��tY���\��KX8\/p�*.q/i��hp��qj!���kߤ��E��ϸE�Rk��L�~c�{O���BG`��^�r�eS>}"#��\ˡ)7���i�9"�6|F���f�SN��O"W��3l)�`uOӷ���6�Zb��I8�(݇b��u5�b+��t��a��]��zl����h-�9xp�б��`:�n�-v^߸�Զ���S�{�1���y����>8/��Ҳq�^h��5/-�1̚ԫ5�V�㬼�[�H�f���-u�r�=i@m�Y:�Bi�j���κ�+�S�ǫ����䕠�:y�(�?=��#v��v+�2zB%L���)*ɻz�E1�6�x�2\�Q�8�A��V��bJ��M��jP*Q� �k��ߢyrp���N?�=)�ebf[^oW5�����E����D�A-�tX�$�-���@L1),��n
�0�B(}���<��׫���YX���,�θ[p�K���d�<���ލ<l��p����R��`����.���GD \��AC��f����?�u�_���f̦~�Y?F��Lu�f〾�-���=�Q�h��1ӄ��,M��-ގ/l[�&���q6���VL}����e��A�w���yzAM�V�{'��~��Ԡ6�Z�O�R*�^|&�	�Q*�h�Z���f;l�T�`9f��a-7Z���r5c�>�G�by`P[�w�x3�4y9`p���I��T��[7��Б��'�
0�li�_��n���d��|�QWf��"�(�vE��]���u�>�zmzv����@���q6�ڳ쨽oL�<�o�u[��-t"b��1?3�s6}f BY&;�:���`L�=-i3*�7A���]�t�'i�u�*\{eT#3�A{{�Du ;Nֳ�X�{HH�[oV��Ҍ��$n�%/��Y�c���X�fɔ%�ے�vb����^�4�>O�z)����<))(2��%a��@������T�W������+m��8YG�-4�f�W��q���Kp�v��`*uyVA�aJ�5��u�Q;F�k�R�ñ���"~������.1�,����h�3�Q����$��"֙���K�{U�@3�Q*ê >5Z�4�J)�"4~�㾃��I�+� �m0? }ڽ�����I:8r�|s��iࣆ��N�uhH�elj4R�Q��=r��l� ���G�-/@�`,?�îj��֣��������7%�@5z����)c�	�Ѭ���Y&���R�P���������s:X��V�$ܲL��`�}� ���s��e���3�$&�p�|�gYK��._E?݄��xi^#�m���6��e}e>��������;@��Wɭ>� RF5R(I�����67�N��\sQ#QV$2�>��BV���dړ�v���%��:�9�[�i������_}�W?�HG4��n�f*fG�H�i�����4�!�3vb0�� �4W�η��iSt��J���S�1�3����;�Ɗo��U^�U��4���e4y�����F�Ht��ryw5� Wz���UY�I~�>��R:$�p�����;�b&d69#	��NQ砙�j�����:��$D���9��ePU�$Fss�z8�29ek��l���ay�+����w��Y��ah>%����tL�Eu]�lJ�ݸ?��N�n����1��M�=	�s���`.���'�]w�W��p�wҭ!+v�����21�j���l#���7��ӿMݔ�a@���._>M��<��	?g����V)\-�D�w��u]�\����