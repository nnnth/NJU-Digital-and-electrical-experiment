��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��X[&-����v|��y���RI�hm<Pi��yT8k[���0��t._��B�k���و:of��A�v��	�d�4��,�5M.W0BL�PZ�����˄��:��.t*�Ddh�F8h�+��s�ϣ2���<�r��J�M��ɞ�6�$�� i��V�$�bT��~��v�Q%�|��+�����B�(���?*��cI�7�C���BA��ڌ�<����vC䖂�x�z��	��L.`nh�)s���khh;�gE\�4x�_|F5Z����ʦ��ح2��������e���ۮ�s��Q�S:��H�E/e��1�����!�7�\�rlHC�bxn�,h���)N�`��a3��訖�(�g?�P�l`�dv����vX��{����e�i��şT��o(s��k���S�����N�����e��4ժu�+5�^�T��5+����@�yT�O���+���xF-"ZT��tQ /B�N��U����m�;u�~둎���M���ؗ-'�|�Q(xV�5�:t1�7e'���d7*�bi�>1�����oD'�R��R���"Bk-���7tA��7�'�o� *�&%���e���w4�5疍�gW��')1�Xq�G����o��� 垃��,�exL�/I��Ȓ��h���׳�Y��rmv������4�r?e*3;j�b���=�.�ʉL��J��{����w�_�g֣��f�?E��VH�@�[fa�Ir.�W�#X���Hdwp�����$�؋sB�qa���u�,�>���a�/��a�?�ĂAA0�}ʐV��>'��ޠH���Cg3���k:ie���d?�*����-h�Sv5n�g��Z��,��F)�*��F�4�R��G- V���osk��5jtW�ø[���Y����b�[�U��Z(���E�M
�1^Hh�C[�kѩn��{�vQ�燐<^;��Z�9�'#V}��^:����ߢ�j��
����UZ*�C�y~a}��[�W��c�D���LB�w�Q���W���s��c�+��DM�({�K�廒��߮��Q�N�ݢ3It��R����H�"x^W�۬�>�۪
 Xh�¼�<P�I�k�.\�$b �r��4��na�_G�%V.R��ⳮ,�t�J��@3�a�5�0T^�ߍ��E��[��;�j��I:����g�y�wds\���'�+== (�0�@�1�?Br�fZ@�Q��u?�.��r�2����t�eF=�n���W�0�:#!�&iۯg��:>��~��$�)!�7@4�40p+O �!�`����ٵ0gz��
�X�@����EmD��=��>�g�S䅳�&��˨��Qa�o�m�3����������8?5'��Da�y��*�܏bm��7Q���]�� �g���B(;O2P��(�Ê��:�����d@_�c���~e,1�&<m9�D5ky�d��v��y�I��Ϝ@�1�4��N	;x0����Ü�%i�R��x���=8��\O��}h�8З)/y�αyÑ��;�"���"�跪���\p�����ֺ��uUA>bC+���3hh^q�J#����gʄDF�ŀ���[$Cy�btrǆ?�qrM�:���Ԧ��&=�3�%H�����>���ʨ�#�9��11p����Lw\4d3XK�tZ�WO���k E��؍�śu��;���%F�#�����u3��j�r�@��xe�f�"&$b%��+�a�����jZ��aA������l[�;��}��DݶNdM.�$��`g{�Uk�cT��C�ʫi�A� +��1b�����b����z.� B��@�
K~Ɉ��� 8�h� սwm�q��m~n"a�W=F�?^2U���TL#��ߗ� �4���3D��>��O�ڼ�&밖�?��S����t�9�ގ��	Ǎ�um��'���/��T��=+܎�����U��m4x�"4�&{�/�(l�{#��r|��2���KW)�U��wX�5�+F�h�����?�l���/%���m�<伅^%�Z0}e��Bե~�l��S�!�F����»�a ��>o���u��;�Q`���(�=_��L�Æw��ϗ���SzlCe�U3g��A�oj�#Ik�ڽ#��|�_m��/�"6��_%V���]a�_�y�h""��iq��-r�tPw�H/r��mP3:�F��h���f��B1 �
,�I�M�5�u�����F�)�j���M۞'��WJ�X�S
)�DG���W���vR�dZM����I=	- �"��Ij�Ce��x�04�� ±z�h*��G�E]p��d��#�W��P`KuMD��7�ְT=EY�M��\c���D�HZp*i�����$������ l7�vʇ����"{+|��11s�M���s�0�%�i.P�7���d��_�������%@���@q�#���{��@EQ����u�}�m��?׍w@��������1~�Z�9f�/ �;S���%�j֬p�ч�N{�׀|�1(��J׵|AW���Ĥ�-�"�5�l��Ipn�G_�@dP�,����/aZ&�oƀ�6���&�|*��"h��#l������X	�x'"����
��)�f0stC/s��iC�c�k���w��� R?슶����,80r������ ����k:K�Zf,��3��vӃ�}㢼�$c4� ��r�w�^>��>C��]`e�,��D_���>/�h~׮Q{��^O�C����*�����/o�#�ԗM�S
h5��dEU�s��������0��Vw�؄��t$a'�﨩,�	`�r�@�σ)��"Ih���a��
�+�t��W�F@'�$�z��8��O��Zkf�I�������.�Tn��}��ܛ~�[�"(��͋�C��.��-���;���d���xM}�}�Z@h���1sD�4P��4��E�dT���9�,2180�-6r�,@�*�LO�c8�rW?�C�C�����껓�C{��$��2b��M��3��'/�~�;�2ң
)o�&�A��OsPj�OF���_��@�������x1[��_�E���>��!I9V�mS[�p�J8������~�T:�+���c|@	ȕ#T��&?=hW��ܨ��1��{_Ѫg2���mEp�Y���x5���+���ڸҹ���O��W�vFQ0�F,�V����^�ϴ� !���I<V)�u���3������)T�?':��$W�"�]�Xa���=��!A�A���o�U/= ���+�~�C@Q�}�Lr�%ke���	>mX>p�A���P+r��s~��<��@I�>{���4e�qy�GtD�Z���&��� +�u��6���7k�;�S�d� �:c�<��z��-�)������
�j�����W�>���$+��"%�I�k���yt3J���"�t����	D.܌,~1ۅ~3���y���2�C�J!�G4k(���	�G����q�*��עi�����8�_l�LY>�{H�l9�c)�0H��`W����D(�}){�#�?�+�c��WY{ܷ��68�?^$��łM�(|z�\�j?>� ��vI��Wwn�(I�y�� ��������oϱ{����ujʰ�%��>lGt����o��Ts%E;�{)Un�E���p�u6l�;ҵ}�mMR�M\�n?~5�52u���p��4;8�M����_����@�9>56<�_蟽�F�:���_��_��ш��uySgG��=ǧw�����l��3FI�6dJ
�`j9gV�s�C:�E�]W��B���~����P�磬�� PO��'�w=iW���^)���
�;�{�v�n��� �t����bk�$��%�Kh��.��3�e�ï Ibn��x���0�k��>h��%���~48���[쯵R�vb�KΈ[��p?��*�e�]C^��ƀT��KH����h��n��+~��Lk��AJ��Jڽ�g�p1��e�_̸ܠ��yW�^�z�UǪ���(8$�.�-0qN���PN2���za/؄gna%�֪�_F!�n{�5�������r���
	���ߖ���ޱ�����X��l��s��@U���p�����6LҚ`�����E����ɕ�����5V�s)A��b���Val��!k>����G�]Y�
r+KZW���݀�(��C��	��z2�;�XJgH���/&�����9�i�X���'����ӂ�:����|����q��^$,"�� �cr�㓟���X\������+��H ��HƑ�I����YH�ļUM�v��_H��f~R���M+C����+Yh��7=%�e����n�օ�X��@�J\�t��/�ZJ��.��-U��g�U`��i�{��ߣʨ�G4w ��Uκ'M��%��,F�EY,��s���U��� ~��Oe>��<Ʌȫtť�!�l��.�S̨�1К�����l�س�k۷�p�^�F�K$3����G/"��u��V#�DJ���P��;��u���:���&�s.�ԚpС!� �ڪ��a:WG{�ރ`�4�F�S�>jC�.!@p�Ⴇ�Oڌ^b-2pD�I�Y�F�O%7���"<_,ʪ��wX[
�Ƀ�b�j�M���y�є0l̅Q]��}op?h:G���s.-��(bjrJb+�L����ښo�e��UudC���A��B��w�D��䩸$1�˺�c]}��`i+����$��f�KD�
�4c�����'"jFBKJ�̵rP"�%\�N*jQ5�Z�4i�Ϣ7�(���]n+֜ctu�)�mr�;ㆠ
lE�o�u��<�	Y����TpDY;����=��T�)�q"6t�B��j����?-��"��� �I� ΅%�Z��a5�ɘ:���k{{�4�?h@�ƏI�b^�Ք�͸C���j6"��m�@�nLA�!�'�~�O OE�.��^��x��v2�#�����G>�#~�2�q����s���0�=e?#FE��N�0� ��A8_��?�&�jg�ڛT(����]������Q�N,�p���)Z�኱ H���#K2��������٠���0��,�$	~B�S��y
��ǄZB����������Ln�u���!k��� �g�לOB��+�ڤ)��F~�_kvNr����
Wi*�?�������E��Y��4k{+�U��h�>;�zg �/N5�6	�g�N�)܃#��I�����-�_�g3�/�)���k�������q���z2Y\�J�����@8lk��B��<-�"�ʳ�S�lc �]]��=o��b��>+Y�\�gj0���)�QXFkN��{xJȏѦ�C�'G�XN�&Gd��2թh�Y�Q�R��@ �1+�)b�޲z$�u���Ea��vo�
Z#80^���J�(8����"�׌�����Nk����	��IЮTQ��^�s�����߰U�.ߦh��$'m���}��;�Mt%�^bxu�Y�]ߗ�:+�#��J!3�j�3i�o�k�FoX�ZO���L�0G5�Dw��_�}"�t2����L��f�4ݠW\aB��i�g�f^��˵��W����B,�H�����	p*�K��̢���o�W���8���ǥ�4	/|-RE@ 5MZd�p�{�N�T꾞���W��D��v�su�)�R�鞝_��I���I
����L�7��}�y`�ĳ�P�
�Wj���Y\İ�t�%��MY��@��wh�[��0��܁Y+�3�Vo�-8�.>���y����a[�c���`�j��$��)/�*GQ���<�����w���RU\�	�E���~���â��m����C�B�F�#��Z�=M{��tқ�T� ��&�a�0��!���@u��3ϲ�l��έ�jQA���<����f�nh�=v?~U�{�Ȁd�5�e�P�T7
h���0��b wb��N��G_t�x�<�����^��$M��:HGj&o�d#/3w���'�����\OƹN:�*����,yދ��������c|o�N<3Dl͙�>��	�[�Ij؊t"N�����a����H�Xbp|�x�H�:���"���{��a*C��brQR�t�)'�@����N��t̔=8�A �e���P�zi��"m$�
����t|0���3�-5iu�ơ#;f�NXA��Z9D&�jd��bj~ѤjJx�Dhl����"��9E�в�ܰ����E�'�(�+���v��`�$��l����q�'5	.(�.�_���.�oğn�
d�$k�:C�l1����s+`��z�Rb:M�(PM�ڮ:��rc�^�]�9x��jn���iծ(#�d��<�P5}��0���HԪ���]��C��Y>�/� v^0`�t7�oU2��8g�p�?M���Z��|�u����`ó��p��4���{�CF��#�P�I1I�Ӄ�I������t$���{����Lh�:��Fm2��g�j��8��@����Sk��	�c'�S����M yQ�)�ǟ5�n	*�]#��i�i�v�Jv mES�7��̩�7e��՗O��L��zt�}%7��G�g�;2S��i��ԫ�OhР�ۦ	�:�"��:�gh�Vw�g����e����Z�~��({�;;l�z����I5w%OvZ㼁y���|H�uF��\+��]At�;�$BG��^�/���$ȗz�v��	kD�nޑ+�nȖ:���U2X�+�dZ e~�M�`�Exf6+u��|�쓿6�*��Z6�����nD.0�t��*����IG���凈��Q�jHc��@�3N�-;��N���a�O�� @�+��
 �%:`��ͤ;�G;*�C���E���|�:Yb�oT���,P~���b�D���8�.W�X>y7��<�Q����ڦ�`f�Ն�Ҫ�`�2�q��I���h�B�/�S�\�����1.�ܱk_qQ�3�?S筤���~���G\��فD�����Q|湓�~&�V'�}�a�z�����<}X]���eǋ3��[^Ye�9�.��9eK���"�!;�*�i�ն�@�QhloB�%u��%-�b�Y�l�~�ڔ��n�F���.;�a:�r�r�)sG	d<����wG��6������Yӆr�*���M+ߞD��&��dN�?�w3��x��,�
4#��i�.�N!�����K�3AT勁��]�w�"���d�����I�+�Z'��0���&!�[�WKЀ����!t������f��������R���S&�����pz���Uj4���L��&���j'dc���TZ�],J�q�q����O�j�+�lj���n皳����\;Ю�<�����"�L�ߗ����ͬ}S�kb������������j�
�u��Z��?��+�V���@��ɨ;6(@�Dm���P�|�Y���`nec�](5����h��t��N��u��I�qb�rg����<�FX���ΔE�^Z��4F�2I4Z��jp�3},(��k��5�i��ָx�\~��Ph�8��<�\Y��')�]j�g�l��x���� a���p���M9��DD�%���8sl��lG� ;e���h�ƛg|7o��H����exS�;L�����ic�X��/dE*���gK��]���N���N[��6��_C�X %�[�1��g`�n)�+;�������u��=�cx���|t�*0�)�8:��F���%J�c��U+[�g�6B���3ι9>I	ȑA�Q�����Yx���ొ��5����N���oss�C[��o���˕-��#H��|C y���߬����7�3�����$�	��a �sf��dv��dP�{_l�QN�����;TQ���L�j<�����o��� �us[�(���	���Y�`�p�Q%K�z?mI�Wk5�;4��
�����Ն�O�H�����N�]��3��z�H-(C�F@ln̂%�`��^�� \EQ� �%�z�X�=(���$bs��f}*:<N,���Q&R�(
ðN�a�Q����E���o����	y�No`
�{���GBm�͂�*�IVʪ��?ɟE�U�F`�gˊ7`�����)t�eB�t�p[��/	BV^,HzҰЫhBN�Y&VX�ԇ���ɇ�j2v�cuϷ�*�j�� C��`�"6���Ws|P䛃B����~?�(�k	j#����YWC5^�u�Ɇ!AHp�s�G+UԦ�#�s��;�P8[��?�w�U������N�@�3:W�?���'̙M#�(_n��0��6�@��j�4��w�g��
~\�vȻ M�:�m���n��9����z��� � ��uB��� ��m2�~��6=���(�=F� ��}�Q�m���|]����C��5�+71��#e�z\�|������/tH���ǌoi��o�^ӱ*�7s�x�*��4w��_Z.����O{��'GT֋B9�kܵ��ޟ��
>,t_O
��p�ͱ�}#H�m)�����-GdQ�T߂���"GMP��z���Q����r8*����J��)4�p��_�� �� ��ɟ#2i��ߛ?�hƢ�%�x�k�ߴ
�z�\j�>�*���+|X��*f�=�!�CK�VΉI&n&:��~Kown$�����Y5%��h���zv�02U�,�f�H�2	�y.Y�@���3ر�E��௃P��[�#5M����J+-L�\�V��7)�#�
�f_�'�_���D�5*�d�N���RI3��A�#���L�ބ�3�cB�k�>'�!��F��<z�[ry���O��8=����`ȢjAˎʐ؎�vN����^�̿��8���:������?��m�JQ~�%UZ$��5�Z�7��"�M9/)j���2Z����K;�[����|��� ���Lore!�z}�v>��,�f��x�b�TS)u��6�w �� �)�n^;:��%E�ζiha�$y�U&�[B�A`��/o�$W���nMN0��z�S��x2Mo˶Ĥ��0jy�? rk��|g͌��O�
�i��(JǱQ�C��Дf�QM9��9� �=-H�3��|�#s�n��RFq ���w"ÿ��UL T�e��?��E�O�_�U���/���T/�����yi�f�&��#��:%�Y�k	�xr���O�b��!�R(��W0҉���*B�c��7 �̍k`e�j�N��#ؔ<��*L�P�
0�0-�9=Egո=��g�$D�ȕ:@P��\B���/�] *���&K! �RE�t�r�������U�j���b>yy ᭈ��f�
�l����Z������U�v��ГDgj����}'��tɁ���3��[��c�kL�ͯ.nJ�fs���+3;��#Q�ʹA�6W�؅o��yְT)Xhe	��KOW��&�Uj�=G���ÿ
� @��9��<��/��@?�r�J�������(J��ޭ7M���9N���`����Д��T��^*�\�s�vG�qF����@� �V��\��p9fg�ᛉ���Cj�Ky�݁�R��5�L�s��L;d�,.����4�dC�p��6)��~"����}�����|@�M��� yomcT��'��oyr7�j ��Ny)Qd�0�Q��κ����&y��h�R�j��J���XL�j�'i��p�\�)��f�(�����P�0i;��wV�zc�{�+k�S�<�/���|�Z~r�T��/��vE����/� ���mR�^�={�4+d!����2�KK��&8Et՛B{�]F<���:<q2H%)_�H�g�njN�/�^��@���q�?�#�.A9m�/6�[�Cr_�XQi���Sf�F�Q�G��?�P�!(�Fo@pB�Ԉ�X��b�?/���N΢�R��6���s��d����B*;c_�z��F��3��](���0�j1{�۝�57��8�p~��1�jE#5�s�W�e`�K�g֪����HV���<�+��C�$bh܃5/��g�4�#�V����kP(ڂ�����rJ{