��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�����U�|4�}��3w���n��B�2�Y��Bر�An;|ܿM�MT�[�=��Kv^��L�`.���kS� z@����$7�.�'@y�>Cf�(t�-߂N�<jľZ�FLێ�"ּ���'�^{���L������C(
�?s�I�D/ܠf�Ӓ1Y251_�u��.���ʻ���-��6��Q�O��EX<D��7����ݞ���1��VӬ�'Q�Z��Us��'+�%~�Wd�e>��jw�k�&���W�Vj��J�cn�]�{��6��pAe碘��*��ɔ�oy��7|�Y7��}����>O���V�h�b2� ���,�a��i���G^�L���x���.�mriw�C���JȦ����ۻs颺�"m��v�bb��s���_�{�0XB7�ϧ�
�(|��Zٻ���9ޮЏ�%W�%����ؗ#�>X2˼�,h�P�m��K���=��< ��G@̇��Ю���B�}�!3��o�lZ�X!e\�+.���R�UG�	?I����ܯB�CI��� ?��8�pX�8�'ѿ�'�h��l��MŚ@6N�I�)F�����aDW~��C�37S�]sF���c�VXys�Gx3�x	R����h�qZ��T<�&[uM����6�4�_�rЈLAK��9L�8��c2Qw��Ņ8)h����$M�zrr�!`�R�^d���i6w�O.4���yz��)��k}8灩㴾�F�]&��V�z����LtpOB��;�=>�s�&�KQ�P�T��k�J���y�����O�p���9|3���9,`��EʝPb:����TMh�}"�K�=cܘָ�]����$�4*W��w:i|�d�3bȐf�S�2=��Ll��e��L�*����(���/E�Q�5)��I��-�վC��L�Y����r/]�J:�K�o:+�QA��p��1�+8uN�zs+�g�������K�^�g�R���M�!4z�U!��{�y���SǼlg���K�SZv�j��` H$���x~�z��G^�P�[cr�A��bHIn�o�l㚵.k�����5�3�S9��WP��^hn�X�W\Z��DsH�긘�L�[�#�A����}��D������2�@DkUfSky��u��β�=�e�0(�G�h�Q�-h4�_���ց<��U�W>��E~�~E��Pҗ�<)�h�Ty�}/� �xzK����9�ܐ�ӽ�5��l�JE[0~��,�oF珑�`ݰ�h�0I�Io�{c�����7�!1e�L}+
��"w�~��(��#ۘ��n�t��VY%t��c��I����D��hE��L4A�! |)��BuXF��_�%�����~`�A�)�<��ߵ�ƚ�4;n��[��L�ܵ�+�D�{�N7zcy��}z�9C��_@t���1Y��Yl�&�p����	vwd��b;�Q��XX��3�
��<���;���绬 |/p��T�cmK�zq���R�%D��>�P�"�TK�K]�e-�3hR�	ɽ�`a��a�?.���p�^vD�8��o�q��ӟx�8IKHO�>��3 ��J_�����h,���82`v"QTH7d��h:�Jx�s$���/6C$[��$�?�ݏ�{9��r<��EiV�V��Sgl�u��X��~֙5��WOQP�~W��cV�^�6��!��uUO��@�=�]ݮ{=c�fkF�f��c�a/?Z�YV��"H�FϘ �cMiS���tO���G��X���~�F�b��x�n�+�n$����&�K���*&Q� �RQ��������q)7 �d/?�|d��!{�Q�v�B�2��S1O����\j�S���Q��n�v�-�y^�����	�~2cc��r�?!zBcx�<y�DL8�$�7�ov}h:��BCm'���
���2w�c�{!�-������"TW��_aދY\�,�oVU�ŗ$AJ-�bBb
�����f;y�����_w���;�ْ��l�a� -Jz����h�x*�u�TV͕A��������?ďDH��q�m��R��8����Ӆd�����I�n�ᧃᕳ�+�\n����H�R����TF�#ٌ�f'�Y�FA+!�o3G�]�>|>�cz���+���m2�4�������dj�Ԩ���}U�z��}�VհT{zK/ϵ��$��7'Bg��Ȇp5���	G�>beh�W�}�@? �.IF+�!0�:~�8��@�p���-�loS_]�GB�,j��Lr���@N�nH��oK~�L�����o`zq$?n\h�l��a�9�-������LRs�S� 3��M��B~�E�{pܸ�E%5�|�c�>(�d]z����T.�m�;�nF�KC�`�H���Qnh(�,,�]��Z���2�=��ѵ��`�ʡ�C}C8F����;��.s�������De�(��uH$��:����C��+
}����..70�#���d��:�nk#��nLĮ}���#�Α����q$`��ޣ����n{YX�f���E?N�T��VL���sWt���F���a�ci*�m�y}"p;�L�ҩI��킠�&������(��N?�2~��ߨmu	O<H�$�M� �l�?f�L���9z}�U(�s�z��·_���;�{�,6�n*i�,]m��H=^�	CrP6�f[��NFkN�룤�ٔH��3!(A�ǀ���e��I=�T�f�72E7���W�Z�N���FY��S5B�*-�+u���R��e��m(���qmJN��H�9\�<+i�F8��z>�#�7Q!(����f���֭c��y���,%�mt�'f
F�{c{?Z��(Y�zE&���M��5(;s|8^�I�7Z$�;��d<5Qr��Id�y-	V��kȸ9_L	oB���ͥ½zv8k`7�T�h�_C0+,P�V�"�b�*�&�{+Q�8|p��=�raͶ�ծd8�;y!�v����z��s(-�7�q�>nh/��K��H��4?U�G��8��e/	�>�~���Og~|�kۭ�z$ņd�K��ZY������ q�;^1N
n���v~�&yA0��mr�6$�j=
x��L�t�T]��w�3k�n h;S�nhx��g��pr:U�r�>T=zl�?�yX���b3���h�����FA��Էe1-�{��gu�)p�����ǯ�v���ғ)�]� ��Zq\�7����a��C��֬Е�gl�Am�u}~q/��$��&f/@\_���ڵ�o�%&��2=�Ml{Mʕ����>��CN�k�L�U��0������m���U���B�1,js�/�OG�\�Nػ��� ����g����G����2��EΎ��G�bJI[ѫ�X=>�U���G�Q<%9!�&�\<.:^IG��'�N֯�N�b��s�Ci�O��[��d_�7�z�pם�Un�=�e�㚴���>{�ah��wC-�L�C�GP�a�Go�����mO3��7�

2�b�'���X����M�������w�uuI�Eayr}��#P` ��f�*%*��⌗�_�ؐQ�ol��b��S2 gkľ����x�O�?e1�����	�m.�aXl=i��{�����4//N�lB�RO����J2��"�e0�Yv���(�i��K�U6��k�������ho�ZO��+ '�+ӫ��>�,8s����*.����T��.&�{"��p��(�@=����?c,�o,���?�bǨ���Wq-v�勂��t��kei�K�+�bS���q"��P�5[6#N�W�@K%��7�vC���+i2d��3�G�i��_�|�Ap��/�TD����d pjq)���A�D�HO)Ϡ���.���z Anx"�7��[=�^��X���?���=�kp���x���P��݋�Ӄ�t��Q��zc�P�jǵd�����<���2ҹ�����a��@�
�4������Ow��z�
_���?��c|g��0��
�~���� �PJ�Z�����tBK��wUS�vs[�#/g��oK!��V��W��π��>�ڲ�ek�>N�=����Y��ЍA|�t�й�������w� ;�g�z�8`)6�u';UY�}G���|+�\���93v�	�B1����� ��9��g&���	���c.q��3��Km��uÉ#���u��0��c͕$l� ���� ^Ml��A%�x��U1�8��/>X��w�������w�=���Q�q�od*����� �j���0]�R�UC�~7^V�K��O6�q�B��2O�y��v��zb��&���OL�iՋKᮘ�Z�9J�7�ʅ2��d�y�k˗w�uޤ�s��W��E�)�G���U3C.��ʶ��E��K�e�Qyq8��	:�f�k5��4G'E$�#�d�M~�'m �z෨�0����YJ��X���.�,��[�a�?�g:�yS!����T���ِq�0��Y��o��Ji���$iy �P�4�~G�$�Gרߨ��"$�m0혻�p�{Z��M��|NhS�����mY��8{m��tLT��p&D&��rtx��=�s�!pV���J���'*����W��&�;��U�$��7S���tx&:i�ۡ���j�xͯo��������dbq+����Ԝ��q�ɥ�)f�]��~V�WC|4��3UɥL�;H(N����	b; �S��%֋�T�=��b�L�q�:}>����;B�V�n�#��-r�P��q�
�Ռ�'`�N��� ��x�MDcE�F����#�{Z�ǻ���)X�2��QJ^vA*6���ֽ�� ���w�'u.�IL'Xu{MW���z�eF� ��_v���?�\:��n°1���Q�ZI�{|!iÑ���
x�����2��=�C
�'�]�TD*&��Yo w4��8�!��|�4����/
U�i��u�39���`<Ы�R�&��2��SI��~%(	�v1�>�=�7a&�.�\F���Z��M1��[�n���ڛ��3�݆�Q�k6L�s��=x<3o�k�BZ]����v\��c���W�F����>�b⫥Jra-��-0W�-āk������M����%=h���W����[��h�A�3����$�`���>�sy*-���VP�����c��s,�Ĭ]�:����$>-�y�8HP�{x�ވ�W�	����I;�_)�������{ �䳳`����\��+�|��M�<��:�o��<F�<Ӭ�#~Б��\����\(iރ��%R��m��vё�&',$�v%�-V��Ig���⢶�OK�r�%�����_�0�s/a65��JU������h�Xc��}~(_v��9<���T���>P�ʔjq��[��`1L�q�ӻ�2F2�'�����3rL�ϭ�f�P�3^���a�>���7�R�����\��	i$2t2��^��S]�*�K�#�ߘyȚ��Xn@Z�s�C���X�����'ś7w�cuk�J��ѕ�~t�E�y1�K��~ȱ�@k�u�$$��#���Z%!�)�6-�+Cu������e]��� @�f��j�7�ج>QIH4�=��>yI������Y,G�.�j��|�e��d�g��ހ���9��N ��E��!��6/�~�x��ށ��;��>���,����N�5�j�;�m��;�x�j�������/�p��s�A�ob�C�}���І�[t�Тe�4/��*꣫D��p5�;�N��Өw���_=����@)�W��ּI�.G�]gCԻ��
H�����4�a�Y��>��~82 K��F�y��l�	��-�j�ug1��xA��2:�{t6�jXЕ��hQ���Ek���J"�ek�j��U��,g��(�^����69vfg�U�!	|����+�:AM��û)~�ZiÒ�\{
���à �<�s��Οb�(�Wf���2���u0�%%?���ʽ��2E���i�NO!]^�ė@��gk[ᆆ�f@��Ѓ��*X�-$<��z�L^�0礕�ju���F�O���6~7[�Q��%�"]�EN´2�rb`ʾ���XE)ی�Q>';��]���)=�ڶr��jmpge��9e[�;O�QD�f�&5]�T�<,�E'8�Sb�#����D]H���Qu���H�ٲ|wL�V�%e�O	Y2��e6�~ි���<2�VJ�BW��{�fZ4Oh�h�j�)DJ�T����QLNSȣ�3x6C��i��#k��m��ć�����LĮb�/SJ�!`��${��0s��$9� ��s~ьP����i}S.��1NB��׿.��+H��w�Y�L���sV��~ �������+峏8W���/W�#U�rM�~�O]k�rh����Ά��K��v�uQYz��y��4�-��!�v��d#�����(���TZE�pv0)t��U2�GS��u�7ui���3���T�>�i��@�(�x~�h�z��,�s�"�'����iL_Y�/��~_�*�rt1JV��� C�a�3	0�cǜ��Xl�������v��^�&��>�i�� �����\�l���
�"#@�q�Y˝�۵bW�6w��p�^�\��j jw�$�X�%�y�l���-�|Ri�3��!gMk��Y6Q��+�R� ,�����mגT�쨦��,����4�$[�Ȳz�{�*7ZV9�أ��,��1�4�S]� ���.�=c?~0�;w}'���+��\���E/���!������\i ��c�HB�-�Y�h��� �sb�@�C�q��Pu�(X5��N>�t�1��}���e�P��.��F�ۘ���1?Gx\�����|��,@4=�2�� Pe#^	Υ�~A�,������lM�V��S��}$F�+�z�Z���H�,����ح]�;5��;5_H� �]���"#o��ӟ^ʔ���|��I<������@���퀁%�-<�U>m;K�1kE;ɣ�됝����L��iqSjk<�Ff�����S�Z�c[�w^�جhl4�#�mu�&�F��x\�GK��@�gøPqU}ۻ��k��[Qz.���%UmV҆�w�f�����P��.��ڹ��+�s�?��'��Kگ86y�����e|ahC!����Uo,��Q�֨�/B�b����Q�4�8����g�=A�P�Ep�F\�+ qk6�4R�R�0��R/^C�@^�sw%�tb��=lU��/��jؾ��ѕN�v��| ��H*9g�R�]:��<�L��/��&P���aB���^fؗ%�L2P���W��>�^T1�'��mC:��� �#��¥����;���f�.�2ɫ�h̩Eƛ݉�'�E������Bh�C*�����#�79ٞ��0�0Ղ�y9�,&bɔc�G"$g鍧�|͸	�`b�����|*���M�c�.�R���n#V���0{�\�k��ྴ���g!`a$h�e5=�Z�T �>C����c�WІ��y���C�P6(!���ob�� �D��8rz���鍄ϻ��qXn9D�~�M3:���?�F�k��O�'�j��s`�����ى�ҵ~��ߔK1�v�c�}Kp�gú<��Ljɋ��|B��N�?�[1�W���ۆ�ye@c�ߖ�**{ɚT� �
谘gfH�rǭ`3)V9�$�d`�:X:-!�G ���T��u(�l�L^�5KQ5w�	t���x8��'r^~&q�tx<�����A�\P �����[&�r9.��AJ�R�}<6�$��l�٦8��(�s��a�϶������;-+��5�J��Q��+8a�>�V���y#G����1�F@�6ǰg~� �|�L��|���/Ӿ~3x4#�*@�C��W��0۾7�6�����8s��O��M���(��ܔ�8����p��������N8ο��g/�G7o��v��&D�� �}�8����8R�{��y��b�6E9/n�ĵ�W���Q����+aEF�?Eڛ�a�]��L���~ �����37þ�B���H���H��2e@� �0m��}k���_�:��6Ԕ�bzW�|L� ?&����$�L�Ң%?tAκ�m�2@޸��Y\�y�[���q�7�1��Q2�Al���~[�'����<A̐?����O�b)c�Ҍ��	Nk����o��r~�7�z�O	a�H��}����&uk��a��ɦ���w�K=�T�S�(m��4Jt\�K����q�'�<��=*��29ōe*�-uH���i	��nQ�Y���J �؝�J�#:�.�M�MȫE
��rP�q�(�-����aL�����@�e�G�b�b_�Z	��8`ƭ��)��2V�4�QN{/��:����Y<2��]n�k�8_d�ڊ4g�3�q<���k	��ا�Z\����Q����ǜté7R����e4���f'��D�4a���(NCWͿ·���<��=�Y�N���(u��p����d�c4r�G����{@@jT���)Ka����J������
�,]��4XN7*��n�e�|��Y���`�������U!�|���VOz�O|*��6-h��K��FH�i�5NT�K�����^ay��V$.��Љz$��2z��ω㲲+7��ב���ظ> @�Z���k�j��-�m��Z��12�X���B:����u��w���(*����V��Bw��DhN�w��;��x�p�b>�V?kb	7&�v�@�i���
8�F#�&�oz>���B>Pr��鬏�i�>o�'�6U�V�5 1\��`.���go$C�n�hX�6�����iͦ��蹐��)�����Pl��3�4��l�D#�J��;�4ČvH����@d�?^�*jԽ��a��*Nu[�;y��~rr�;eQ���I���7��imRC�������f��$��YwӑR�8��������	����Ώ�r�����nw+0��pE���|��/�|���Tt�g��z���P1,
��"��r�o���\X�H2!���gED*�����m���	�
և�X%��c��8'_X�`�s{ZH7\o5g�UW��?F[z4�ۅ�g����?ױs�0!�����L�h���Ɠ���8�~VX������|䚳��d�������2�E�;���	
���M����4�}���a�����&�E�!��v��ssw���L�D3�����܅li
��3A0R/	��p/�%u����h���q~�;{�ۀ�@��]:F�Q~"Č�A�.Ԙ��-r�^�,(�4���66�ꚖׇD�D9m�h��4Q�!509�,�3��V)~y���ePW�`���ͭ��X��G�ڒ@D��;^r����G�FmmU��]1S�|GqF~�[�dM�	����0M��u���E4�C��/�D����:�Od<� ���t�Z�)a�8�f7�7eeۦ�H��
�\�L���e:`�h#A���|�G �y:&A�G�}�ޥ(��=�ľ���	�/+�0[}�͍��:zx�=_@�^6�T�J���R�)o�����)�V�w	yή$���t����G?��t����=�M��q�^=�o��RW�;ඦ�M��a����E���CY�ֆ:s%�jJ5�fk�A*�ݢ��W7YY�������c��X�\���^��ˆ	Ǵ�Y֥\���(�r�9R��j�)H!/{��=�
Gi:�d�����xi��"2�#wÞl�0�T_&l��/&umVr
 �IUm��=A�C$���Sup�UW�z��3}ɻb���qM����-����~
���
�r�k�����$�zY3[z�O(�*A�F,�|XBǙJ9��1l���=�zH[W@�{C���J���Y@A�͊c,6�:cmJ�,�UmcWP��Ա�9� �{`�2�
s�	6���T6ʝ|��% �� �W#X��0�kX��rs����8/�^�'��U�m�+��r�_�ե���|��+��o�M����+>]�w��k�k��APS���p�e�����-��#�U2j����Z��RCr0���������n�~	������K�8��,��8�pfF�ǧ�U�ԉoL11��2j.w!jԌ�o�������,4�*��1�j��������Q��=�j+;��j��e��6-�H��.�������i�1�L�������F�É�eW�bz��Pԯ����8Q�m�m�E�a���@˄3P��g=�gB	�����jN��`����nڦ�v�Ƃō[!I7w'iID���!�>�X+��70���{���M0 :1Z�l9D�J�.�"e�3S?Mp%c-�+]�W�o��,\�F��i֌����Q�Og|�����PL������8 &�Kc�=#2Rm$*.coRc�X8�����:w�h���+Ti&�_o��	"����/dcc���C�T�:�ֻ�W˂'\L�����p�|4P͚�U=���,��v,�>u ����x�W����?E��_p�`�M0t�vf�jl%�A��uK��f�Zn�O����xԓ��L�a8��g�.6F�Wz��дgw�N�\60���,wA�l���+��/d<�������	��l!����#I����Ǟ=�/�|�(����lȣ�=9g	c�*l�?zЮ������_~�ZK�⇂|K}�U�Y��};s��	��]���^~�
>�1� %����RQF�ޯw�ε9�)hW��xe�p��9Y�%�+����[�ި���ۢ?ߤ^^���-����]��Yl��G�ـ�Ӿ���#.L���Bݸ���^J�;�+�l9�%�<H���u���U�JT�\~���g��s��<M� �TG�[��v�֎^!�d��x��[D��\2���p9\/kƯ�7���&D��rJK��-����D��8���ab��:՝�.ݹ-�X����_F�D���=d`f(���.�XI�}O�Jg#@��2��ԩ�׾Ǝ�5� ?����8FWn�15!=�����5�l��|�{
x�������A��"V���DT8�A��]yVB� ��L���ر��D6ʲ��Z��"X'oI��mZ���Qb���'���#ݕj��,\M�����1;U8_�}���4\U��Ðz�L� :�+px����W�P�+�i�>Nr�
Gb�`�E��[*9w_g�������(4��R$�u	%�l6�_I�犠I�rA�_V���}3�ɴ��I64s=Uɾ�+t�z¾Y\%\iMr]p^ϷFk��(���+~YG��+Z��*���{ȼ
���b_���F���f���0�� OF�޳ ���"���f���t\�b��/�Xn�.gP�\~�L���Vd��U�s��z<��KK[UC��Ǵ<PZ��'1��9��S�h3V��� I�����6"�]�K=;�[evr �1+��y8�7���L�ń��gyЌz<wĞi =Kzs��;�����{�H�Ǡi��	�5i5CEp@H�t�8��O�����gƵ�{��A��vD�����c:�w�^��ӉZ���U�{x�:$jܖ�9��p����?�8���&�e Y��3p��|�ȋp��Fywnb�K�s��!�m���F���E�1��VL�350��DێuۊڦLYs���r4���`D���
.�p/��7�͇�>�V�%>X��"���d�=6�pDE'+�mPi��s����@�4a?Sd1�A�uIfE��n����3�l�j�㑐x��~�5_���DV[]m,_���@����� �?�y{9�V�=?��m���w�]j$}J���>R�Ej��k8�B�Ŕ�Rk��H�^�l�N������e07P����K�qo�Y��F��Z�[.8�����*���$�/:
8CD��Z��-�1�6Ż~�����:1i�e��gox
\������H7)�#rg&s�R_O��j�S��6!�l��,�h��zB���w���Y�Dp�#�	��9�HV���������>҆g�Y���s�A�%�)I{?�OAZ���٭����	bIS�뚴�˰M�G�Ro<��r���"�������P���A ��Y)8�I)��HW�@�l(���/��f%����� p�þ�==!�7y�����7
uuUVݧ"����C���u��8�OdF"������C=n�h%�ֽ�a�?����q3Zgq�Wr������Q�`��/u��Ք����Ԇqb��`)��7T^��a$�H��Z��5%y�.{}���/AA9�eN���������$f�y�� ii��g�\GQ�!qL}�USXn����s$#��3]�0b�y�C���X���+E��q�C�
^����:'UUC�P�*�w�'���\��]�+��d�K�nV5����D��Z{��&�:z�!�3���a��tX���z���h���m���ҙk�N'QX�(��'J�[�V�����Els}��@T�Q�����k#�t)�:���rW6�K����-Ij�����ٝ0qX��i��R�g��A�s6���У��vW��f�g�K����u�Q�g<����u����g�z�C,Z_b����q��5]E��}mVi!�%��땖�_V�����9�`z �ޕ| έHe?�+M�%o6������!���5�z�溥���h����iJC�0�h^�d68�dN-|�V-���j�:�.Z�Ck�w���]�`�(�G�%�P�?��ԄA�1>T~(������
�R�=m_�؝9(�ƺ`��;$+MK'g���kdS(�X�e�ۢ�?^�E��Ǿ�o�H����u�ڞ�`נ���C���&pcd�L��!�YG����(@�v<���s����0�;�!���4F`͝v�/��}Z#�eޒI���Fͬ��Na�ǋ�d�cj�;i��~w����&��a��q���0*{�b.:��k�^j���i�-u�`��j"zN�v������ې~R���W�\��\���źO6|�_�δS����Yvޒ����E4"�h�4A�M�m�� o'J�h��J�״1�4���@%�^�Ûh��;�!�L�t���ڤ�J�ML���T�F���"o�N]�qc���9P��N[��Lg$:��ۑ���Ư��l�m�v�34�Ǐ��g�6c����ˊaw���(k�a!Du�4��t'=���dŊ�%��1��tiV��(���ى��|5 ���6��C��U+
�Z+��Q���o,ujҝ�
��x&4�j�Av������'�y3b)��y2��n a�J���
-�/�^�e�~G��m��Q�dj�o)h̥�=�?Y٢��*1�Z�R^�K/�C��h3��7L�W;v���Svw��9�\��N�~��IG/����(��رT^�����>�y��}k�����d�C��Y�Z(���������?P0O?�Br̼w���/u��q O�g����t��C�F
���� �q,�N����uVUM��n�i�[af��a������zaj"�)��su�K�.�˨���kD���6��k��z�%h��d�̠*�]��`j&a���|�ë5�'�T^��m��h�jz�!)Ւx�Ɵ�0��Lm�G�C��%@����һ�������1{�4]P+2`��a�.���\���up)�7g��p���L#�Ɵ�!�s\'�x���r���_c�b�.XY�PC��Ȗ�t����M�Gx�Wl���]'ޕ!�%��a-�QM������<���~���u���*�����ļ 7$�֯��pf�'�ށ�A���U�Y�2�lvA 1��=��;I�1�/��o D�a�Y��-O9�����Jz�d���Ҙb�^����1�0�5��� 7�f��D[q��y��u���}Q���d-�NRjz� �X��Pt��%)����������souV��1�Cz�X� ��Pa09���#{Pe4{˰ݶ.�T�G:РDm��p��t/9��i�-��µ�{�w����-+)9�"5��^m~�Y�bO��'7�@�1/�{
��ў��9!�?-C��`m㭻{�w������c�ꌒ�1��=�ZT��T:�:U��"ܭ�T�{L@�a�%�v}t>"7런zf��}�<M�K�o����7S�5�V��G��E;o;q�Z,F���Y#sm�����$ᵉL�g�#�-=ַ~��\H������[M��Uɸ�)ۻ����s� �o5{:
�=E���ڥE�i� 4p+Y�p�~�A!�ʺct�r[0�a�������x� �?p��N�|��p6���b��؉�k��!�������W�����	��\�uI�g~_�HY	�W�w��Vr�$*D!����6l�*
����L��,�[��u��{*alͽ���Ca���ϴ� �s��L�G��ɡ��&2p��w��wt�)��Q���IK���V��~�C1�G�L*R��	D����E���Qӽ Ũ �~�.����K>j�����+��
�� ,C'������#ȵ����qZ��@l�@P�̟�"�{L�t�v�D
�gB���tm�jH/[���n�z>��OJ��V��riD���A�k��
�Aa"�z��̪d
u������}sk�T���f���5�0��/������PTq�[�&��OFs��a�` ���%����i�UE��q�"ș�r�;�f�e�\���N�:���>��L��r"a+�57��
�f��W#���K���@��3t(��-҈���?Yp��5C� ������[\D �"����_〜��O��y[��*�:q�W�*;I<��K��pc���o�֘��Ԋ��lڴ�.��I��
���R/~�X"��E|	���;�o%���&dE��:�R `õ�D�(�>�r��e	�H��)��1�G�~�|��s �%�s����!Z�(G^<�z�I�(�:�5�~�>`ؠP(#�	�XV�/���XV��
;���s`C������wPH����>=�}��E�a�{'k�g�ڇ**�]�_��/.������=`��g!f������������P�\Ф�!�������*)H3{Jְu;�֦����Y[�.��	�|�[���&��Yc�X	�'懀���:���/|L��Md�(�7吙�{<�A{��xN�0�.98�g\���_��޵�	(3c������h	V_�� ˎj���"΄P�q�PIO8~�Fa�2��4$�ո!�5���a�&�j��q�@�^���C7��;�1���w�G��˒���F`̐�1+�����MM�#<��P�nd�f �Ώ��)��`[HJY����_���>�e�ķ��k�
�S��@���8�Q�Z�����6ֵ��aBh�zaq����������9y��Y̜�}2�7{�O��W���^x`"��0��s�gW�iqA�����pgȖT(TO:�C���_�I�|�nⱶ�6i��	oM�ɣ���&*[��7,����̘|�������8�"���3�<Ն���S��Z��e���C���״Z���t�<�U��p�(#k�u�nR����\�����&+-�,ҭ&b5wEH>ţ��>d�Ӝf)qg)#�	���q��J�5䉽��"�|�.:�����%?exT.`�2��یi�I$]�6@H�K���W���euΎ�(wW`*���,�Gߏ�d��LF޴�z�$�IyCa�tp�M�������@�1팿T]��V��ltQ�pk\C�0IQ�j�%B.�#/�^I[� h@��>1�މ���X����(��AH����m�+�z���+뒻M=Pxd�w
�������_c���s�>���-!��< ��H�s"6K>�J��{�A{~���~P����W{�p��}&���w���vb��s�ӗ�!YݞI���L4k_�+/�yq�>V�
��bY�4ɑ�n'���
1��N�&���<��4�A]*du�1�li�~�'D.��hG���E��y��AIQ��d�{�f����$�r�}'/�V0���p��x����AͧA9;����!����m�Ȗ84
�_�����*0���������˻�<C��m�`
A��Md����^�9�̕��C�A�@W�^Ǽ��U�2��$
NA�����ҿ�j�ofQ]�$��ȶ3��C#��n�oFn�E���#ES�1੹������!�Aw|Ϥ/��2�q|[U�TX��u̸��:�)�r���0�?�.���b�K����s,�^�⠆De:�Tܘ_�S����d9�����ZB
�o��ښ�0��"�-Bb��X��[�+��Z�4�Z���jz��'X5���/2D)J�6�5��`l0��A�B.r w�2H�u�i&���	>�Y�}߃ڄ���1��э�x�>9�w:���Vt }f�@ v_�������a ���,�IZ��q�^k$H��M���q�����TM�M�
]m�aΫ_Y�Y�N�Hr��.O���	T���98���k��_vDؽ24��蘎<��Wg`U�]Ӂ����1(��yS�h�B��^-��g�>6�Ͻ��$Lw�2^����w�ǖy�K���r<{{h��
��#�W�,pA�c�(�Q/��ϵ��?�S�G���f�G5�z�i��|b.�\��C��M�gެB�h@�^s�8����
������m&@�԰hMUV:�L\�i -a��y�.^�A��$P��W��<�S��c{��xw%B( �	s7ڴ��8!O�2��B7;�eFL�JA�5�W��S�Px'���Q;��x�D4�� d�=f;�nr|�֬N���SU��*��hC��C�>K�5��#��ts�<����!��_��#	��e�����C�С9Y�?�*>�p
�lIW�E4�L�
4ߏ K	V߿��e���;���'7)�������w�_}����aD7���P�Ě�~���(_s�N;�{F�1����Ig�)��W<�&���p1i�'3�:?�|�XAlx�%G+'��x���l���������j'�,Y�-�2?�B�I7� f	4��'�C�AV�lr�c��2KXI����+�o�;z>j+�L�T�H�2��擻TȒ���Ka#���g�0�/�k�3rI�8B�=�G^`���,q���R���ƚ�8N ��06A�.X�<���5���ӥ�v�XQ�f�v�M�M&��aƱ��o\�+]0Ԕ��f��i������F�����y�Rk�����P���ȧC,gV�b�c �r�*5���$f��W��"i{Zo���E-��O�[;C:�u���A����u�;�&C\�Q��P�%*^���`xC�d��e
��YH���fWڸ��G�]�|�CE3����+��yH���;d�C�ٟK�ƨ��!�5�5�[���}������n���׬�U���󽅾=r�eH�A�hj��fct���\P����EL�q�f�7b��^�g�$tk��y}�xL����.w-X�^��T1��Ň��įe���kڎ4+�Q�� � @\|S��x|����k׈���.�b�Nh�qI�@x������� �M3�;~p6�a�B{�n�����D]�/����N��X�^�K9N��Ö��4��w`��p?�u�z��0�Np ��'��Z�(��b�"�{O`^��ߌ�w��k������2����ĽCJ�2I�;��������5�O;)�r���a�{{�w|����󔠤�/O�=�}��Bm�xt�L�w(�T�E4� ���><��^I"AT��;��MŠ��3>�������WԄ~�b��}�q�I�㶊��[5�-��b�ħ���1IO�5z,�>*g�(s�[���rt�)-J*!�2q�A�Z����~�,��w�2�c2����y����q]Q�}�~2��RH76��=�o���2�t�h���C�E<�� �	ѝ���es��nHU�X���N��vMA�Hˏ�s!�N�|k�Ir�zrD,��O�䒂+.��</7�A�=��B�k	D�v��H�6m�8܏�y[�\�{l
FC�b���I�m%mZ�@��x����gS�/R*�p +���c�nA&mFc�S�&�\��T��:��B�O�\W��*��ZO�OC
iP�o�X���kJ�/={��Ǐ���o|J����WW��k��7���w�/���&/��%S��hP����V���ˆ*
�������և��AB)�0������F�PA�n��xQ���y�=�@�1%�����r�ˣ����m)�6�ұ��<�R���$� �Б$���R�ɔ����p}�!�D~�^��ϲ�%T�
 8���c���+2�"�@-9��mX{q�#aw�.L�Qy��spH�I�y-�,�R�;�c`0?ؓ
]&��W�Yk�U���N^ z�<ǿӎ*�]�`.������Ё�雑��0��;o ��I��,�Rf�!��˕ć��׋T����������b�8����+�a'e
�$�B��\R��\8o*$9Wm
�뇞�F���c���7:(�K#�dv)9���&W4��K��Ksv�t1����^���5��8�����_�s>rqhUf(��9�}ʽ�$m��8+���
�5���
7vY���U�2�b���t��X}g�@�i��U�Nk��{(���[k	��N}*M�&0�$�Wv���nf8g�~�W��3��C$+�/ڃ�b�CHR���X�Wn"����%44{/�?���7�&�B�9x�����2�U�P
:VUA�9��i�ݫS	>�%�QP���Njo�|��A}��=	H;?����ar\ �W{��� ��I>�ڎ���>�%r}_� a�O�U0��	J�B��,��q(ı[�.x8$c����y"�_��-�܋g���	f���u�ac�D&lVF�\��8կ/Y�ZN��*���Z��� �Ş{���u���vB��>�&��G+�6!�1�"��o��+���(�g0i�>�R��q�6��=P��;7�����ߏS�f.n��|-���P�w�0����T����-C+w6%h�2�'�ء/<7,A�I�yjzQ�����=�L54?*$�b�;�`��Y蠡Y�q8��|����cJ	\�Ԟ�T�)O�W/G,����E[�Z�qqq�/YM'o�f&O�?�:3��@�፹�'��P��AG�L_H���~.ҕq�"��}..Y��=�����?�[�\6n�V�����޼�6��\3v����~	�,:���kOk�P���@孩9�6��ȝEe`8�旴 �Y�Ҫ(TTa���W�#vr R�����yw�Z���75��`MsUJ�d/m�Q�B)VR��R�nҦ�@��p��N�U��gSL���?4L�	������=�Wة�,ꄗ
(�o�*=�����5�P��H�+PM)|�.��h 0X� ������-����h�>=�z��cgL�@���{g���ڇ�鳯��ۧ(IEV]�Cp��������no�d��m4�\(%�	.i�ݼ|0jJ��]�?d�]�
"�19���N�޻=)��V�h����B�与�:�Y.қ�}��I@�Q�1��Un����qN
�Q������=!���F�g��tfx��Cxe7�C�����W���n�2��<�=��x�ty�h}!s�Ʒ!�S�箁�|�T��@���~����p�2b��6��6��!������(���ɦ���nQ��m�Ӻ�:"�){?��rR�Zd\��2*�]��dwNr��^�\A�B"�Y$j���$]@zR��,���c�P��|�tK�!��N�&s��c��Bvm$�뷋.��� t9-#�^��[��*{ޯ�T���3q��\��#O�m� @.fxTf�����N*����.��^}m�\��1�޼�VȥY9���2����ȥ������"�o1%�O����Ʌ_��|f��
g�ˑ��_�	���ۗMvn������
��|��S��{"=5
�5�5P ���9fB�xMLkQ@����T�Dc$ף��?�}���	�r���P!X�$&�k����=bx(Ys�[�\B� ��[$�K��w�����/��/�OJL��IyH���� ������<	ϐ���%��T��O��A�d�G$R�ax��q��Ҥ���Z��6���BWzg(HK¡Wc������sIuZL�\�&�%�#>x�~���MrTWiċ�|c񽹑Dm���D�Y4�
����k��|�ՂO��X<��-A���=uGx��'MX6i)�I$Ow����;�P��h
� ��ݘwY	�E�j�o����x�EvE|�%�����_�sJ��+���������*���Y&�N=�m'�7+jt��K��T�l�x;����(<�_���w�ym��n�����"_�uՍ���cL"���C��D��q]l ���� �+9< 9;����r\N��/�9��MBE�g%�j�fs�
����΋��M(A⻒��J�� �v3��!��|��Q�j�I�U�b�-����(�>n:1zE�GO��T�O|�p=s$�b�#�WI���kU�aTXjT��i��G�r)�)+Wvv�"����f�%�fYbS���s4u�K/yTL�o���lM���H��X/�P��C�F+t����DY�6G	�(!��Yz;%�Z�?�D�nt��^��ʇ�R?��/&8#̷wF��!�%�r#06zW�������~���VD57V�jOݑ�j0�8`,&���)�������es���r�179sܠ�X��&;�H����E}I��ꙁYۅ�m􇁗����M(�ℏb�.����s8ڤ�g����$���~%�� [��q�Q�o���O��J�;�v����j�S����#�b�a�^-��\\��P��r�ٚd����{Y=N$���z�L1Y��8c��6�4��I�z��'������+a�`��ÅU�X-*@��\oS��"��'u�v��$�I�.�*��X�u"F �Hi���E}eP4GK�� .�������8R�NO5�3-����.�Q5r�l%]��2��p�y� n�0�B���, �r������:�sf�.�?���s�pđ�WyAm���;��Ė2U� >�|�7�B?�[e�䟫!�<�
u��bA����8@�Β�l�D��dEb8E�I� ����_���N ��̏8Q�R {S��O�1~�6�䬓R����#2O�Z̤��-���&YbeF�rA[��I��%����8��5�6^T��W3\} �:m�00'3�4pߘXkn�T�~E=>'��]a���%6���wO�C���p�m����47}�����(�8-��j�T��Z��/͟ �7j��e,D��~���b�[|�E��6E�"WƯ�
��"��1 4ɾ(YL�ȹ���2M�@�� ڲF詜35�1)�g#(���9�ӵ2�-E�{�Nƿx�Qz�4K����v?�[�އ��F�t��U��l(��o�H�=.-v�,B�*�>c��#��=�"��y��~d���Q�����_��ȡ��j�����a����q�ɷ�_��7�&�t͌ZG�D�j����#���o�ϗ���@��K��;re��.�]R�K:wm��V��X1��lK��3|���z�h�@����m˪Á~�<�|�-Ht�d`*��b��ǯ#¾�b?T*P�G\g�\'�.p��&3���7�~Π��I�����Gw�GOՂ-I4R�gO�V��
{�z/d ���۔x� �s�kq�T���S,I�r��5Z��P��
l�A�K�8C�Y�7�N�wS�t��{O�׷��DF22�Vdբ�	#����+���9�:*��d�&�=�f�����$�$���&��ƣ�����,�~ 	 q���$�����>X�6_l��b2}�����GVHJb�`Kd~yiW���!� �Eҿ�0���w�����{!�<+��5"���5?У<�H�yV%E:H���j�3%S����_#�x�����4]�+�%{(C���+7r�@��x#�G����Nd�0uG�d�ЮCs��\N�䰻(��p�dV/��Ami�eʑ�<���
���&��8��vM�����i�L��7�F��-��{�/9s%b���TpZ�c=�@)U���K��W�9*�in��1Z�J�܊�h����� ��۶É�<�k���/G�~��'Kn���e���"�\!��=|���"�D�3J�o��f��Y-�m�,w�\��X�N?�s4fZG�~�9��ZYm�nC��:R�ڧ3� yڮm���wF:�h�|�1�[3`y��b� ��#�9^,g�۱�·�d�ib�G9n)hD��΅��Y@tb~-�&��%�p"��ك}���Q+BY���v��\��n�.�� 8L�by5�n\��lf�}ž�}����P%����Rh����%[5�v���"I9Uh[���U�VJ���-mxPQUAᅮ�eE��p��u���	8�D�min��D��*"���2�}���i��[���z?�'s>�Az��2�f������ "�dͮs�cUF3H�>^�i�u�CY*�x�tCvo^ �wb^�`X�_zr����d�l-�9c�f�3�v�id[��9<�r&L<k�o!v�e�7*���"B+�g���]\ܕ���7I�_�o>���3hV]�a���d�kltg�"�LJ��@ՁB7-U��.[^�7�J�h���Gc"�'���L%@����w�"@�2�+� �B���A$��fl��d3�ޖ���ea_��Fm*�ƨ~�{[�&�B��>�.f������136[Me�~����Ɂ����0>��*ķxpD�/�w�Pɴ��d��?>6$�'^F2�+S�?��T��q�FCnu����d��N�~QDR�	�zrxH*��k��Zs�����i�"D�&���.^�J�� 0����۰hتT.�ׇ�G𮲛@U�hZLu�Żu��nf�%5W����i��n<Q`�a<�Ԭ�~�MPl��!��K.*;6���'�^i/+�jE)ќ�4$"�vF6�_������S�p����w��WW�݆���R�q�%i�|�f�4�	�6��������|0��0/�;�U�8��=W����\3�I�:>偵�JP��q�2� B�
[R!��Χz?��	���.p�kQH�3_�7��a̳��e����~��<�[v�B���:�`7P�uw�±��[��R)��0��'����YL�\�~	Z�.�M�I?��B��]��
�w"�6���� ���M���&yG�+G�$)���k�dN4�J2IۄopUb1N��>�+�T�W�d��v�*��_;�4�X�������>O]4�e1'S'k�Q&�T���������Q���{�2�f'�t��\��W��ZV�@ԢMEn6�Ѩ8�����W7���!~�0��/2̤mH�vCe��˔ԛ������߀0츙:��~F礼��e�<�ȉ.<xL��� A#�=쥞�����eX2,���7�9G��P�Q���=���'-ZO������	ʵ��H��QIm�+7���w�q��1���ڄ��Sx4�J�4��Q��a�
<k�C\a*){=�F�s�C�`u m�*}k~���q���]\"�m�)���� �+@kW�^�$�+��!�Uݎ"*��&�"������]����d��xr��&�oc�JjF��wb�K��ۉ��oD�!�i�J�[.�jً8?�+���֨�%W��*�5F\r��j�VdE��p`��6�+{���KgXY}�A.�]!;~r��	���ht3�+�[�� ��!l(_O���	}KՆ�o���|�*�� ��>5�D�K�f�j����̈Ky���\�%s���Qe��,��*�C��c�?|���I�cJ饩����	�q9��;��V�����ɌL�����E\Aƪ�Ѽ��(�{>.Bs� C��BV�j%|�U�<?(�7�^���%���f�E�ho&7L���z���s �0u;=��&%�k5PQ"_�G�<����9L0j��v�臛�����kd���5��{P��a�����-�kĪ���6���Q�k��^@�W#Թ.�fݬ�[;�#'T���*��*�_bVC|p]fIп�F�i�a��dG1����dw���&dG̛S\`�y�CV|D!FOMQ��ٔMGǿ�9b��C�'6�����Y�4������+��	���Q���Qx���fN�6���F_␳�{�s~��ͮhG���	��;�5`jZwkIw�R�s���k'�ǳ5@���ҵ�d��Ä�wΖ�����Q�gN�y�D���TKU�i�^��|�>�죭˱PI�SWk:+@���#*	���~q[,�x��A�fVŚvJ���t��'���[xŰ�+�{���9R�Ƽ>;�UY`�((�J�Y�`dI�=čQ%����a�C�(׹��N{Lâ`>`C��"���8i��1����{FNBH�b��C�8f���"���!5
�e���֞WˇY:1� B>n��Q}E�U�H:�̱yJ$-n��}���|���t��
�"�m����ɖ�����2�s"���F��%���V�g��>J�ʫ�ل��9��i�jS�-X�O���K������5[$�Ra��㙭��!�:l��c/o�ǂx��`PF�37�~�+p\O�!��[;�8��w"/��7(r��� ��7�����/]旞�$��U����L������AǷ�I���W��N%�8�M=^�2lT�s:�<顫$s�ܡ3��잂�5�J?�/Km~�E"!F1v!MU��sؤ3�� � �dcR#�|�A`l٦�& ��'W�68	"�]hҽCg��B�%�{���!�;��8� ��bYFhJ�� ʡ��+���e%��/����W�Q���<7H+�� �-�	Qgߨ�zvο�ȟ3��1��YFI�[���(U�� ���֜Hs�W��{��?�;��|z���3�V��|�5h��mnq�J1�8�@tVJ������*9�N#"��|��*=,M��g�B��@��)�ퟎiH��*�%`�V�ǡ޼��	����e��Rfq笜am0�%������I�j�r��P ���	�m5�@3�='����v��D����k�%�%���LI�~Ơ��+�)2�w��ү��+N9��9N�����QN�G�g�۟MW�yNm��g#	T	ҹ�[V�$G�7��1?dr�&�ı�QaV2{ӯ�W�T�͐y5)��ԣ����*�B����.�ܗոK�4h?��.wC�>� �%�S
>]/��.�g��M>L�[�±�~��7�8Iwl65S0�Z`���������$���[��]W���9#��Y���y���[`���If]��N����!3���[Rj΃���:$�'3����?���|���ܽ���[���S÷��ϊ������&M��d[6\�Q
F���X����!��E�ʮ�!Ļ�9@��Zl.�/���`�R�;�z��4`�J����N��m�"q�gG���$�d����+������"����O'�P�B��o��'-����� r����d��Z]�9m�5�T*i�b�k:�������hٯ��[�&!�4�Z��@�AY�I�I��U�/�[�'K���ybW�8�p������k����a��B���Z���vx�vn�a\rң��b5:̽cg�<�|T%$wG<����yCN�x�8UN(0"��GpW-��s�zP�����Q8�iAT̮1P]�:�)3kt"`L��bfm�z�=�X��p@�y)�º�E��������yP�=ষT��p!̥�g�҄��ٹA��c����c V�;Uၮ3�E"�[���I���뜐�-��(�ճ��&=���Ѷ���s�<���e{Ea���o��U�1O���J�%��g/�t��Y̈�4�f�����_p���}3eWڼW�U_��^_f�ϣ��1:]�~N퍽zo���D����1�Е�w���<�
�(U��PQ[��р�|�G��<_�.��{pXk_���S��n��O\�W�&�h������4���
t�-�����7���R�'0l�AQ���N��T��R�z(�5�J���}�{��Gi�pRpبB�g�_�E�4\ �/�E6_	����b�$�sf˒ť�Lqs+�Ɋ���Z�w����	�;��p�q�k~���,Lkƃ����g	�G������o���mf�|��d��*Y���\�Y<ȋ,S�w�Y�7v\2��Ϻa$A(m���ǡt>`]Ө�R�⹲���z��/,���Y	J��A��ԗ���H�v�$]�~j�����[jx����G��u<�a^R��h ��)��|BKY8���\rD�H�Z�l�W�=>3�H5Dؕ�n^��US+#^U��/ۛ.p8>���н�C8@���
��)���M؀ϡ��ZC���#�y:��i/ ����Q�0�� zpz��9^�̶d9b	��"&��,�(� ���|�x94���4�#�q���]J�۽j���!҆�O�,�����{�_��'��'�Q�F&��Q7b�;�ұ�z�y�`jۧ�&W.����V�G�s=����BuD��e|I�z��}t�x#6�b��p��%k�p����m�D?j�+7�ڹP�P�p����g3��<�O�Q_�ro�_��s���;��C����m��j�g UF����*��rFn�lZ@�T�|��<��U>?�u�p��%U��|�bV?? �p�*�*u�_��4�v b*�"]��`�+�@8班��S��� q�!��_=�y��Y��s��)�F�¹{��nj^�����؎��Lbl(|���3��#v�`X5�"���?�v�:A'��}C��)u����K�_��8�+ֹ:���������cm�S8+����Y�f���R��Zca=8T.^�>G7�J���ۚ7�����h׾.m�7��8䤩�W��p]�y�2��6u;�R�e�8d�&ݽ�_��0y���y�[d	�Ə.��[�Rג�����W��=9J��³�~s��䘞d�x�I�a���$Y^-m�2���>��z�`U��= ��~.x��w��pV�0�#t�󅷣��%��jܽ��9s����6 �!Ă�1,f�ǩ�-+�Y9�8�j�w\��h��Ԣ��?�{�z�CJxJM�5����4B��!�3�Vy���^٩�p`(&�ӆ���'=-3���tN%k��2���R!��#��ε0����M�#|��#$���7|�=�� �?�SS��X���w���G��	�cl%�/�� uJ_5hٴf�r(�9zQ�vpiĤ}�dw��ʫ>9�N%/���.�, n 
TU�)zuܼ��/X+�
a�k	��=\3Cu�׫��4����GzU�;�
*=����P�֘�2����!D�uj[�w������g|�'�RK��m�>p��7� ��pPadݲ�{�����pZ��$�܋}çk�.4��Ұ�s���6Y�I��/�{i)��|{44��z�޲�!x>fhOt7�r{�\����L��G�,6��� ˌ��Ǫ�8������+�d\+�|��sư �/R�X8s��m8��N*0|�I��3��)��=�~�p�0X3r�6�mſP���b�K�-Zz���\���95�Y�j �<���K�Z��C��L���"g�B�Xܰ���S�0}�n�4Y�Sjv�iU���������<"W��m��c�l���y�f�]����;���r^��W3_���A���Aɫ2�z�6M�0��r�Ow����)l��`��mcL"BDy7E\�Zfq���.��?~���AP!�T���/�$�E\�B�1>c5�͹X
ŋY$��@b�jK+�6�@�L�|�|���}������I	���� :�db������7���Y$TO��t��|�W����~��uJ	�m�3�|n<IS'��P5t�:��Rv�F�w�H�U���E���hi�yI��׈�`.�hp�ivxۓΔ��9��Y�h�����KĕEG�&��N1����K�rS�H���u���C�w(����u������\.�T"e�`���5��ڋl���lob��Z����Lc��i䱪H��1�U�=y��nL�h�@JpkP�
#ʅI��77$HYy(��BO��@�t��3���ȡ��S1o4E�W�^���<�Yd����o*|֖�F+
���,h� �yJ�g#�$'��(Df �<����B���>|^y������֊��Z�i1��D
�^��F����Y��1X��.�j���|\������Ľ>��X�P*��&�y�[��$WU�G��;a[����� 2�n����Ω�J�?;	��&�?��"��p��&e)K
R�9ۦe��G��,ڌ�ֺ=Ei���	����%h���ճ!��@O�엲=�=O�-`��V�6���K���K1Z�e���p��>�63�A���K�A��?\��� rs��V'RTG�5)l����b�!���X�6����0�-묜���H_d�y��t���{��gzVy1	�iV��sq"�$.�܈-��e=�)�G�χCƓv�nI��(�j���x��)�/zS���U�X�\l�<����߂��!0l��<�
�Z�(����,���m}��^}y������ ��Sl$�p�;�Iο6���3_Oe)`�.��ӿ�]�G��JOG�N�u���q�}�.�=;V�N���Ռ��Դ��g�cS���0��v�J��M��e�J#hU%�f+����T�wBbU���� '�K�!�FM��0�d6t�zziJ�nS�%gZ�%�� )ZR
HX�a��v�^*�f� F{����>r������S_UW��1��KIu5�$u�����r�����Н���� ���PV:N?Μq�Se���0��S��	��q́g�ƪ����V)#E����Y_|I�nIC����
đ�}ϋ�+2fϡO� y�*��r�͕c���rd��9��-�mߵ=Zr{��w�#_ �����6a*����ե��-�rc�4D�('녻	.m��>i_��iP�l~
�����qY�P?߽9E��Mu]X�ʮe������H,�YcGnl�gȏc�@"3Y{E$�����ϻ���|��V ��B���z�&(����������G� cs�߭�0�kW��c����$�*��w鬅n���QW���~�Ox"x��1ɉ��7.�*��B���PjU%%�!.��|(���1�H5J�\�����$޶?�b�2B��.V~���-�w��1��A��������j�%�͢3�b�\W���T�+�+�N�yw�k����� �!H�ň7�W�5�xzS2�.� ٰ�1��
(���ߚ�$��O,�Z˒����M5�ތ��"8�+��tJ��<�Ѷ��rMk�	��n���ѷ�/R44�ʾH�G7�q �e���%�h���5��� D�����c�|�͝������	��f��3���U�v���W2&&[���}O�ͭ<]ޞ1g����,��݌ 8��?����)3��z�*?��q%���#���S| ��s�*��`�(��7�1���qo�ቹ	�(Ώ���Z����5�C%,�D&��Rc��l�/�j m f��Z��`�-Mŵa�T��`�E̤b �a�-}��f^�==�3��×��Vi:msf��|u�K�w�,y�*M�2�zjĮ0���3�\큼����ϖϮ~��r�;X2���i����mQ0Q{�kZʣ�d�'e��Buğ�#�m6�ۆ����Xb�������*����� �i*�F~&�ئ?o�S!����>x/�&�}��vNO���l:�Bj7�{��SD����V��a���e'O�@���V��=�%���5�A�e�	�g��q�k���DeJo��0�E�x7s��i��0L]9�j-Raav�V�B����g��Ա�DDCT���._�qOB ��1�Z��:K��.�e�ax�O� 1�/g�
Ч�޺2�B���'�����Hʆ]�����a�i�DR)]��3�Nm���\�4;��xr�{��D�����|�e�3��r`��x��
C$B�Y�}_�D�3��u��N�қ���[���u���'�҅]8;�
|����t��f6��5U�J������oT�u1�F_n������A��	lu
��K�K����^��y�A��I�"6b�y=��ιA�e�����\~����H�؉�Wc�>�Au9	�-d�de��y���������򯲸G�"��m!���]ی��8�p��WC��
=�� �Gzi/3�"���$ȝ1fn'��эF/V�%�׎����'\i�����Q�8����d�75�n�m�E��*��7�H�q�/�38�/�;V�7�鼜�j��ʑOyxy�J�ZXBk۠�nņb�?WA|���{�|'����`���n��O��I	�%O�K�{j݉5��OF��3jTص~㓡@/�R��0���r=T�Օ|ָ8�	,�Ku1Ҡ��5�؍�^���e����x��~ ����y���R���@�J�:�#�a�x�>�]q0ص5��9��U���zߞ�q��% _*R��C�
 �ZT(&�N����B��v�I^Z�m���ĬD�&�W��,�Ѭ-�-E�� fh�� κ�۴�5z(G�_v�N���B49:2�l�T�$V���%�<����¯�lצ�%g�B�:�A���g~1�\t�*F*ݝ/x���(J���AOEΫK�|�]TLRn���m�Є��d�s8���ǣ�N���!�F�rxFV1��4��3BW�|���
�q4�,���ޟ�y[/|��dM���k�o��2,1�O�� N���P��ȝ7��	��e�zq����p�S��L'!��M�UA`I.1G��֗@���1�hA�c�h�?i��͊&|��\"
R���mT����s��\Gӧ�m�?�{�3����N���d�}kɫޟ�3���Ⱥ�~$��#�Fy��X�>�D�C�V�#��/�4�,ǖ��ʚ�`E��K���@�"��|Gq4�Z�#oe,��4"%��/������ n��v3OΦ�0�y3���aI�O���"���q��C�����>?ct�짺*p���Q2��
�a﫼�1Hy:K��ˏ,��`���q���e>���l��_Jl|W�k����Y�����2n���enY��}��K��Sx�e���t���g˵���}Jj��;=�Gɇ�f��$,�Fv��N�7GWjŅ�yKN�
�hw}t��G�[���=|Y3��=��4�����L��Q Q��r���RKb�N1*�Y^{�riH�#*��|�����/�e����,cHw�xd)v� �N�鴎�5�a�aE��W�˿ĕA7���C���<;���\3�yĝ�l Z:e9���&���+����>�{��������s�a�/MS'�1��j�����i�B�k�j���t�~�s�oӍl+}����+����t_a|�Ƕ�2o�0 g���&muuFo,M���6�֒ps"o���Cpi��.v����<;����ϡePv� ��u�Es�T�R]?z�O�$�X��'�*���������w~�ώk%y1<�?�`M��XZ"N/�	<8!����<o�E8^��"���W%l[�
�P^̓H�.���á�`-������E���?9e���߳�C���:�ύ��Yd���"d^�h*��g�ې�['-�\<��N���$��G��W�ú�ol8�ϧpHsu����(	��$��LẊ�҄����=z+�8��/$��ɍޝ�W}�����"� ���n9�yP&�i��� �m��q�>�E������"!
�!ܒA�#x}�����q��Z]6�k���MlEc�U��Y����lY�j�#i9'�Hd5�ۥ���J
��ʟ��
�ѲY�� fǴ5�z��-��li�cG�{v��	(�O9�m��(�,;|٠�P�� >n��<�����_{��'�R�`u~��:�U�5��L�p�W���6l�+u����_#�����=��&�3�s�������5b٠�E�-��8K��:I��g�ٶ��mT�*����E���d��F��;2]�� �Bp�խ����k#ډ۴)M����^V���X9ךϳ'Vq�
ʉEhT��!��Xi�'B3�ޗODG�t߱�K�Qj�t3Dne��W�0Z��ֶ z�nU`����>�}B��xrO��ĩ6���0�<8��5�z+��h�U=9#�C�+ܽ��4&�����5���j9��̦-"�M�H2�E[��Ʒ��/�� X%?��,y�U:�E��`��b�xW�艞��z���o�̈� �K�d����!]�}��Uz k�?8�~<�%2�
uo�bЫ�Q$X¸��dYe��K!v�h�fH��	�h06���R��r����Yo艵�o����h	l�����z�К1H'ߣ�
��	6�}�?�	�{P�H>���k�6�`Leӻ�+T ̷�S*8��������Y��>9��u=����@���>"�a0��ce��I���t�9�qk�<�"a�{[����H�MZ�[��p�Z�:Q{<��p#tA�Ad۱ ڣ�_B� (�Ymec��W��mE�[B9?U/��ӗ��BKLA+��d�4r���jj�� �b�0�v�5^��������%�l��Aku �p�w[G�9B믉WE�;;����䒧����'��/%��I��-���w@�+�n�c��n�����0�j2���!�a��]K�waIbMjGE��Bm�~N'GP��A��J�$�K�~6[�2���.(%���0�Z*��#���5�^��X&Eb\��X w�G��U��O/ƿK��r� �B�� pl)�|���뒅N.�-�a����B���4�O�~r�K���	ݬQ+���a�ƒ���<툝�0K#!�R�F�m�x�J@n�r�G�pdB3�q	���?�,w��f�@�0�|6u���e�D�K)!2��dbN�����kB���"e6���z���o��������rY��"�����p�q�3�G�}�� X1��ֹ~j{�&��"���}�zX�_K��)��q�<3l�~�������$�����4���on��-�������ѵ�βp�b(�6 ��&fgKw �ŜHJ�<���<tA��|p��+U)����+�j��Yi�и�r�ةީ<�bxA�[��p�f�����l�)up��T�eJYC�C�f[��z�E �⩓� �
z��:�w�|���q�ܰ.R"��^�$(��&�%$ΗT�Y�͍^f�}���� ��3��5R}�Fn���#ue��^_���|�����N���ԑk�*�����r7�T"��&/rn	�:�_o���,�����/yKw
��,����4z4�A�����@��]�Ɯj�&��R	.ƥ߂����`G]K��F����H-gG��D����������~xiq>��.��>��+{F�G8��C�TMS�F����N�Df��HCyi,@��"�h����ۦ���ص_�@,��\�ڦe_[�N�:5��Yn�BŜXc5b�8�Q�T�b���3l��m�FVȰ�K�w$�?P\?��z`��HD��Rzd��d�q%lM�4�k<x�Ϭ#�p�m�[���÷7�N�D�>�l�!�	��Z���h`6��QB�����E0����=��d@�Z���>�VoG�z�_1��� �N~�N��e>,���M	`M��!��Q�S(�h\|������#h����5;�ل~�ox��Z��x���۩�N�ˈޡ(@=E8��+:��y��Ғ�W �Y(v�|:��bQ�R��1���k����4���ep�a	dq:w	�KFhI_���/_R��=�~�z��J��6�}�T냾�+�	��~�7|��RAI�_�Ɋ�z��dX���1t����2	<X»�Q$S/�QaN�_����-Z
Pb�\��R��|*ǡ�"���=�Ϻ����4u�����1�}m�^U���#]k}�$'��:}5K���S�)u4���x�C�W.���79aK$�0N������J|5��Y�j�8$_�E�$`H�}�$���S�-0�C=r�K�m�~)`a�H�Yp�P2X*��윖
�*��wפE�o� 4>���-uo�Գ΍w�E�W�����m�� q���_4��=�уw���G+�Bq��Y�oK�]`��0t�T�?.K��-:Kmzv>�*��+�X�ƺ�$$�}hp?���~֩vAp��'�3v�ܔs�D:�?�O�ר�)��m>�ǁ�ku�����W�~��\v�:�`u�ңs�N���`̑�}�[V�JƘ�M�$����	ᛦ�'}"^	r�*��TS��q���
\|p%�Dj3S�lrxY������z3{�8�*q�jⱨ[Z��Cɢzw(:��)߾t5. �l|Ȍ��(>C��]|@u����X*�`�zK�y��d>e6��mn�>�S1yf}�|�*����R-�Fè.�x�9Q��9��T����8��f�n��Mxb�e��WbÙdf(2�qU[��a��)o�"{���֟��s�mkV [� ����}�$U���KA��%��X��𖈓!�J��H����%̟��6/	woX=� Vv��Z%0z���-��S��6[�ҕ���F�<��ƥ�Aq��N��T �%	iy��e��/�2}�S�}7�d�0��,b��������8�=PvČW�Ys�/�}x�y���L=t�m���Ljko�C��������A�8}Y�|���rp���	�kwN*����(~L"#1fo��)XP�a+E�ݖ���W�Ǟ)��k��Qgf�����4"����b2�$>qiC��%��W5R0C@�j@�JbG{�����L�
��6�Q�+Xd9u{f��ȶ�
��K\��wKT�ԛ�YznaJ�MPB�i�_���HQ��uEq���PS+����»:4�����M�,KY���Q�����/2q`A1Pw�W{L韏����".;��kf����4�ڈȊ:ܞK�%G�xl����<6�14����[?g,U(���]U�%�(R��� �^E��=ָ�����bd�8���G��hA�z�GENUfS��DrZp��A���ÃwɄ0�(V����36�UB"�IBg(o$G'Ĺ��M%V��zU��l���Q>.��_���'X_��Sυ�c��C��aI��Î�=��L� �\�
��P~��gv��q{��34�TE��?c*[�pf��cy��g�������Ua�.������".�ځ�ͨ�t<��ya�M�*]5�ʲ�}�.����BC�q�!$C�9Z�P��7B8�����"qe�~��7U���~$B3�M�w� ���4~p��[ʟ�Nʡ�!8��@gMZ�Q��/��WKYi�rJG�2��~�댄 ���Y�{s��*��L ��ϳM�Y�e�L9��*D�U���I-Z�?"��4%|/��jL:}t���w�ƌ�ӎ�� ;��D��.=���Ca��%LO?c��)e����{�jj0y@̰u�����!W@'��-\{��� VON��\�@��X�vT��G2Pa<��K�0���X� lD�{㋭f�v�}	5��a� ��^����q�6��9l���6�d��Qs ��$�?� �2W��̊R���Vn7�KA)���q��m����qg�y����ȫ���?�疺E�7���8M�"���N���?:���!�Ț����o�����9}��N���ߦ�Я�p.���r�he,!/��R2*"��Dԋ/c"�<"m{PS������[�g�ʷ��ւ��H*�U�/@&#�g3mF�o�v9v1Ǔ����=S��-D ��9BhB�FP5h��֪V��n2�(n2)ߥz&�F}�G���3�^�'��}�����6i[���7��������?��斯�G�g�^�`"ռ�MI��b!��i��/�CZund��tR�j�P�<��D[��Wj�#rn�D�u�N^ڣl�rcS�<u��s�M�d/����<2$���N�UL��/� O|� �O��Ԃx,X{fݐ{�]*���ʚ��'���O*ԥ�Ԋ�t��#� �U����s)����v�/z��"����g��A�����z�6��,���v@QS�Nd�1p!��d%"b@�4 #&a���s�rw���0 i�Qm��`�4�%��\'1��f�}��/2�N���6'mr���pmWYm�wV���ߥ��cA9��3+���0��w{�ö�)�``m/{��ᔹ�z����A)��
0p�QUp��F=�U��Z$���1��Zm'�����%�2����C�0v�_�X��=_%W3�o���sW�oYr�ydl�s��[}�R��k������g`�S`��� ��sJػ��V�=�ěʽ�`~�m�}����(h��_$lЕZ�d.A/����ѻQ��+e�-�TƨaP$�V?K3�7ŏ��d�U���]SW2�S1k���#�>}г��4����@pS��p�Q�8J
�����T��ϳ����c"��D����?� Sd��B��P(^���g�[*Oo[1H�怷9-�&̒Ŋ	X�9Ĭ�'}힢?'��2v����$`�U��J�9+���FJ3�|����4V�5I�����!Q���7��hx�\����A�k-
Do04`0�7î�l��X@GƜ���΢�ײ���߬(�MS���3�DV�`~p�g �ga!R�$��J���fp=g�0T�}��@V5���SA�L��B��Ư��cl4M�	4�w$oWI�Q-e��u�\����(skM>�W��[\\Ze����5$]�������W9$�-��iCo�Tb3�)a����3���Q�d�@c��<����	�=��un��8C?�,*��AN��#~�{����Az�z��af�l�T�J�Fo���)��O��s(��Y���~���o60�'��*-;S]oS����+�6�j�K&'Q1�cfNk��y�-��L�%R��jb��M�O ����d��"�ةL�����g���O���h�j��,k`��ώKS�����R��AT3D`�b�#�����fǷ-�e��D�\E�r��B���Η	��5a�.�T�]�b��94�hʀCؚ'�*�y�ͅb��ʂ&V�h�5*V�.�E?���Ѓd��T�a�I���W���S����o�3&g4/�)�q��:7INx={Ji�����Ef�R4%��)��U'`5�#~�S�kI�dj�󒱎�>� �IC Yr�W�E��
ӨSNUM�(����I�ϼ�T>��8�-�zbb�;R�tT@�6ź��kJ�eR���g ~��E1����%�;t\t1amO��cIM���1vQ��5��.�螠#�����)\,f>�Ѱ��x?(Fcs� �l�k�D�"�M;�++x�l5�G���p4��Deᚽ�m��0�20��F8����h��\C���j\�0��_��Z�(�H�Mz,��y��5}��idO�?Y ��Ť_��<����I�Jy���gece�u3��^��m����!�Bu�	�{�����Wҁ#J@�9ٛMI�G;��dX�~�@z&<�5�<�z�%�
Q���W2<����D{^���&��0ʰ�Uf�%��z#�^��׽/�uQ� ��T��H��r/�^�K�Q��<�"�ߴp�0���@?P���L%��i'���ӟƼQܚf�TE�J�ݼ�a�$��M��|d��K�V蓚�d*쀵o�IC|яvD������ f�a�I���C�O��#+騇d�cpP٣2s'lw��ٌv;�w�#�#@?���ܫ�w����%Vx���ny0�s�}���߫@�6F�j�m9�CG�J������n�v�9�s�T��G�"2�Ƀ��0#M�lUw(s��*jN�e�K���zU��$�H��ڊ��앹�DAĉ�Lw���8�� �
�b��S�u�\(ٟn�۵��ק 0n+C��D:��_�4nBJ��-�<���<j�Z�ޘ��?BPv����ҥ-BIV�lz.Me��?��ZA�.�7�P��T4�V3��.uPJ%����)u\Y��Z��Z, �<�m&F��T�uV ��V�JV6[H(�>�?{��j ��w�T�N��Vx{����.j��!��ƕ&n����6��Z+M,����eS�!Xq�C�Ŕ�tfC|vS$�]~�;�ߠ�SMY�BՕ�$#��qF8��Bq5uO�2�0�2�J�oZO��O{�\]����蔾g��c����A��˽N)N�~+B; �c��WYsA��"�g�[	C�h**|�
M%7�Y���0RU�'�
���F6��>���0����Cct�e!�P�<{9f��)����]xz��l�������56�I*�;��}5�R�Uz<F��$�n�I��x}��u�����V�R�,2_51~?���I��а��;g4sPr��@��Ά^wd�j�	O�»�|� Z&�2"�\� N^�D��]�py[P��m��K�D\ژlc{�0~#Yo���5�ϐ����E�C���~e-Ax$��sQ HiR��HOO*�į����d(B2IЫH5;����e��)��;�Mǉ|���:n�CV�qM���C5Q�W|H
-b��+e��+��:N�0�_~�^�0�?�H	�Q���ۥq�CU���++w�H�3F=L/�Zϣ94������r�	B�)�ć�<�>S׵;�6��[C�
�����-'���s��2��C"��"k2�>s
Ǎ�pq`�+�����H|I�ZO�9C+�ƍ?�������o GhX�/���R��]Ҥ�@����.p��u�u�L�Mc�!<ۓ�Sy�8@3.�j"׹�f@\����;�bO�M���۬��S]��ȗ��\3Q�g�
@��N�<�Ϝ����en7�-�E�@�T�54�W�r�Y^��{7ܙ�����g�������S�Y`",U'j �Cm����Md�F�;�bR>\���:��&����䆱_�J���+�ś��ˋ#�_���t �/��aQ����ì���������)�LB����.�$C��(�G�&kQ���+����A�o��ލ��C�I�QVC����L�7{��͐^���<A�8�m��BZ�]Q2���	���Rp�$���x�lA.s6��1��]�l�J�O����M�����?A)��6fxb �DuT#2l�N ă��Ȗ��v��Փ��RAW�p��(���~�̰)u�4�����i�]�砪���J4�#ka�me$|W�.��N \<�`�Y�s'�-"*@��O᱌{;�>q������va�U���a)�z��)I�%E�q���������9�XF?�*4�Ce6'��dو���ڣ�Z}�*�K��2�@��l�Œ ��!��I����2s^��d�͉(žqY�~��x�bz�>Y/�����x�̮��Yۑ�����n�X�Y�<��ۃ ��Y*��\G��U��.Q*��@�'&
�Ѕl
��&~�;b�M���e[-�����s�k����Eö[��6x�1rR�H�U��6����f���	S�ZĜ�,��/W�,gέ#�D�b���,��	�>�x�����,��~Ιv\k�<o�_�@�)�������:F��XRtKq���rA��'o%�3��Q�ξ5�Xx��q��OX�%�U�0\�v�� g"e�l���^��/	��4R�'@�z>le��ڵw���9.�90���M���=`	$^u�4�'�j����p?�̥���̬'�)�	�
����N����p�_����Z?�$^b�8�
�w��zG@;��HL���В*����ɞTQ��(�� �������ggo���F���E�]F\̔��gv+�>v��%�Hހ��}p��sХ	���T�қ8s��ܔ�۶��7�I�G�ޞ5����V��Й}�lR�"LMcv�=� ���c�'X��7�lS��a�ް�;�N��Х�>_:b�_я�T��?H���7c'̬�:�A�?B��g\�ۦ�R�����0�r�A����[4�M�ni&��i\yPTw�y�=K��:%�Ц��YE�&:ap}��ȍ,&)ig/�����x���Ǳ���,�-��v5?��F�"�3�	:�F5>=_\���(��X��i�>"
-���R�c3O��������3XV*�+`�i��AJ�Jx�^2�_M��.��-���J�LV).WQn��֨�j��Kf;{��it�j��Ԗ�Wkw��6*8�
� �~��r�,9��Cm�(��"����G_�k�T$C��Z�k2� 67H7	P|��fw0z��]�~�h@Y����q�IS)���6�Ғ^���5�QR��fx�F���X2�m�kd&ɮ�&o��6,"i3W�����'bmQ�yO��3�R���ѡ�w�<�A��%[Ai�'�-A�!1��b��I6_�m���%�<��u��}�M_�5R��1��\Ο0�$�{�Gํ��$
�.�R�i4�g��w���N%S/�X�E��yPY��i��E
2�Wq������I�����"�Ym�k�R� �|�(��L㮃�,��lz�`Oo�Nw�7^�"E�/Zx�ܰn˝��ڋ�,A8\����UH��H���I�J�B�����fǥl�O��?Q�B<h|2�f��}�Ȋ8x�{u�S��U9ds�O�E%�Qe�Q<����7H�G�n�I����)*��}���c���:������N5�������j?��j4G'�P�TI�h��Wba�4�waH���	6l��8������mY�\��:�ۑ����D��L��.�4�.ڭ�"�
��*�4�>����~2z�Y����t�hr��:G�y0�Vm�fM��]�A���q�M��#��t��\���s%�#��B�ۚ��U��&.a�N��Y��6���ڿ��� ��:3��+���?K����F��m��Ր�Q] xw�^Lu��0�������J\��*�X#���A��]A�k�(N�	�,�nap��	s��zy���b(��z)A�����p����jL_�</��ܥ��C�1��βOK�S҄=�y���!r�F���2j^�6,�u������dn�9*����J��G99R�/q�z��������R�z��ҕN��m�^Ӥ)�)J�C��CGZL��n��շ����I��ĳv?HA�j�U8yҝ%�J�ҰUL�K�1�D��V��-k2}ڀ��G��,ޡB}F�?qglbZ(�CCډ�E�#u�EQ�D��4od�q�P~̸'~I&�Y��c	?h=!��R����ǇS�<�jq�Z{���[�Eu-h����d�E��p:[J����YgRR�#���T�TIj����8]�6R*�g�G��?2��;JW{�jPbj�d�,��Qٲ��C�:�ݨ�f��ǥ� �f\���Sj�xX56fu�g����X3MO�q @T�6�Xi�	����2��V��>y ٛD�fg���^3����~�``<^��<�t:4�ř{N�1|�@���u�a`~�Ò	0)����}dp��ĥW
�&b��0��ƹT42<ó�0��ȧ�$5�i\$ԫ�u�|�ߍehU<Ԥ�K|"���'����TcG�D��v����z�<�ۛɿ���ǎ�a 4��C��>�ɃH ��/ţ��>�x�Ӌl��+�2*�K�}%V��#��@�K'4����V(�I�V�j�6l.��5{rGXv#��_���-�d��*���&j���2�����1)�g�~���"9��c3���=�i~ֽ&h�U��fG��k$�c��YI ��"�L��`�;��ާI&M�A�������kq̯Yj/��u#��^�BԞ���jl.a�f ߧ!5ZBH�ia
[�t�:i\�����׫.Eh)�w�Y������x4{ktԴ�C�k_3����ˠ�~0�����aǈErvRȱ��%�r�I��.'�0 ,��x���Ӂ)����6���#U���c��k���P]2Ӗ�շ��v�ӨQ����hP�,E���ڪoQ�i |���jB�H��<7p�o�a
���N-�iO�h�G:��O]q|3�6	D��~0�ʇ{�9I����v��˻Sӂ�}���#�̀n����6o\xr%��9r[�,�S:y��k���~�JB��ߟư�Cġ�/n~��X!�gj�pS���)�l��^af��ZT��l���.���*�����v�\��,v�u��AСE�Zh��\��nIx9Bh��?E)@R�jF֌��ĿtD�����}�W\'����Ӟ9��TM�_�N�hA��Î�~�9c���+��,3�	��_ˏx��h;C��e���y++Ŏ_�DE ]P�M���s�O-�dBq�昦Hc�QI���l}��*\5�+��b��ʶ�a�V�Ԏ�y_㜈h7P�?Lb�2�L���a@!�Psg
q�M��(�7Ȅ|�n�e�WA�,5X0�����KG�Ib�����:?T��ؖ�P|B�~�k��E��+>�z"p���z�P�ʿ�d�g��*~s�F�z@K���ι.�L��V$�d%��g:o�*��F�wG���&�������Afs.tA��Z��10U��F=�(z	),��o�C,%ωg�r����C�(�$D��='G��Z����+��A���<w��~ݢ��%a�=q�F;����0�,�|f &2"c��@ej�1(i���}"^�aƸ���(�r�T�����?o\H|��|�>�����&՟�0��Q�5�L�B���u,�z�u���E�<��)�H���Ft���ÊV�N�E����q���g�`��2�g@?�	iZ�����W�} ?qf_�LV�^q+M�=��9����8!�-��5�^��
��C�r �V3V��i�L15����͕F��O�*���s[
�I*p<�A{��p�Sc5��-��">{]빏𼅤��|����A�'ao�֨?deN&p�Q�dFt�H� ��
&�������-�8֤���o�i�ג���*��)5�Q�>�`n���xж�TC��p����F>^Gf2���.53ʊ�Q\4ъB2��K�����s��Q)��1��L�{3|���dt(�.*�i��W���ŧ���@.l��!�T���;�Ձ��
��܃�k8Q`���pP(�|�;g�(;]ӎ�$���dS���Ξ�&�N�4s��w���I�h7W0����DvT��X!�JK��H)z�L�#�R�9�lw|u0��΁_]�1���*BF��Z4�J��O����(Қ0���E�;K 
����XH�(�&��#C��k�iK���E�P�YA�,��ÛP/a�Y��P���<$�4bI�ܬ|��cFWj�����&��N⾐(�0P��,s���v-n��в)�}y���h|Р�#ZG��!\����U��]_�����f2�"U�^�5�nb��Qj�/aK��I��l����p�T��,�j���-����>J~�X�2�0�x.�_!�\:+��[����/B\?��aB�5-��[5�l�[�� s�z��ڎ�#K�deT�sv¦-[{Y�hJ7,�&�� JP�M�]�3�Ao�h�N:����#U��Z�vJ1��4�8���kaP�����!
�)Kk�A\f��ؤ{���[�mT`	L@��2��e]p��.^�0����ړX�},%%!����g+{������2��~,=�s(�\��{��q��-��r
\�$�ҸFx?إD I�!�{܊���au*�J���D�(�����*��>��y�p�� �I����Vz
}���=jN��J�抈#XW���y\5�my��$hgu�Z��
QL"�h�:M�8z- i��
<���M2��s\`4�w�.'�X]C��tÔᨦ��▝�}<m��)P���7���VEx�i揄�s �H:+�_�11��3rm��^dw�
^ni4ܻ��V(r�����~4=Y�7�\WU�g/L��i�߆������7ӷ7)_��VI�v�<�Ր��n~���lNXb�T�ǔ0;^�1�0�39�y��{*|ɻ'�Xܢ짧�ƽ�'^p4�$�Y���f�7��Tܟb�>��]1�o���,J8oC���ir<8IzŎ�^���A�M#=}��U���{6���N
tnSͭG�#�#��U,�f�� �	�h��Bn�1�|>�؈:�S��9�ԯpx_:�XQ��ŵ��i���0` �dXJ�פ���Z;����.��/�ѨƆ@Rn�z��KW���c�-l�KpJ�\�!@�!_UD����p�94��)���Ɍ�5��ڒG��[ݹ?w�ZJc����N1[|��-��r�φ<M
�/>�|��X$���6��ϸ�{AL�O��tY��ds����:��`�]��� �o���L�"#���򟃢�eU��J�k #�lJ�Ƚ�#�k��[i�T�DpӰX����旱wc�sz@�Ǵ�4Or)-7��uxD��-c%,�1����@��] bfVR��r؝��l�2�6��EP9� ��#��UV?˓�UFl���
X�2O��W���BS��8�)�����:����y���C��~��O�\RִB��Ow�.]��q�!K ��+�sH�Xs�b&Z���Q�6�4��uhB���
�?�5����B2��E�;����k�w$��xo^�>/#���\��s��X�wY��j[J2�ȉ��z�y�ے��]Z.`V �
�8��;�v<�F\$����ڐ�b��\���iFF5���K�M���R� �=���c��ުfT�n���`�c{`���U�,(|�ߺ�.��;�M� �7����FY��0��[Ƞ{я�H�ʢ,�;G��;{M���B�Rf�ľC�U�� �x"��-���v��`�3��<���C��ʃW�}��~.�E召;��)��h�����K�ۿ���Ec#�P4�%�o�k�`^P���D��d���x�bi@�r�Y��j޶�ڄ�ܡ�>8z����Cq�v�_?�g<|Y� �������j��N�
2#Ԑ��9ف���0Ӵ�3k���gV*�������}jEz�8���?J1"��C�����ut�g�\w>���|Vhx�x�2Wy��Bkv�O-�C �J>�{��*� Xz��ԍexY?�y|")���\�ˍ�v�Z��Ki��-��$��A�,���$�YnK�tAgY_ղD��l�Rap���e@��\|ݱQtEl4=?�6y�0b��:�x�no�[��5aeQ��fg�l���
�l�ߩ;A��Fn�t��f��J=�͔Ϻ�p�^����g�C?��B��W�t;�����s0��V��H�^"��t-q�0�Fg�&K�j�'����=�X���%Ǯ��c�4!e�,�V��(i�p��>�!�M�'�]6=� K�g�B#�9a�åL* W���;iP�oG����"J�~u���:��q����7�+��bSɟ��@)����)ɱ����)w�Z
�[[Z��e�:��3B��^�;"�Ԡ2׍^?p"��ItY\7t/���y���U�"/1�UsqB
n{~�4g���tf�,P��q��Q0��ԯ�����0H�h$*��1m�E�N�ew�,j}鹎���/�ӣjZguz�������c�'0y�b�	�uB؞�08�J~o\j(����Q-b��ET4>���&$�]=:���\`>���W�~F���`UX��S���c�@���y�Y}�>ve�Y3�|��,��_~蠇��g\���C��2b� �-]|�ׇ�Y���-�v�|)��Ԑ8�Pƅ�)�ʊ�q
s�!(杢xh%%�3��O��h��I����n�~�9�Ɇ�s,��ZVHif �wJ�_񨆥��fЗ"�y����gB��[�>P���We�R.l��xaňs)��V�Ϛ`� 	@ЃF�,�Я��<���<��ڝ�B�Ǵ5C�M(�pZ���O߹,L�(=�|�)`�k�N�%F@�����ЄG�{�ٵ?�����С��b�Mu��U�֚:A���>H��hi&��KRr� �Z��Q�X����l&+�=�+N����g���a#Rvԕ�M�h���	Ym*��.90-.؜��2��Q&c���fe�*L�!�}������zM1��C�~o͟��B�8]�e��fD��~7�6���SS�^3���EHX$ֻ1�� /�Y^,����b��0&(K�r�8��cE�"Z�|F�!h�����H�ӏ.n������p�U�}B�{�F��zz1
y�~�`�#6A���b몗�A%|4����=��+��S
�L� 2&z�؋LF`�H i�%��8�n�mg�:z��L�v�\���}T��&�|�3y�0 �6�H�h�ȄT}���G���Q�T=wr��r~U���^N7:�&���SA��V��r��������#1n�wJ矧�f�q�ġ�����#>���e&���@�%3�_�=ID��o�(�V�'kF{'������ԭ���CͨS��7��)$F!��a�>[$bJ>/4d�P�r��ݗ��<,�.���:��W|t.)�|�ƻP'�T+��QR�#�MJ:���Cj������k�ܖW�/�V�V�^p<C���,��Dv^��5y��R�Ti���#h��kWR�]�K�ˌ4� ��4�����v� p��r��b�zd�U���I�x�%Eǆ Vv�~K���mw��#�!�&��-N�_�͔�!�263Nz�ټ���.�+�uU������n]M| ��_�e���A���� B�l�D~q���ƺ��{��V�@W,�6��@�����,��X��ĉ_��	C
}*�ޞc]�5(׫�y3`g[Q"W6dT@PZЅe3�ŭ��� �1���$0qY	M��mo����k�\�f4���Z�.l3�V%P��Վ8ԛ�g�:�]�Q�Gf�&t�RB��Lt�Ż&�~�6��%��yty�.�-�o�8�q����&Y�ް�7���:t�d_�Vw���[3 ���) ��̜�6p����e�� ]�Ϸ)E����q+vX�	]*�$����_����g�S�z|���ͫK{�%GK�������:�� �w�5�RY�!2U��t�eo���q��:���l�zT8��.����k��S�����V�0U�1����<t*��\Iim�z�����̎1�c99�뮴��,�S�T'���4�
�BD����z+e�q���q�0�f0�rJ淅צS���	8���
�� ۨ>Oڿ���0���
x��Yh�P��aM�D��x
A�SBb�V�sٳ�ל�/j��f��N�}׸��p[��ꧏ>.+�5�d���ڋ�VCv���Y��Ժܙ>��p���8P�_]��.,�������X&PZes��$Y;��ϑ���_�#����u��;u�U��v�"Z-�,v������~x�YPd��9�����i��q'ҙ��~���t�4[�����O�u����@�gH�� �\ߊg&�jr�lG�D�xWa{���{��8Q� :J���Ԕ��_f�DF��J�Y��n̑X�/�f�J�3�o*��ڬ�`���䓸�=�נ��MBA����o��V��YN����`�[��`Z��,�X'ȝ�4P�+��j3�\R��U�c�{���0�0�t:qc�HV ���yZ�ve�<tSܫ�P �#�D�{{8�_9��t:I����a�oHR":hO:�)%���iQ�#E̄��p,|�dDJB�xy���U��-��d&S1�,B<H7tV��}m����,�&t���E�i&�us�dqMt+ ؐ�u\MO%ܚ���F5�M�j���+Z�IZ�|I�x��5�l�l��Z1�6F=#2�O/n��=�r+�NՋ]���@��jcT��=o��hWש�����7��^�m=��3׊R��ǆU�K���fW鋋���b�w��{qt�e��n��t�0�ҧ������_����Y<����~�/	��!��;�jd��G337(i3Y���Ɛ*,�'A:��'G} y����|��Zkݕ_Z��V3��!�QQ��Co�J�9D_�E�_�}�1�d�j#ۏ��f$��c������G�_�V��@7��J��K]AE[�l����i���U�$L ��
}|C�~'��0�s�g^}mX߰�j'H�ރ͕�皾���Z���Z���[�8�q8�U?d����E����`2�S���ǥnT>̜9i9��|P�7.
����s���D'��i�9�jI-$$4y �1?�e�G7[7�7B~�	���������&�!U��}ty!���z���Y�y�F���S�UH���X|A�m�1��b��ܭ���'�`@ok' \�Ҵ1�R��2�-��||B��Ŕ�:n��wto6���6�1��Ϯ!���)��n]�wǸ�Rb"�0�R�1��(
��%�lX��`}�-��0J�S������������N��v�G(�1V5�"��U饾po ���{܄�/J'��\��K� x:hB�H4 ���]�Gņ�	k���9ّ�K\ym�`��uMO6�^9��I��v���?��\;���~\�-�B:�7%�rm荈g�\�ϭ78��;~���`�sx.�6Csx���H��'��罷�:��\�L�¬��&������]P��-��Q�l��� !r@�w[��6��ցUPWE�C+��tQ��1�딊9�0*:��K�?h�A��y�m���S��+^�HU���pHf� ��6U~���
��O������d�.촘*���]��1u�E�o��`J���L@���L�����@4*��ӹK/o���J?F��knh��߷�9�&}��.��	��-�_4w�9� ���O<��~�e�[��xOH�?S�`���7��H���FmY͐����j�>z;(~<k*���_�KJ��B˹|C�����A4��C|�,������ddL6�%H�f>%B��'Z�)���B����ة�0x���u��y�E��4c�ٛ��@{����&�}F`]Q�j`X#�S�h�+'�R���;�:n�<�臤f��G�o�f;��$�:]���,���+�,���@�:=���D =�,
-tPjQ=h��+�!�0�ލ\���Q�z������2��pm��8Lȹ�rQ�=�a�K��)iG���S���w�QL��O��� ������ڭ���C��䱮V��nf'����>��9�<�l�x��T Vf�#�w��G������Jهk9(�@CR�@�L�[qy�t��ޡ��B���{�b���=���ñ�&�3�/j=j��
d�^X��J����14�8V{i��&D�qu�G\��n[��"�+�!�(�0{�+��H����$��ٕ��T�G>���L-��g+���4Jw�ZeO�tW�_�����Ʊz�2�&�"��[P��z�(������z:A���?�m����j�;v+0�?	���l�܈%� �}P�e��?N�ny��ޛk>����a�I]��t�S�
�gi��?��+{���u��3��z7�GҮ�d}���;k���P��V�!�/��-a��#�~�&?�+!ی��a �pϊfLNZw��>Mf���L�t�.(:�k�(���oE��~�Y; Y�۝e��Z:SWkxe�:'XQ�Ĝ	c:4sZ�|y��;��8�� gJ0���
���T�ϐ�k�;��v�v����U� �<SU{j%�-C��s����
�/]�3�F#F�����\��-�sjT\���4�e�j6� ��t�˝��z���g�M�C_�����HUP�*�GHȢa���:���V�����
|�:@�)gB5Eu��j8:xwn��j�=Wm+`ebap c���D�&yx�E��������9�F
b�����Is�x��b���Z�Uk)~S�H����=R�TP��j�<�����������S�9�6��h�g��-����!���GI��&+��Q�[W�Wo�6U'��{������˖$�?ħ�ⱥ8�}���3r��ܽ���|R�%� ����z�k������[a���U
G�>�f=�qcd�{�!��8�%��n][�*@+���s�0�C���k��<��w�f�J%�^\�x5����`� 02B�C��h A���Jլt!��*��+  Ĳt7�3�]��Ej�X4Hp��ckC'Xٸ�=�	I��Ģ�&��lK��MX1�R��(S�aw��v҇%A�o9�=L��3V��|� � M[��m�-D��EMU��T���щU�z�<���~6B�l��U]���h�LR<^C�Շ 7eD;��ĵ��UB~��b٭ut/8�O;�M��Ui'qʱ%Z�r��6��,c�%������?=�ie�O]'A���.�íb���[�m	'� �<*%�Ȇ�N��4�՛���|��Bb���u�CY�dcE�낷�5��XRs
��G��ҏ�N�t���N܁5;�LQ�#�>�u��2�|�����Ws�F�ڽ���j�-2�������x��:�⢫yp1�B��5e�(�,��X�kj���7$����EL0�!�a����#W��ڦ����f��%c�!�J��)nD
�/1����Nt�nV 0<��*m��"��\8Ul��M)&=^�q/�D��{�j��nH��V���(���'⦍SK�j��)w��i֯zc�������<�Po&T�-�E6�U2�p�J���y�u8��{L9z���\�UN��D�z�����JA?���(U[��]"3�ȉ��h@�,�𛂌����=Ԉ��r�5��1���ipx^�M��v}6�����~�R�>��S�Y����"�������68
�?�����ti�>��p��T���U���u��רf�^F}��Rk��� �Z��Ď���i����M��yǦ��Z���YPW| ����[Q�C��#'t�L�z�B0�xt�
�����B2�B��B�����㭋X8Y��[:��$UЩ�U��ŐQV1GrC N�wV��x0!(�z�A!��V�|�ɳ{\_�(�Gd}42�qX��)h}ϰ�Pd��J\����ժ��`�2�	��/���$J�����BS��[~o�~�������?��2pC�����8S)훪�1�-7�;ڗ��H!�n�$�: ?ؼ�����S1�6�X�<�H��,�^h�ڋ��aX~c�f����
�BT�A�� W2{�%,m��m� �*f��_�Sc�
�B���P���KM?�<�B�Z�z�8�UW%2G �`(��Z���K��~��Ɓh��9ķ���>9����֤�U�ω��[����B��;yԛO���:wAe�y���#�����"-f�yBm���j�x�u�W�Pn#e����2>7ҧ���A-g��y���4pI��O�c��بk�7^�"a��?��������-}^ӹ5���v���m҆��D���) ���ue�6�e�k���{+�v�DT*��W�S*(�� d=}* B�?�PRey�D��EA��9<pŒ�xE���ʝB/�0+茊@�wy�>��f0�%4�F�Pp'; {Qk��T���A�%���t٢d;!|���ͥ�Ms����ZK�]ޕ������U����p��pxp����Z�Q��Jc1�2V��ly�a�R�3X�8�oq�<G]�I���	i:�,���� �^���ډ�����Z�����(�)	��|2��F#�	6N�9���ٖ�0o�n�����^�t�F	2���j��| \ca'^$2HV��\ho�8��n��[_Vg�_�ۍ�XEB0�&����R̐�9}���b�#iT;\��0��k���(��nD���>;��W	?��y*; Kb>���X��Ν����kN����"���p2�A�pO��ځ�P�{:� ݋���ߞ�\�3��R~D#RM�)x��W�3	U�z㡕�^�Z���2W��jc���es��Z7C�Ø6f�1Y��Z��)2X��zy��%&��7�`0
E+���U��2@|��kv�}���:�d���v�`7OU+����D�M��)�n�Ύ* �d;�֤R�Ջ�P��"E(��%*����ԃ�#�]�G�nyb;mc��M�_}���"|���;�7g��0w0��4F^��}��L����.: 6�nPl(�\�H"J�����xn�\a��5Oz~�� �z^7�U��ԅ�ץ�q�=cW"�.����=�<H�o�b���w��%
E,Ϣ3�.�;2�	�o�6FS~��)�@�Y
�&$s��U�ڼ�=+�Y��0G� ef�0B�3���a{�uԜ��@4J�(=�<���I$b��f:� �<v֗I>Q�������Ћ��ÑB��Ǌ\xKT;�D�~*u��U���gm��Mԯ�Y��l� ���4��X�[�[�T�߆
Ɇm
�X�*���R�^4������s�6��A�L�]��wX�����MM����^��j�R�a��/���"邨s�+����<;%k�s����=Q=�X��Üf-I��hʁh�M�@���/}�7.�����"(�[B��Ͽٵ�gU�c����x
z�.�pn��I����,��b�4:|�,�o��;�z�u�W�R�`.[�`����f{+��z1�D����=6���$��i7�.�����] 9��t�3[�,_Ce۾�G�P�+dTM�v�D,�#�40�&����B�4���~m�G�"������%OT�p`��� �hĩ���R��!���?_��j�n	�x_2�>�~T���
���'Q��>�j�F�" �H3���n];n���D��w`�ړ��5�7鲈Ȇ�a���p�y9����;O�F��  �\�;�Co�S���������ؒIj<�#������r�Yj��y�1�%K9��H����-m�HZp�dE�K����fA�x���k>5�����ό�f,,G!/�¾������l��OMS����ߧՄDB �k����6��ii[?T��͵�UeB�{\�L�V�:nf�8��Y�Q3���a�seZsHu��~�]�'��i������ׅ)�0��y�b>U����;���.Bz��om���:G,�h�f�!��+�a"��>ň��@Y_Jfz��iN�.�>�$ּj�̼i�XmK�_��tڍ�K�`�����J!�b�m����`��t%�iojA�Hq�Q��sO	zeY�M�/�7��{��35?�%��Hw�r��ֹ�'����&w�[�
��3�H�-�0ҵ�����?<ri�mK�B}�bN ��B1��^�0�U��QT�V�� )+;~4u�x�S@�p@[��}M�����t�婤k�-�0�kp�\Z�Y�1�|~�L[I�IWc��ߒy8%��X�Hx���K���i��(_�?������z��@b�_A9�I�*�&��#�CLHY�LF5cR��Z��d��䂉#����je��g c~ۮK���]�/��9���v��q1Z�[�m�Ǻ�����gw=/�v��2�0ө*(Ky\eJ��3�#�'��^!�-�7�>Qq�@h!��_�8��E��?��{����H��������G��ۣ$C�fߡm6`�������5rB3��[+��c*��;6Ä��wvOQ�ޢ�Uy/H���r�_����P
����l\F|�_q�~|��K���η�> H��h2w�e{-���w����^ �E[��Vr��A	��=y��1c�O��:]֬�<䮙�=������8��(��!ϨU`e��4���]��f�<���Z28��?7���.��������C�|� ��'Ϗ�5j�~|�6L�\��Q���x��^0:� c�8�����hl�\�}lTN��WP�W�y뺘��+*�F*�����p�Ӑ��%��D����^����N�X]��[L'\���q�j=�{|�ѡZ?!��k]:O�P=�����_;���Bz�ʠ���4�[�~c�US���M��E!�Gx�F~O,^��`�љ�0�t�#���r��|��Α�=L�Y����N|�t�id시���&�;�ښ�,[��:y@�3�8Rw�2En N�	s�����Z
��ȵ����B�8'#=W(��,�L㶆�����[^S^5N����^ ��\�o2�Z�O����Wb�eWb�0����LF��9Y��"
��I��Β3��9s��A[�>Cmg�gMH:3|ٕ�W��3vx�=��F��d�>��n�1Ak�r���3����+� �|j�i�&��]˸�E�S4�5�<!:ś�ӗ���n���f�2e�����;�F�'�^�qZ��W��X��&/�;�|�ʙ��f�_\,�z/:1U�T"l������Rg�f��h�{����y���Ab����`�|*��8)��~Y8����"ä�cP�R�[-~^h��]��>����a��6(5���R�
�I��9���B���^��j��&�A��������Y�vM���~l�c��<�k欇�M!Y7߱bR���D/W=��3���gu��@|�.	G� 1����_G�V�#"�~���_U�̹��E���!��kO���\�w�qζu��{d���}xB�c�����R;�6V#�O��N�ʇ=�˺�X����R:�bL��u~��S��e�g�חj�nU�s�Mu�+�9k:Η,�Ú���&���a��1?:�߂�\�~p��C1[L��%t2̟�+0�-����@�P���Vđ^`[����
Lv���9��.
���o�M�>!�T���6tLw�0g�#B �����I�Y�#'�fҹ[u7�M�9�+zhqD�,EQR
�l�Kv�(��&�j���m��pA����7K����� �y�1J�$�M�X��J�V1&��� ���5!θ�Er��{���K����{�4h�L�n���/�.�M#K�h ߍ�VH�L�1|�}F��g-y�)�
�0:|8������nle�3d� �V!a�����C�{�gt{h�gߘINI�p�D˿7���zƣp���Lo{}�
�GM�ZyA�uaɚ�}�Xd]59��LG����@���%�Nz^J
���#���ƀ-�5)�a}�9������O�՛Ɇ�h�0E�7��T7'!�e�D9��@���a���)�xŢO�Ⱦ��d&G|3�O��~���+j$�_i��z����aˍD����B�4�����v�$��� n�4�:�G�铸����
`�U��:��:�rL833�=&��4Ɍ⩛�V#��E�M��Bzt�� O3���,��i�FoFw%;P�T�P��+���ԑI��dN(r`~�����3���s�9�t8=�}3`a�<�0���E'`�
:=�HCH�c�Q�Ec��h����趠<���0�����F �T���{~��8�אy/�����5)|S�M��}�};����k�┪��X�5�{qfZn]���t1O��<����S�u�2�G`|QS}�Þ`�Yڬ(Z2/=ޝ8`I��|1%B颫�G�����F�����rH.�j(��G�Iv#�h�#xm���4jO} Uⱟ�5�����r������bL��X�f�Y�#�\��c����!{ɵ(�����,�Y
����/����M��Y	:1�r��˶"��j�4k���I�PշE�Xx�ϯ�j>S�K��Aiԃ"�}��I 7*0�����뱖�<��DH5�;!�&�(�������"�ڍ����p����W�t�\g<#gEȣ2��w� *̳�/kg�p�~b���6���?uk�����k{=�cr��գ�q1�,?B6�7�}78���F2N�����YY)��띋�<O���6�޷:�������Z���� )mIZ~�c�*I�+/�?�#��*�������B�	tk�lM�P��	��Om�0�6�4�daцL�e�Q��������MM.r�����1LN�î�y�-�f6���[�&��i�}�`� v9���,��l�;�ia �e�L�s+��.�+k�	�����V�":J�"�2�tك#�1�˯�5�b�q�k�h*�:��޺V���=�I�ڸ�|Ϗ�x$�e�n������޹Q� �^���c�0�w�.ni�>�7�A�-AD#
�	�ӳ�
�k_��5�X_�SB�HO�	�$&%��1K��o\T���'�P����	*�H
��vf��io1�^YD�拿J�ސ�-��(�F�3���T!�P	2�|v�v�'���3Ϯ����x7m�p�El��.��J#�+�O/.\�c�6T�� Î�7OE0l�-�ltٴ�{�'�v�vL�[8�� H���n�&��Qꀊ]!�M��G��T�E��G��
"#\�@���BDF�UD����v���O�73o�����a���|;DMF�c���^۬!��20���zh"��3η'�������1�na�Ab���rz�Ӻ�p��9�AMm���5��r�Σ��zGK�������E�L4����F������ �y7[!G�j0~�##�lp����@_�0�j1ŀ�B���0p[d������y�સa��sG|�����颍�A��]��e�C�z8�xg
���^'��4EWq�c�9�TyuSnrN=�uL�jۮ����x��Vp����]'�^-@��	�=�����6`E_��B�;�N�B�R���i��sp]T���'�Ds<��/�4���K��w�~�£�a����r����:;����*f��6��
��\�z�vZ�3*���n�}��d��B�3n��uo����R؞y_g�:�^@����F�K1^攪{,K���Si��r8�@���US��.FY.�D�͖gv�L����Ӂ��!�(��ڂ@lV����{���s���>�jr�Z"�k�����Ip�8�+"�F�0>��{�0kN=H��1�k���Fu:��IU/!T�b$X��m���[5+�k�Ê� �O��%Uol��<��A����?{��>_e-�2i��m?d3W<���:� �n��C�ъe�# >�(�X[�v���v�<��:�v0I�3�(�ŭDt�o�E	ς�;P���@�e�z�B����R�m�w�� �֥I�~c�m���ҳ;�gV�P��'�$@l�JP)���L�d��|�m���:劗�	@���Jal
;�w�!&������w9Po)B�.ù&�B��,l�����K:���:?]ۋ�����O�gY��π�=?�|�(h%����G�x��Gf��W��)�`Ek)Є,v[ǧqb�o���
�Ә�p���S�%�?�\�;񔤟^ߍ+�7����z��<�T�l#"֗ˠ�9슾�YvX}h�x�"�W���<1�e��nʑ�3LWɧ�pg?Q�g�0f]�� �տ��W��2	�� a�~^ʷB���:�[���v�@�a�֊q�Fd�"P�2�q�c�����!дN�j\����\TA��L�6��>���Ӓ�'t���\0�^��/d��'��5�r}{��M��.@<����?�C�(y�;ݹ��{��+!�4	��fUdY4ю�۪{�}�����:��B�pXp�~B�.�j�����Ϯ��n��W��=g7�Yƹ��O�������ve$o�;���Q[�!���[��<�|��c)/S�d_��j|����->�~��컹���O���4w��|�i�?�q����9Vh�۷K��s��U��1	Ѥ<��ȳ*6'�,ӧ��Tm�ڛo7M��}�n��|F�(40�hG�Cn�J��˒����Q� g=;CN�jN�h�
��+���7��m[�����_9���׀F��R�,*v!1��&u�["b2x��o:Q����݀y�a���bg��B�*�z��t7�W1�{9�y�}�q�Y�㜂��]��t�6��>�9Rf ܰYd����6ڝ�>�7��L�[��,��X߬X{���y�H��k��B%����s��?���z�us�U��ĉ&��[��!�_��g�'��F��,����jVHS��ir̾�����̊Rdx/m&�Xj�n���}bF���E?�u�J[�s��M���:LI���c��<�.�r�׻ORo�N�,�2�"3���� ��i��+?�z|qB|�/H�o/$ʏ�Qk��F�bh����N{���^����)�>3�������&��S��V����=a�=5)ulam�����x̯�X2PF7�(�?�ZW{��b����9y5�������nk���+�����R
ҕK���� ��gJ����&^=?b?�/+U�˴��BJU�(F$�#r�gص�!b��xy�X8��%�&- �3Q,A��7��)f�-�q����x.��xE��}?0��Y|��N�	O���u�w`^��f���5�˷p�[Z;�㋧�/8-�lw;�+�6˚���-H��GQ7F�T炍d�]�&C��3�����Uy�� [��z�|�2�F����%h��Qo�������F���� ��; e3�՝��lғ�/p�$��><.5�v^,�&����W��_C'���)�>��L�A�����Y�~��X�Q\m�{��tS��p Ѷ�(g�[[��+�.�rA�|5f
�C�d��5yq��@&;��Z��G(�G.:�Ӝ0g�3c7	�[.�r���a|�Le��6�M)�K��2���+�� ���[�Ouw�����q�	�f�'d��V��ʡD����6�2��"d���-.��z~Q?�l��(ڳ�$\?������N��(�(��I�0��5ҹ۶:k��T�ɗ����Q,���v�G�\� c`|OW&8��P���;E��-B�@�ݍ�$+C�Y�7� @=ZiA��h;���f a(���D�/WU���/c]�|J��ÖD6�����]EV��ֺ���c�>Y��;��gTX[��8��(�d�v�#�x��y��o�N�����^��߶�E��%�cFrz�2�L�G13�a�*'�R�X��Yݚ��rWmݩ`]�g}�ݴ9J�Y���"yd7��J��[6��F6�k��@$zH��������&�^��2|��m����Tp6�/un���J8���Rgf�F��t�&`���0�X~���$3�fTNۛ��<l�k��:�ѽi�#@�n炞D&�z�����*G�9!�@�=���0vZL*t*ñw����6��,7�#��[W(�ߟ.�>��!�T��0;0<#�z�͇�'��06�������3u�T�=��V�_:?��:�ή��(�nҵVKA��)L��^�t+Pi `�<59��Z�8c�"i��j�o3&��Z%	X7<{B�y�ޖp#�J�\`r �rp�]����FV`g����uL��	��w￈!+��`�7�����2#@�Y��Yj��r�p'%vG���<;�C�|�� ���>�h��g�J�R�E֥�Y`a�呩|-Ue����IfVW	C1\l�׍N��&Q��M�:�7;e�K�l�W�K\�4� _�Hy��E�OP�ۏ���`�0���%�M8̆�Vz\&{���ھ>��Ea��Wox�s�d���T������Z
e�Ob���$McY�kF!8)��g�U7���oQI�n�d�T,e�D�����MV����)Q*3�Vz}� �O���v�X��`���"��[7��@؄]��sP�/�ή�G�&*N�/����;~w�V͐�r��4X�mN��ӆj��נ���'��o��3��kҩ;�fڕD�$E2�$D��e��rw�׸@G��1��RWFu�&�X����(���C|?| �I@G�����V���t��Sx}���~��x���"��ܹ����s���q��I�U߸*l�f�����G��A�ڔ"JI��}H����9f����sX���|J��p�|�s��
d�C5�i�H��w��g�������5�L�-YM+e�:�&�^��4���E<\������W��y���0 ��=�����:����iB�H�3x3�C�:�ڽ{�=?_�9��ذ�������Д����������<������b��)�\�1�H��l�:c��� �����Z�C4��mM[��v�9�L����f�MC*/�Y�[�L�kA�^ՙ��38���*�A5�@�6���j�J-2��1ՆCHX�9qЊ�� F�rqM��-d�PƵ��	ë���c=����/o�[��P7d��QZQW� �y��@�h&˧PDEG�A�4x ��,��z�Jia��1��U��EځI�32t,�rop��{A@thE���H<kLL�)�觴�`�lD��.�h�!����I�:;�#�w|7eYb�I��=JM��¡�w|C�_A���dl��Lv=�&z�"�t�/63��I�c������!^=a?r�˫��1.�.�k�:W��!c9��B��S���Xoi��Y��x�^�����7<��ţ�x"� ��8S�ޭR`:��r
J�˜�Z-H��p}��$��� �Ӽػ��l״��{�����p�8���X��s[�5{�z9�o;�-VA�8m�?/b��l�6Vio�3���P�*|�o�����H����p��e��l�#���6�p��/�2v��vI３̿�y"b�UhUQ���9�uΉr�,�Ί����F<`�>�5����oA�vɠ� �g�Ci�nr�ꅡ�MM oCNxI��t�5�1ݑ�:0Qlz?>':��x�Pi\J8���Ӣ8`��rk�BַpyW-oD�n�73kP�K;�q��t9kr�п��@*���F���T��T^�B\8�Ҍ{r�k�t�,ᡶ�?ʏ�s�"�_@��d�Q�W�'�#ν�z۵W5�o���ɢlʸ���M����ɨQ���l��p4��=O�/1�&�P�T5zvB$!�IY	�m���1��4_��q�"���e��O_K��A�٬GCك+��f`����r�!�j���Ё���<}~�9��-�~]T�����p��s|>z ��H�^W٪7ֆ�k&�GO6��J*���L}�_�(@m���1�V�Mj�)n��'�]����a�D1��0����T��xq�S����`tЂ��K �@6u��3H����_�9a�����ܖ4C�7��/�9���d(
��Fb�.��/B����T�x�'�yQ�G�,8���2t���A�/\V8��'��9ۊ����o0e����`�6k{V�m�_��M�`���ѓ��,6(�K��r_ߠ�˟_���w 0'�Bs���Ⱡ���Nϔ;z,�C(Ƿ�X�����R�wc���	�ضq�)��?���"�8����� /OY����|ޣ^#I��]����[3�D�Zg|���l���Fͱ�#��`w���/�`8p?����V� ���^����
3���K���/ʠ��d���Udq,v=�3���
Q?8��%.��fh�8�Z������C��.���W;Y�I��eL������{d ����4+���i*# .ZԌ����U���p�������NW>+|b���,̅��꼠��gǲ��B�oL�߯�ڊ�y����.6�)j��,�A��y	��P�}Z@6�t��}5���O�e�"��d�k��+.gJ\l���l����ɚ�M����- k��Dߖ ė��jN�Ѹ��f_R��O]��QXHF-�\ W9r�	��KĦ��}��d�!�c�`���u8ů�]m�EZu��~�j˼n.����,����៽�_��6��9�f���p7��"bA�7"�Y����	C�b���c��.���[�u�%���7j�����)~�8-��ٝ��y�ɓ�~�bfg����?�I^�f^c�~��s��z�;��_0݁떌��ީ5�Ҙs����.5�����/�@��;w�op���6蠥I�b�����O,��YX�GZqG�덢0��W.�&���"�:��xi��qӥ>vi�>= w_��?[�H
2����|Q�tNK��_+?C�OG�Ѿ(&��9� �/�UA&�D�TD��C&��(�H��:ϣl�����z��ʚx\�L%&x�̣�Fx�*�./�H��i�r�P�0fò* �p�Y|��>FfQ��H�a���lX[��r�6�E�%���Fa	�ܖ�nF�{��Fe
H֞�:��al,X �_�a�~��I�]�\�rn�B�"E��n�S<W�1��wc5��+��tCƣQYw��|E���d����L�q�;�B�;��q��,�Ka���Tݻ_��٫�?����3� BK�F��~W+H�R�E��v�~C�q`�h-�M�I��{�|���4б����Q�?�f��J��Eo�TY��{�_�P;�I�M��s����@75�	~���E;��P���a��6��B����ˮّM��M���ξt,r2z�ѿ�f]/EL��S>���z����lG��iSv��/��_5ш�:�������B��v� ��9�K�����,�= ��g�f��c��9�|r	���4�� M�ȽnJ��Ho̴��=Y�.ho���Tt�ˠ1��\ӆ~�H���|�^|�受�yO���b>������Q����v7t�#1���}!	�L��,2�����Xn�O��\Z_��k�R4�]�^�2�_r�9�L&`h-��L��X�A�L��k���<�G|�MK�
�*�蛱�2��h![,{�	����	���5�; ��!�D�3�Ȝ&o�Y�]-�0&�\R���]y2�k��%j��(��{^���5m��{5ׄ%_e;������Y|��!����9	���6��(ඞKe�~�c����B��쮽�R:Pka�f�160�kF����E�=�k��j���1�3f0X�x�A5��03(B��2���&�w��7�Q���<�܏1�inI��,�b�����*PKux=� ��jx����S��G����A-vТ�����K�ʵl��=�e�c�-�bq.j+��$�&D�~PTƄ.C\4}��qg��a�{~?�x���{�C�ܜg��/l�#�c�L�d6�r_T1����zp㻵8�*�r+i��NUf�:�[�P��bJ�#��0vȬ:)	>�k�Bɩ?~ ���3��~Yua��k;��X�M~d�+�-n�J-���cQ?�N�?}�kZ�/���"��s|�d��8�B�M�^�6.�q�D�����b�`��.Ė�>�Eh������W������'�x�e2��9t�k�y�	jQ�G0;4��t�|�oǕ#]��y�[�NaEZf,a����Uk��+�%\����a����1���j���O::�sǪo����`��⿜��A6��yO�T�ã�ƹ��oRO�ыq�^�7V�@	�3&
�^�����?:�U�Lr��,4�Ȃ����V"�?u-����[�-j�M���]��EAW�� ~�3͟6�l�����o��{�=�;�<~H��r��7 ��V|��ͣ�t*�/2�W.%f��+�`z���>�%*�6m�rͤ���q�	�t�Ҙ� D?���ZRN%%l���]����5���L񁤜��L�[�B���\=�Y~(��� ����߉��Z|�b>��h�ȏ�0���L:O�l��Q�p`��iI�U:����.�x%�-և�� ���	G�X�-����k3��9��$E�d�96�o��Ȩ�7�d�9R��e��H:�:���ēp�	MO�PV���LMl���ͣxx���K\�{���(#�n��7�����N,ޱ
���d$����{���DM�4���m��SX$wzL隡�*eX��q�q7\�H{�`�y;'ΡIn�*jÉ�X�z�f��u�jSlB��z�S�C�'4��Z1���Jc�wEkf:�+�4M��O�����m.s���˞�y�jr,Sc��}��g���VSd?Re
|��K$XH3@?��H���c�>q��Xtb�t����1��g]0�Ex/��l{�����O-�wf�sA���r/*]C�u��O�]�GEk�Z�![z���v��d��~p��bMAo�����27�W�Ϗ�:B��ǁA��K�z,�ĝb0~�G��U�9:¨��--���q��&��\�+�1� ��Am�1{(�Ի�m����O�,ۄ��3�B�Mȿ����VC��UK������Y�ں<�C�qf���2f�`���)O��́o ������� �;���D	A����ɠF�!���v��^�q���	�9G�7_gꅙL��GG���fE0�X�-�I�~����+�v�o8ٵ�����,����kL�o��zT��쮺}���������dޒ~�����������u�q�įqS	�{(�5�7ڛ̨��O�c�4�Fi�xk�����#e�Fࡤm�g���Z�UOܔVx
���95�u~���w�{���f�U�a��s��_j0:l�ܥ"�W��3d���7�5��^ �El��� ?�wޠ�yy��f=�@���[���l�C}�
ZilDtq�ٷ~_Gt߱%��3�A�5�">��b=a�0{�&��`��?��`�^*T��@U�/�ك|�ǟ�h}e�8\�/	��a0f�99�<�ç�sU7��oԓ�Q�[����J����qKl|���jC+�k�u�U}��)�J?���3����F#�HJ��AqIrh����e���熟��r���L6��!�IWz�1�Gp�(G���7��Q?��QЋ�x����&�9繉n���ɶ�l���ty���4��^`%���Z���"��1qIT�6�f/K�Fdܨ���{�*P��tn�z�
�L��m;P�MG��7�3�T���[�I^�"z�АF�0H)�l�����CF䷌ .�q9���V������7{�R���E�ݘ����v�p��������
��0I��캚7�t��QNL�e�c|~��.�}�^շh�ꉳ��jK5����a�@b;�aO�a"�=Y����<�u��o��V����r��d�Ħ�`lG'�X�h�<vTs��Q�Pj��-�c��Z6e���_A����o5�� �[�	��ܜ�&���
D�`)�D	O
�7Ig5*��d4o"�1�-�".#G�Q�v5�%��,����ke5a���$>���Q5C��&�qyY��m�ﾞ����/)�b��U>ݢv�0� fӞg�qO<ّԨs������h(����r��F�dD�q� ���m��nS��h��+_�#��E�e�k���y賌-��B�������u�,�"i�EPܶ�?W|�6��OK;�w�%����i�RRfrR
��[��
�-�l_ ���r�$�x&.2�C���?/\a���/��ZØ��O���1;nx���$P¤�n���+�y3�XވVL@Zg��|V0h��k�b�G�ڪ�[��#bz�x��;�����I�d�ZP�k���)W�r��vD�*��V��B�zi5o���> b��n�d���'P���~A�hӖ���&�cb�ͻ��`Qc�5��2pq�d�����;�����ָx��|��D@�i�T�P��(�bV!��w)"I�5�3C���1�(���c�Y⊹�xt�QA����Ez]o���%��,�)yqo����[݄��h{r����t
���l� �MEN��s��^�0���ߕ���O-��X��I����;�V�R�D0���z��+-���"�jM8��CfS�~���*սɐ;e���jd�+S.�47��fX����x�2�;��k��i�i��(���7�;����%�����u ������g1B �T��0IX-@-�!�r�o�E�Fz�3"�{Oa���e:b>n5��='��Q�]-\E�3�zU����&'��?���!Y�B!�K��O�tzŬ�l�x��e$�� �6\΍�]���qh6�ڟ~�͵����.�F��@#�%��F�Y�hj�E ��$�`}�;+�d�z���=��{�n��GB��2�[cB�u��<-<	���b�>�9֧����{>��8(�l��W��!H��;�*�7?�ZO��,G%��������>��J��O��O�0���x�q��҉�����V.{�Ɔo7��9�7$���6Ma��f�Oj=�G�ڙ0�	<���RK�'~0��7Ձó�P���&�[�b�w�7@vݐj��̆�;���U���#�?�"Ж��/u��D��[m�l�f���q
A�~�0QEM$^�lWI�C��^	}o��d���4@�)5�@9�ˮgd�������B�k�]��+z�3���z���/z���g�n07���Z����}v٤�X�������/^/�ѽ�� �(0���g�!ޙ-a�KY]��9�\����?*��ۆSN���g��B���3���ZͶ��+'Y)�~K�#��/GZî�U�D��6]�]7?ĸ鞱働�A��M}e�?0/�j���y�#��$|7����He�'b��e!��r{��G��x#�����Ϊ�ړ9��22|}{%���Ĵ��P�-���ALUO�!Q�+��Z��v�N�.=�'���zDW^�����FV���˕Oߥ5�Ʒ?�y���+4�m5^+e�܇���$�h�$S|��c"�2}Q0Nē>#��R�T��>'㜚!u6���j���Ċ%;c���!ڹ2�_V*�?���d�B0��.Dnf��at'����c���PzǬ.C�[�k�	a�{�i.[�l�V�M!;	����*$��J�z�#�=��B�C�8��>>�S=J����Ϧ�%�>	��Ri�L�öQ�Q{jZ��o��j�?fl���I��o�N|;'$dJ#N�S"�<�gD3f�H��5[���r>�>��{ 5�����E��tz�sK}/7�.v}1�z4� �O�A�X�@�Z��Ԕ�.A�x��R5 ������O��~1�G��v��@yѫ����N4����&2�#�FZ ��v�R1F�B��H��0������uL��V�8}A*!�U������#]��d�_t#h��yp���ʶKlI&�s�ܠ��3�R���b{�Oԗ� �x���p�\�uN�;e9��9z�uy��>z^w+�ñ�:O}�z�t1�]'?=g��˽�����E!f�TZ�M��ggq��7��l\�����W�-i���~f�4憏���A�˻t��1�t����&��7�&�Z�/�`�vt�7jotvP=2~�WCj��K��`��͠�$���KE�}(�O$x��T�O7�m�L 3����k��0�F��H��hKr���ki>x|�0J��w� H�aV�!Aq��ZPJ�uJ��7S����{�[C�3n�<��R�rM�8�[�Ih;�H-�;4;t
�91�m�Q�Euc�P$N�t3�=vΕ1#�FqW  �*�80h;6d1��āe�E��t>�1�:>54�V��Q�6##��`(�Qv&\I��VZ�o���^
&Y>�+��z�fw�
LM� '��섿x���~� G4�F6i�3Rfx_����]d�/b���yb�bm��S�4��~fëSK�h.q��3���Q(¦��`D�M���}�:z(+�x�PN��G�u$��Z�k:���BK ��~�Ǘ9�,�B=I�tz'�Z�.#L��DQ�]��6-�}�@`�?��U��OQh:<ca���]9�ԋ�{+�U�3�_Q��ǒj���,ұ��V뗲�'V9h���5r�����Q��\���&�>����+ŬQ�����/�uE?]��}�~m�KG��Nb�_W`����]K��X,q�>�Æf�S. ���k+��&K��h ��-�`������,�^���Ӱh�w��G/�aε�^�e `�M���o����g��M�Ѱ5	r�s�W��|��-Q�Ѯ
�Y�H�X3�k�bGoEzg�JW�������3d����@� �i:����|�u���H�|Bu#�I�SA{�{��
��������E�v��ܬӑ%V�=��X����Fe}�fz8���r`��O=��ћ��m.���3����Mv��$ �B�MG��Ϛ�65>���8�8��s��
��j�pV��#�q��rC�jr�d@C�U� �oK��&�}�ɇ�*&�Qd�g"���_p��{���>
<�Lw�j�`X����kN��ح�,��~��/��6�V�^�|-�!�fW� �L��d�1��lQ2�֭)��&GGϒ�ߣ_6)����T����c�l��C����7J,��ɦ�%�fj�2�/>i��s�[Gn26٭���:��pa�^�'0FE쏢��6Ý�C*�zWB��R�Г��Wj�|���G0!DR��@��|�)o�bĲECS�^��Eb�h��ؓ&'5#�h!H�Y���y�� G�K�& �X�<�ߗY6�O6�a��)\)�^���Kz�G*���h�YD��J�9�����W7 "��sĨ�n��M�u�ë{$���\��![ۀG7�+�_:�wl�BF�5�#9���� m"2�KE�wwM�7
�2�pz��16�zS�`(�=I�;�f$V�EaC�Zol�@�V�8![��>��Q�Q�*���LV�e-f����1dr��)�p	�0v>��Q��hN��J�a&��j���х#�^b��
�C'M1Z��tz;Fx ����OJk�k����o�TF��C 6����X3�j!B����t���Ʈ��X�hm��������|��}(�k�c������I�MspSH>���(4T~� ane[*��QG��+XU*�<��Jh[������A}��-,�"��"=�[x��I�����NL���Σ�]�c؋dw}�?E�3	9�F>�j8�Q96���ۓԊ�ϥ�J��A�~]���x�aӴE�yF{��{���w�� +n	t��A�z��K!�~�^N�z���z䀻�)��%#aP9�p����r�,�B��F��RƵ;�?�}aHM��!�e<ױ�n2�t[<T:��*T����S���M���!0\C��*�8�nHPqfhw��8o]��=�@������08�-�a�z��L�ߔ���K�z�@$Z������t� �a$�UrJ&*����__�������x��z�A�
͋��[c�C��c��O!Z��������=��	���&d[�^�������p�ٽ�
ߋW8k��Kn����ύ5���/S��e����'�إ��,[��`�����C!��P��$�@t�PC��L��&t����Y�(U�~���eE�>����'CI<��@�O9!���DTQ<|V�۫���|���o�17)�Ily������7��2�F�<Ǭ�-G��F�fʹ�k��;�Ǭ�g�~�<u���{���eII��,o�{6(���"���t��z���ߖ����s��P�g�G"_��|��~r��_��ץ����*��L9S����G�c���M
�(��3�HR����>�S~T�E�%���n�E��?���.c��w�ɲ1uj�o~��1�b)� Q؄/XG���P
�J�p���
�]���9���~�);�/Ò��/G���� �R<
�v��21t��E�HҦ�W��.�i��Y*�#�M�1|H�)�l����|�d���۳�7��d���Z�|@u���R�]y�/���0�����QRʊ����"��	��4k����^��f�d�
��~R%�~�U[~���z7*���z�a!��f�+t������%�fan���ʕ��u���G���yrؓ��3:�2���z�_��,��	^'0��y��0#����&���{Fk�[r��G0eE�,�Bo�_�Vq5��>�I�`�^�9B�7�(�u|H
��nܾ���N��R�E}�[��C�C!q��� �z�Bw*iKl^�:L�Yy��!����J�SR�B19�}ju��1�}4"���� �~��+�k,G9���X�=o�� �+mYS�4���s�bx9j����3d��/�=�ך%�L|���6L���|�E��4�ǜ����EO�P����8	)Êr�NM8#/�(}|tf�)?�C�!�[)��HDM5Bm��Bb �U���07<�!��@h�F�ŕ�Z�UWJm��������C��ݙ�}�y�9)�������9�W����?y�0�3��\E��z�(��;�P�R�>�G�-�rk��?nkL�ZSd��d|v+p�UF{��_�0Y�5�1���������E��K�mO��l&��]#���)�9M�$&e�]�#��o��Uh�od�&�&?�NJ�וy��O|�,���B���+�:5`w�j��������s��]x����W*��mv'$�4�N�b�'�X��5𘊼Tq�!\vk���2� LF�}����:���en܅���qa�������Ȯf�m�����r��S�.������G����6�q����)s	��%�\jw��A��<�X�4�����G�5f���D��?�J`H3�k�Y����dn�
�	��c�\/�/D�Ӕ<�f��Ka'Ϛ�~�rV��u��q�pe��������v�Ų-��U�EI�o��YU���l/�3�O���1$W� \w�����W�����>��` �T-���s2��M��)հ�[r^FoP�(�����)$3��L��3c�u~�z_���,�_��+�w��v�3�A���&7���e�tZ.����
=�J۠�ޘ7M��,v��WoF�Q�`��䈼%3	�v�n�P֧<��,�0/z�_�E(���{M��%g�\)'&S"�F;������lO�_�u��Y$
��T��?�[�/ɶ������­�j�r�B�غT�E�HNbtU���g.V�7g&͘ �J[B�T��3>9ЗWi�#&dS����Ȥ�>WP"W_��yx+qpTW�!����F���,��;�M����2A�v��3�X��6�\#�"%�>|��r�
'�m�|?_ۘ�"���8��Z��A4���4�r�*Ɇm���V�Q-��|�9��F����ڈ��S�����w���{��QƉU�_��^�$����v<�e�����_X"�1��~�4�@CW�IPҊk��v��ӿ��im�x4��r�ˊY���}�T#�)O�4�1kS@�^�9�ܝ�ϥ��p��m��'�E�܋�h� � 	�����A�bZ��X�`�)�r�U�S�8���zw��Y،��e��6�dZUA�+�_2�d�Xl�	�:��z.�ܟ8��t���zl.l!F��M<����5�`#�Pu�}�4�(�$���q�y�/�Bg���L0��T?��Pi�x�0�E���_K��j��ڔ�9�q��������Cd��[O�v2C�B�Pz"R���s��T��J^QJT�g.��=1R�H��s��h�C�jޖ�^���Ӣ?V�O�� �9pK�O��1m,�� �r㖣}B�5���+�=�Ht1&��^h2Z�wf曊\��.��v͒�g�2��I.`fvEH��{Yw���$��0���ѝ��Y`��{���2pn/�:CN��z�pǹ0W!Pj��P6������) �wy(mD-Q�E�)Hn���Z�v��8Z�l�N^yq##'�b��g�˸6��ˍޞ|����n����U)C�fu� 9D����B?�$�y��hC)��E�� r9
�v>ͫld�tEQGw�AA-�,��J��Q��m����������a�mը����uLY�EwY�8E��ÿ�OO:�pMq�o�`�R��{5��2<L���#G3Nͨ������,@���R+��ȣ��/p.9.BI@�T�t|C�f��ă[�`Ȣ��H�W�]߀~[��H�&�y¤��'��!�yN$A����&�T��@�1� 
�Z�`ф��Ln�XY���8-�1���L�*e�'l���2#���L�T��A���]<]_٨9�_�S�+����'hz�� ڶٟ��2�/l+`�l�t�C&?L�)�ycg����L�����]H�mu ��ѧ�'|E�;�;�RQ���?T��:�O��Ų�����#
�����sn`��`��Q���>�R_K�����4A?I�����ж�`�.{aie��d�Lmqs��c�6-�Ĭ��I���C(����m��б�b�zN��L;k*4��T�i.Y)0�g�w��$�(9���{�6��蝄,�Ν��}�K)u�b��\����('4_EFN�g�b�?�VU8���'SaݗF��(��]/0��P�X��m�
���b�2���_n�� ��Or���5�0�^c�Tt�������֧d��|��4�2�
_P��X#>�Rtl�N@����/�^�}И����=�����pŘXJC�@�-�t|��au�X���S��AI��f�Y�g
�
��w1^F{��&��GH��b��OFp]��B���&��`�`�=)���n�^��k,�G�����R7Z�r�"���$���>29zW$��� Ԏk��=��w��Wv�\��f�N}��H#�����m�u�\x��U�qn�}1�[K���������\��8��O�K�R}�%����-h(X�"��$�s�R�FV�/�)���^!�ɬ������"���C��z����v��J�D+MJ4��^r���b �H60E,~Ћ�Ğ+�##���Pوyt�p���En�9�'ci�)�:zS�����pz~65���/'��r��*	�\�v>SN��g�ߡ�6N)�N��h�TQ���;`���Ԧ��ۈ��6����j�`nԙ�8[wnV�JC��)Qن�H���X)�b����˔�S�B�x7������T����cQ�$���,B�g\��P�ԋ�a��[�� �4���%�d?��9F�����M�z�^2c��Δ�GT��Z�:�-	/4̬��ṗ?���5����QF� ���T�w�g���D��'�)����S��HRi�R�@�Z���>�,)�!�J�`����d��l �D��~���=�5�a�k�V�����Y[��Ph���u{��U(۰���1�u��.�Jd�s�g`�8�?�VǗm���L�kRv�S�5�s����U')ń�y��,�*#1�=��(��V�m�sy�5�t'�	��a��H!������λ��2ȼ��BjɌJ9���.�ԁu�j<V�Az��.�� �abx�E����^�e����WН+އ 7�����6X;#�y���l̀�Sգ��V��f,w�����Q�H����0)yI�3)4M�"�-��t�e� i�T2�!4�����r$ �Z��(�2ܴ*���K�p�{��C��2<pFa�A.M�~W��x�ޤ����ָ0�^4%B6D̀!�VO�$:B卥��%��~�9k����[O9�3��a���A��f�]?���CM�(2��Dr�8Vؿ5"�I�����K�����CO���FhGJ�ȆҴAZ��F�z�Yj~Q���E�	���7.WC�i*/-�OJ�r2.�Z~q���V&�ܫ�uD
yz0���l��`�L��Q���:A�g���w>�Qu��?��%�*�@߳����<QV��@���D%�6���2��v�t���^D>m�� gQ�/�S	�'X�E��(}����i��G�R�߷�>L ���$�n�₇w�|/���, �ϭ�-��G$�� �w����،��r�1�/p좛��j��@+�ͧ�g��!׭=W)} k�;�6�U���(�vԬI�
���0���N}� �I�mL�����!�)���_��b�>�j���9#�>�� b���xj� ��8�jρ��a���^u�H5�����4�k��J���.Sos���![���l�U�x�+�5�hQ�uq�?:1Y��5[��ˮ7b���,vq��,������N�n��B

�Z��k
+X�,H~8T"
v�c���yo���M y��^�l�U ^j��M�{��6ڛ���9**d�ޖǌ���{,��9=̅F�L4�4��,;��[����W��b��v�SK���XQ�Ha#b�?
zı	�����6��/��4Qi�B��R7�Za�%L���&�Z�gCN�dn��u�B����r+��ٺ�x,e���^�X��*O[�ɋΈI��y��O����u����v��>�T����r�l|1]���
h"�ye$����)�66h�Q���������A�:�?��k4�B�1�>�	.��R��n�Q\!�#V*I ߌb���]�ᩥ�v*�5NǄ���ײ�䠥B���!�[���G�J��$RY)u�,�(���m?��� �z���&�]�GR�s��[�DޟOx�Dqi1Ű����mD�F�c�����ھ'?L������e��@�4�t	k. �E3
ˑ�+�25FO�NO��10�{k�v�[|X]�����.��4�E�l�U��L)e�AthVղ�[hش��Z}�����Gv*f+�lx�J �iP�:&�6!�B��ARwVۺ�O˘	�o8�y���^,+�]r�.!\��F��KB74ѤJ�u��=Ǒf�@�w�;��
��T�P|�����	J$p$ȡ��a]7��#M�q���_T���;��`��?J���?�|!�V$��Wκ�u��ݾ�/#�f�
�{�LA�A�*6�d�+K�'hJOKV���*Y�>ܗ{f=�Q���u�IP���ڲ1,����h�e�����o��T�L�*Z0�f�����沒�$�S�f�{��a3�:k>�/v�0<�D�:M1%�`oۺ1%՛�
X��pY�G
����͏��sa�M���Ti�mme�� ��R�܊����Z��|v��:bݿA�O����u�7M1}�r?F?�%��\uY�S��NY}��?c����kC�%"h,�~~��s'���Ї't�Д�vM*_5��t�}'&>���V��N'���)�= g�ֹ�C)����h���dl�nC��6������uE��'�S�l�(�{�혝�Aݝ����t,��4�T��۔j�<�T9+1��8��5�n5�*�I㭥��@�ܧ�q0[�Q��ɺ4,�	���m���l�'B�,-��J����ջ;��޹ �4	���o:��3f��֪���d�
����҉�� �|��>����'euSf�G��DcJ\���]��|o��_�%���Ja"�!k8����l�ki�zg��92*�Y����KLz����
��ѵiK�D�n���R�7�r����JW$��Vn�iJd�3LiM��Nl���Zok�D wj�(c��\�/�˰-�?kIF�!��*��B��	z�lN��ҢDzS����E�;(��������e�c?��Ѫ�wvs��|+�<uw�A�W�#�O�[�c?Q��As���NY��dö��j,M*$g�t���~�������ep�����g�F$�ѽ�Hyس}��YTI@,D�,��q��q9���Gc���hj/�Fs�y���(���]6L�k3d��������##��}%�Q���OçOo�n������db�V:C��XnV�BJ�����#%��V.6��ʴ�Z��\�X��i��}��B�l�"�j
r�e`��%����[x��a�G��0�%}J	.�L\Y�s���w�ǖ��F�e����f�y�Oi���\� �+o�^��!\u�^��?�q��Q$�FErj�J�]��P��
^�ܧ��~F���jQ����WƝj�ߎFǾ����0c��l������Q�?������M!�u�G�g�l��!|�`��du��B~/�<�ok��0�7jM�jf�Weq��C�%��!H�cnEN��(V�꛶��cU6E�������7}��-Ֆdל�:���\��c}��*�㢻M]� Pr��}4��9
�L�S�,� -�i�S3�^p�A�Jm$b��Ͱ=x���Śo�)}J���|y�:�P���.$d��đʷ�M���DĆ��и���YR�{/�PYԔ��6���YV/��a]��
��|�o|����C�IM��
���ր���PYͣtF�����D(8�z5;����Z7�Ոl6���<^a������^�2ˀQ�����}��[��D��)�h��'�o<�������X���;x>�b3�a��r�5�W%�2�ntW���+P���z!NIM��E��$�)Z�+N�A�k��F%��ò���=n��؛o@Ѩ?*6�-5D�B��9{��0]i캽�o�W5����T��s�#j�c�ǩ���A������@��v>&��G�M�4��++��Z3/O�'	`_���|� �uǩ�)S�_KL�����+B� @���`w���v��x�2�2�֝m����.����웙Bnr���a,7����������(f5Q��mB�h���$HkV.��o�+YW�+�'��VXt����FW�*䦍�`��cW/���` /64�p&̹�P�~�qS��G�\��ء�~i�\�?�����T��Ja�$b�ܺI�S�m�&����$�WIZ�N깩��*!ZI�kb�<�{V_Ǣ�	�Fs���%�?���0�N��~_�s� �Mk`p&W�A�L$����m�F������N�ib+��z���Y� ���&��k���ѧEK��v�}�B���uU��rn �*��%W��Y���S�ۑ�:���OP"V��y�����+UG3�^�1d:68D`�6ԁjMY�Ol����,�y�v
�F��yg�����jqǮ>��Fk��*�ԗ^j$�����������A�=���*�|K/��)�Ý���z������L�7�
�lM��D�v�E������A�u	���̓F��52�����Hq�2Bn\�����s���a�L{4�+��i�-��i^%�g�-���	WŘ��n斈1D񁄠�Ε�y��?��vJ�6Ѹ�&��G����{�����������i�C�{�?�q	4ք�C�������:��R���U�V�#��$��O�}�z�<~[���?zBKdy�I(�U>�A!�N��"��o�H�;�wD�E�9H�{���(yM(���$Kȳ��T�
�J�81��`M��&d:_�����N6q�ӡ|�5����7�T���>(�7�P��݌V7	J �}r�4L�z'�Y!��$��uT^F� �?��R�B�9�ਦ<+�8���iYD����!Q_�͔`WA��.C�t�<��4d�k�j���C��Yj�/f��~r+��UH�o��\�{�7�"�AgZL%P(İ��>QpD� S�()�"�%8zE�Ԅ<�˫;Sl��(P����|�e��7_�����h�֐($��V�O��Y��=�hZ� �cp�p�wr�E�)<��� u?�ɺ�����BЦ�j����〸���Ji3H�"<*j��
ؔ�b��N�ֿZE�����[��v�Q�m��mDLbe��������7}x� �����ɖ��i��cC�����@'_����N�Ǯ��#k��;t��@ۀ��mӎ�E��9�
Y�Ӟ%��S �@d���=j�$���_f�U	�P��XF�1��ݪZ����ѩ@�"�� #�?p^,k�0 ]�%۝$���Ur����U�i��(�w1#�^o �޻ܔ5@�ܰ�g���ǅ)�����6�j�I��/r�T`I�30ػH�snR,�_%|��zY��^��=��k�e/���eu�����]��&�ZL�7	�W�x���F�=Z��H%�-o��Z�C
�����eT�R*��Ofn���x$�{�>ϰġ�9�$�ףǁ��[G�N>Y3��<j�'���H���NY6E���v��{f�J��x��T�\�������n���̈́���\_�o�g.k�^x��#�4d�9��.]����{�_|����W��ޭ���Nc�@�����D��qP�-�Qf�W���:��f�B����E!���^8P�U���\E�wQh8�W��<$�=����q��a�G��ޑ�ތ,�A�po��h��Br5xk��H�����t�<�{�m�t���I�H����U���!���t,�tvC�3�Xd�ƽ���9S�E�ǐ�ع��v���f�,ڞQ	�w��aN���52n��<7=̣k@���s֏�MMAtiƀ����z؃���54B-6�D����K����Xd��e���Ry�W�]6(�QT��#e�[0�.�>��̦���=�+��jM^�v��1�SU��"�����
0
�m�>(t�Y =���q٘Js ��Z�s&��b�5	?>b�e���nJ�w_�m�~���«�P}�R�_�����9:�Ɣ3[VH�����ߝ*M�Σo�pu��L��E�����E㰐ð�U���:uh�=���u��W�)Ӄ�l�-���߾�w�q�Nh��Z���8b_`���w�%R�3�l��& ��Z�Z��r�wM������Rj�d�nY��J6iڜ[Sh��]��Fmyf�u���C���'�"
�fd���3G��ʑe$1Z��(�s)v`�
�P��B+���U��M�ji�1���K7�J_o�S�d���h���A�M_��7��=Zk��<��<u)�g&J��T���~�uwFMCϙ1]�;��ES1�s��[L���[���j�?�~��>��I�����V��n"��D�bX/_C"Kh���H��,nrЬ�~"͵��@��s���4��T{�K�$�H�.�e@��Wwi��\) �/Ə���ul�6�@��]pgw��X�`r�A����{V9���/�;���&�U:�M��u7>sM(�gTZW�ދ��; ����g����0{}g���
� lS��[B�d�І��	[�K�����������[��- ʠ�mg��s�`-&=5���|�/�1'��F�:Zb���l����f]�|��R9��-�/�_B>�I������6��S�u�	첝.��^l�����"Xc�"T.�v�T݇�̌%̉z����6>��I��!�b�{T���?��?��:�T����l�P�u�m��Ϣ\����T(�#v�ip��>g����F�V����� T�,h�s��(�@�;�t��&��.�Ә���1��V_�oqC�3o\vC^�Κ��ֹ��R6p��N����>��L�>��`*s!嘃����cн�V����z�Ћ�:2+�Y-�F!�T%��F0ML;�ʴ
�ʨP��`�<��ab���B����T������i�=e�læ3�
��4B7S�?%��yo�&��?���0�W��V�p�	���[�#mc��x!��Ϩn�l3�V��Y�E���d��"�^N��u�G�9x*rnh���C��M�ݡ�jWKK�T�ͫW�/箌��@Ms:�g{�!��-N�ؑ,�,�����8!8 �\
�t/��_��P����W˾��$l%g���l����QBX9яQ�W��e[�CM�)Nzt��ԧ�JRZHh�\o�l˲�l1 ��󻋰(�<,�jNn���b��ˣH[���b����N:��\����eg��TøI/u)� ��GRy�e,m��ڣTMEF��D����s�@%X�ߪ���ا�8�x���Px>IDOщ�%a�Ȋ�U?8���D����ю�e�7M2��^>�f�0�o���nz�4���#��%���\�}>1(��� ����5�OŨ�s��g��5CU����7��B����ͼ����&L�QR�;>�U�c�F����N&z'��_(�Y��n�-nȸ̔(�O��>�V�E���(p��O������E��؍�>�@bm�j}�W�k��������G	���s�x���I�ӱ<O�}���Z���b"��|���&��kI����µ�R;�f�8P@ LEC��^�NҰ�&0�5�#<�M�Ӯ(�T�&*�ͮ3j�6����|��L�얂i����ĵ�d|�.?�XR����ceh��?Y�Q}��A4����Q;��࠲�kЌ�����{!vR/�k��a8��|Εa޲7�YJ�q8��8�L��1x�<3$�)�_�-!�@��@�
�ž��|Ck��l��wa�
N�|��ƈ?��tA�V��]�|�9Z�4�8�9�J�Q����r���Mۑ�``7�|�%�,���'�+���B�*<�<L�B_��g��-�p���ܯ���Kj�؈��5�;e)���fD�G�ml�N���ĺ��	��L�i���@l�X�%�S�gzC�0�r��R�P���^��iz����=���I��;��Ц�`���˚S�)��q	�^��;9��6DT�7����Z%� -��z��WE&�u�(�q�e�M�l�Cٞ�OpN�����N�m�����KÁ��J�̶�;�1�@c�+f�����؂� �e�ۇ"v���	�؟�9�}s���V\�\SG��K&�h��奒f6�S�0p�c]�I)ھX��r5�3-☀q��͓��8����2��s(yX7o<�]�����v�Z|�14ɐSW�z�!�a��t���m�;�s.�~r������g ���^��%=p���GI�9��e�٘?%;í���Ul�-x3'I��b�^����E�vD$'jPS'��6J�1�>J��Io�N��c��h���T/���Q�<�v�ש�^,��6#"��n�.���x`�N�����L�3��I��{/����DC��!N�j��N�%��ê#6�M��b�.�>yNs��[8�d ���\�������Z��-�w\T�����q�@wE�\��h<ꋉ����$A�2,���������~&W�G\Y��J���!bh!k���r���%A�2 �^X�Q�9v�Z aV}Oݔ8И-��D��*���,a܁�G;����ԥs[��'X�&)��B�H-��Gkf3�î ��0#<�lG��7�	�/�٣4/?�3,�m��i��D43����i�-̔���x�8�J���v��{*���6��	�/0i%�B�H�Q�gKT��QS�/0 4�QC8����_rK������Ry]�f���l�}��"����e/�:x��a��c�e�Z�CDQ8 d�P��D9^j��@�+�x�Ӈ��6��V�
�
��Pg���ۅ S�^/�ۥ�ҋ���f��I��(����� k>12"�9���5>�w�<�;�P��
�%�1鑯���	�C")��I =�ix*��,l��kV�q�_�7��	���M��2B2�����<N.l�h$YC�L��-����-8�+���Y�#�s~X���R6BH��7� ;��Q�1�a�1�g:�WՔu��3��K�GT!AsJ��F-�b� �9�_��˔<`��=��@e�?&���b�{����`���R�j���_��k54�i?�;��ʖ��x�)�G'^u��l��8���2X��n��tPn�L�V*��Z[-bɪOɈq�脛#$� �pzE�
�~f��	#���'�|�(4���_w�l�J$�g���[̀� (1[&��X�K)��m\o���Y[��b۪�Tz�0���;U ��7C�p#�zH�8̿C�><%����-����y�>Q�����ڽ��tC[,j�3K=�*~LX�J�T1��0�~K��%o8����J��'��,�r͙\�_?m���ݿ��ni]:�ü�1s����(��\~V%��9�|�\kϫV�R�7 F�g�-��û<���f1�gx�0��*���G�����;+i�Ѷ���9���o5ٜ����"�H��r�){*-�P���"���cIaF<=A]��?�ZmH��i�[�ɳ��c��ݥ5��>��H>�`�L�ȳ�t>�(\g���y���5W��c(�7{ә�
>A��T����Gx���������C�H=�0�#�}�����tT����18��Z`�|���p1х+�b��^0?��tc4u5�Иv8���8�B��D�3�CL*�V�������)@����\0�?��?��+E��A����1 �dm8R�OxC���}*�W����q�V��;N�w�<�>��e�����:����7������X�eOJt=7�����73��σ��1U
t�%� b�N��}����_��z3b?��6W����-���Ű 0m�L��&��HC8gB;+L����]R�0��,r!� ^ߵ/s	�����|���X�V�5��/�P$e�?�Qށ�^���~9]8�^9/���H�th�6�������\N�Ċ�֝�#�,�Ud�8�t��<Ֆ��Vp�$w�y���U#�x��!��ţf��^�2�$i2_lj�"���ֻ!V�$aysA'E&8��#�M�z����ڂ"�Lh����("���:�aV2�h��m�b�j�}1L
�?��e�u�������������������MD�*z� �]�Q���/1��b�N�Aõ	�P�:�ߵ�<�_���sZ~�|��{���-�SX7����"���/&�!j�]�I��[p�,�:YP��	����j�wg(b��x
 v��b�S4�pgiݹ}��� Ѥ�		�­���� �E�Y����oM`Ac�yj�34'/q�X�h*+4�l⹬ˬ�v7$��6ų7J��nc��B��TW�`�z�^��γ��'Na*�#8��Uh2˒9kũ�m,����_|�o��d��՟�n���v����	��W��%���X���Q����̳���(/k�*3{?��u�T�Kz��aq���:'��Q��&_�H��g�&�j��%<8Ӏ@�bS��q�|��) >�w(�����,�jT���+fY��s)�9</��<۷=�Q_ϯ�Vx�e�+���+)�3<^��$B�';؋�������RT�Kz�`߯d��V�����_�����B��N����ai/�����i���E����p���T;��1@ٞ���.�Lg�7�'�`��T��M�<zr�dg��Œ^�����r���{�-��iW���jݪK`-�辖��{��i?��-�sx�Σ���\κ�:<�iUɎ/�%�K?�щ�%�"ȁX�Ĉ��v�?���" jD�r��YG��k��pN�{���pEl�Ê�jЫ�07xI���OXҊ��E*�I����X�C5���T|�t@��UF[�RR2�����:):2q*R1"P�ћ��_~B;�;�Cj_;	,�rHU+�:�!{����M��__��c[�9K�o|\�&�Ы~,~���q/0 T� �^P�`q��m����h��h�b�k�%x�VZ`]_򀰚��)��fǱ'���%�J`��R��Ś9/�f\��~�W���Bo�Ǒ�"'���SY����A�}1�o�c!W����l/d�!Av-�aq֗j*vz	�oI޾�U��E�I\h�%�#�tE�����r���sQ	���ȴ]x���|mzZ��ZgM��m&�Q��}���|>;#�vw;՚������4�ap����:���)�p8���zcx�
)��:�K@�>���6�U)f��d1M9�	F>�jo�6�55��S{��Qg6��պx���h��M��Q�Kn�!��`Cj���Bʳ
����J��ʶ���6�����>C���� 2Ɣ{ѐ��z���?�*К�#X����D��kT�{�"s�0>l,��!xVh���J���zP�G��51��d��"#4C��MDa1���V�wQd�
�c���&Z0�w�ļܛ���5�)M�
j��골g;�PWY3����	6��LU�W�M�8��og�?��ࡒ$F�>j`=�1i
�ݴ
O�P��r̳�C�V�3�K�:�t�(�}��a��GO�����H�Tkn�w����A�_Z���C]�W��b�u�0�ʏ��B��B��	Ę�K����V�lUx�p�A� h����3��K�Y�3��&K��z_�p���V���,�Ea��{����e��8o�:���-w�d6۵ 큋�eR����� �[��_�7c<T|i̹��&x˭�ر���ؕ��݋R�2�U�F�2�-}}~�>km�V�w�ԁ�,�7�ٰIأ� FZ�2�}�r��׬�.���P}��Dڰx�us(�v\1ǘ%�,n,d\[��6���ʒg���s���D�a@�T��k��*x����[�wi����N�^��%T#3�O�gݾ��~��,����*�1p^�C'5����6������}l��d�[��ҧ�j+�1PPqU���Z���.�0��@o���2�����_�JɊ����l�#/�@���b���	G�&Y�aj��`Gp�Ğ6�w�Yt� P ^48�&��,�����S���#ƣ�⮏~pqKޚP��ܮ�Ϫ�ŏa��/�vl~�'�= ݖZ~�������
���V׈�nWaCD�)�N 3�S��OӔ�J��GA�T�����a>S�Ft������Z��U��G���-����o�~�(���e�ә�`w�6����"KZ�
��S�K�$R��/�L�����w*�5�I��_���@P�����>:��|NdL#<�=N#��%w�l)ġ9/����*X��mmLR���p��,��B���m�
k[�-K����X8�����i�~"��s�PN��Vy�2�N�9���a*x���F�&Ƨ�J������h�!E�o��l�+�����ü˝��%�^g-��\V����%�3WV%8$��.�"k��;ʃ��f��D	� >��֓�A�w�Jf�����=L���j҈{�ΉXĔ� r4D��'��!����>�x��"H��4hx8V�ҧ�{t�S	�#���9N�}$$;�jP�%9�[����������j�򦨹��  R4m�S�f��W��6[4[dm�+3�I=�6|�uJ�Y��5)�x��l0SY�e˷���|�v?�R�c�i	��^".&p]���&ya�nM�,	�PE:���Z����q��Y��7/�>E�?D�E��mǿoF���&J���.d��w��to̒�6�H��!�1��Nz\���"}���̳"���Ǭ�^���M:�LW������"����b�z�z�!��d��V�0��E1j����q�-��i�X�[h� 6��)��k�a^�XI��ĳ�r}�%�6�K�,��"���.�4�zriT*����UO+��{�\�g�����NT�y&�Bt��;�LWg�T�r@YZ��Z/|(�:�}�J���`fe,�K �`5�8N�C����of��t���\vZ���xݵ�so���a�4:ɕ�{;�D��k���ftv{�h�_�ʽ��\�GY,�fI��8��GP�ٵ���h��ÝP5�G޿2��[a6h��]P	g�
�ĵ���<1,*pfE7d��v�cH���@�!�}_�_5P�1ii���a]$����}�Z��F��Y�buko~K&&zH [��{��fq�)d��%��[6/�'若�x>a��U|��t �:νU`U�/��]�HZ�XP\�M��5���H�L�C%#����U�}��G�D%�nÔ��
s�7�cQ��L_��55���{��Rz��U(%g�yq1�`�H�R�1�!.u��!�9LJiK��ń�p�9ʦ-p:^u~��*���5�Ѓ��S~^�M���I���{�nΐ��bx��ʈTe1�u%y۾��2I��Z�DH�&����xwC��!X'	�ѱ��T�d���S8zq;�R	���I� 7⤐��  g���ؓ���o���Ĭ��PGc8��V6�p{�hu+ѱοV,��4��B"P���k��+��k��I!��{o�0�6�,�{F��C�u>[r�3T�-6���b-eٝ��W��^0�w�x^�-���한�}qN�[(�K`՟��6�@�����x�5��<��2�6�#+c���s�8_8��|/]��/) ���k��N
&t�zY��kF,���e		������*��]0�M�dK0��U��	X=�R��ϡ�'��j�̫��o�Ǆ�Ѧf�X�|���leh���Oq����=�澏�J��	)	�ؾ���[�
��L�?=d*�hjW<��5p۴��r��� [ L�O-�ʽ|�C��ߏ�I|	��g�BCeMsT��H�Od�� #,�3����Q^$����	����w���!^��W' #�`J�c֠W�5�d�_�3QT��3���|��� ����Q���1���m�f���+�G:�Ǵ������0G����Ij���&d��41b��}����}~N���ۻ�v�ćp�OdjHp8gy�QF�#@��4����mow�"~��������Eߊ쓙ק�k�:b�9�������v��F�!�ZHWA�@�2�򽪕����n�z��7�Å�
i�Q�,	.ȉ���"\�!6���2qp�oT�^1�ۺ�)�	4߭�잍�i$���.`�!�]�\N_�W��^S�}����i(���կ���Z�#��$�i��_�d-$�M�fS86�`�?IF����Qcfzb���7kVt�jϺ�[�M,c4�gn�%�n�����ݮM��]X�7��q��ԛ�Ɠ�o�e��O�Ur����[��`�ú����|E�'k��°��ݕ6���3Z�u(������[�8}�D�.��T��ru�=]�Q�+�?B�GE��0��E�u~���3ی���n�#D�nZ����8���?Z��C�F\%��Ԅ8�[_�c��e8�w	4�M�0bc�$Z���%��J@$ Lx幵ؽf���_,0�$��z)�e�9���
GI�m��n���D�pB���ɌXU�ӧc~�e{.5�G�nn��#�����@<	��aqGD����l8�Єʞ���{j���M���71o,�g3����6��}��W����ԹvST~L����q:DT����?-
�O5D��&�����ߖ�HZLV�y�ڤ���=;
?���ô�w�w�Q2-��J����B���{Dr�/�$V�zs	�BkE{����M���Y���tl�P>�' �s�x�Gfu�� K�W��H2��ަn�1�P���z��g�W	�i��F��E�b�:de�W�P����2���hjh��,�<�f)�f@�e��A��v'�(���� L�$�)�Rf&$�c��7�$�w����9�b��!Dػ�{��e��r�.waۅZ�evXM�j�� �G��_��jܓc�~Cϩ��!>��G�?qe�����ץ�ޔ�7i>)�T��ĈA���,��m�R�f)�*������������Պ�]v+�0� ˒����J-��c,�b8
H�y�|���t4߫D㍞���Q������J�s��5/�1�8������)	8���S0s�%_���d_ݻw}�	��|�`A�dչ\�ʪ2�~�G�3H�c	'<�Cؓ��I���;�MP��u�2r3M�߭\�A6P�v�x�m�3������M��-��Ol���Ď����k-^�}�����K	#���^Hd�	A��Cb�����l������|�%�wl��.M|S�)�`-�Q"ҏ�l��Xck���K�����[�p,
Kbޜli�Hv5�֢�%�x7v��=3��fO����`���I��y��C<�iY5*��F��&����N����T�f�3qO���߻���$��,��3�	�g1@����k��h���>� �y���w��*IZ;kX�2��?񠵦O����?&M\]4|�S� ��4�)���y/f6�t��H`�Ә,�b�1�a�5�,(}��(}��7���G�)�o�Ԉ�?�i��Ɏ��8o�4p�]�t��̾�%��=�?�����z�,�ļ�������N�k�z��ae�a(57����h>|?�O<�S�r9̇0�J̓N���n��y�xX=��V4���U��PQ�<�R���L|W?�O3�3��3A��]6�i��oY��B�~!�~�eOF��4Y|� "�v�V2���1}��i�kV��#N'�c��v�T�m,��E�s~�|sOw��k�jQ�i �T��@)Jt�듨�م,v6�ZvG�Z�˶�p�[�����қ���Zakz���,7���� o��xp1ݧ�^4���5�_I�el뤓�0�U����o���,��4����	bQ{��&�j���q���_5g�ּR��rT/�QCǜ���H	>�Q�RK�]��%��G.�`f�:��P$$�#��o�A}��q?�=��3u����#�kpKi����tC�"�Y��������������P��g�!ˉ��X�vv<Z��4��'�eڣ�'����I��K�7yD�x���^%�s�`��{?�����.�p���ۏ�'ʠN� �K���[ �,z��؄�a�0>).�]k�'o~��Ut�FI��J��Z���g���@��4�?ˏ;�����d��Ϝ���[9���[��6��>80n`��|�K�k����#�߹$V-�"�����Ӣ�w�7T\���d� Xnh(/�v��Q)а��k���5�/0L�`����� ���>^��pRs*���;���r�{�W·��5Y~ޮ>�8��[���E�^z�O��z� �a��jt��h��|:�qP��5_�t&�P���(ۋ@wA�u`f��_����!tt�O��r�,�L5��e��u�A������	�轔Q���.��A�����U�H~@Ld��ur[J�阌�g��В�K~ �q�l�-�s���+7�ŉ��>���f?�6��+X/(��;j	�f&H�����'�y��>X]�t�b�D,�[ZU��I�$k��rd,:|�S�vܛ����a{�y���r�.�ji���=�Bg������i���"��I	�����MH��?mm�|'|���_&/�;��p��ꊡ�� �M*(�8O�3�/S)P���.��kE��W#��"++5�$���u�N^�FdQ�׀O���d����-�hz�� ����+׸�8U�c瞈�X�`|L��z�u��s+�?�d���S�����;��E+�hv-p3�_?vy�4�1�����-�x�@~����$�7���gx�gY�pD�[�aAȪ2N���حl��I;�8�R��<MX�hy蟎������o:�%xE`��%��ΐ�K�����F/�S�u2*3vU��/ܟ0%m���L���"�pw�G�kF�h|e�!�p8����Yot�X�p��Y	օ
����W �~�&�E=4#١ %c^�2J`#���P
4�NJ2A~�L�ωp��OL�z]V�T��q�rOۈ�y8���^��[r8�yk>���f،��;	����sy�u�au�<Z�/i�I@�K`H��l����WAj�C|�X�����VhE�&L�O�!�� Ɠ?N�}b�պ3�Y�RtHU�w�x����N��p����ڴ�ji�^j���+�I���~������#d�y�e,�����s�����|ֹa�{��KT_�>f32��_��ү4�MP0��m������Ini�]�D����'����]��zМc9��,|yDWr~�4���t7&����:,��Nn�V1��V�����j>��)��j���������*AV ������N��;!���B��j:g�G�_�B�? ةU��`�Ɠ��ɇD�?t&*��#����JQ}K���qD���K%Q���[�Iؓ�Z��&ss�R��}��C�=�
�P�W*�����g7��Tm�
?
1����~��$ɰl?c�A�,S��9���h�*��l�>�{w�Oq@:�:��!Xe@��dS��Y�oC�5ʔ?���AS�5�B/8%r�K5���|�,�4�$,-������Γzڔ�7��X��V�����5�?(�b�R8��<3K� �}��B�M��`�|)�28k�[j��3�Y	��ތOj�4��4Q�F{�uѰ ݗ���4�އ��[�� %醿�HNxk����ta����l^�2[Y5�3T��S�)��(84GG]`բ��U����HM�:� �=\#��n�[S�:�3~/3�~�A�0�tYչ�@d��1�pr��4���S�OY��Ek��?��+�;��g�O�.U��'��^َp�8#yL�R������KK��;�x�yư.�h�I�=�{���am�_�#GT�~mg�����[w��r�bS}��.͕&���c�Tv��lQ^k+"���+{�C��ꨎ�F<5���#����Qi��+�q����_��.75��~"9���~m@�B�)wv@e���iGdr��?�9}��%�O�.@miw2SNg�:�`�b��r�D��la=1=)K�?s��g�8��(B��ұ����ˀ4it�aҰ�`Ƅ߲��"���
��2}��6�ܿ�+�,�.�.A��ᝡ�Wx+�C�P�e�����_<�:휉N-0+�E: k$��6/ic�?��
1Y�u��>�޹F�,�Bܭ��;<�	$���L�{�����ʰXxV2�=�v��w���v�_��M�-Ƃ�@����d-��X<��9�6i�����d��@q"�����65Ϛ���k |�ɡ8w�Ap�̾L�1�lG�j�lB��0	{��b!�����<�� cl�4-"q"֗p�͞�#g5���L�
�[�p61|�����ls��@��n���	���>�o��0�u�jH��љ����"UOH�Xn�R�C%	\�(���s�[�⡔��ژ*�]m�$]u������It�e hІ0@������&�5�������3Ty�$<��2�B�V��#���2�'�^A��K� T״B�z�<�R'9�,��$_+H#�Û�\�&�?���K�ZEZ��b���dgS�L?���'�]�w�< h�����ԲT@y�j�-�����K��a�g墅�gLA��U*��P��u�u
#]Ol6�B��L İ9ŋ�z�d��i;�WX�V���fIXZ`��:�f�L�s=��!�M\r���8�wQH�<q�خ���Z����	y*(�n��W%l��0y�/ȌaO�8���:4.���/
�% ��R�/����ėo�`Rm�Fޜ�������[���(���%�P��z�o��=l����> u��a��n�|t7�W���t�����WC_�B�B�������r�`ǯڹ@̾���1]~�8.��g���_�w��]fZ�cz9�q�����+/��FH^.���?6�6��G�ӹK��5����N+�G�ca%75U��i{��/5W��Ӵ�t����.���qx�(�����R�<:��G���!&M�N���l
��&��
���A^p�);޺	��1�u�d��Om%0���
O׻�y�֙�' :�!s�i��NsI���`�͎�`��삐�yd߳�V�DS|���U��2�K@*/�o�p���5B��WS|9���: 1�ns���9�����iօK3�y��3��%�������G�W�
��;8��������o�#aQXMC��v����K�q��x���_�7j�
*��:�*J�s.�`���êY`z�xa��`��Q�Ǽ����v�Zc*�N�-��_�Ӂ����"0���!&A�RQW�ZC����Qp�C%c�>)C�,�|Ȓ�_F�0��;��'�i��ݝ��")}uU���hըl���L'I��h��VA�1�Y0��g�)aӿ����E	���N3E��_��"sY(rs*����{�eIբlR��z�GU���ƾ\�ܞ!�=N�^b�t`���
�#ZO�*k�Ȧ"|��d��K2:�5��Һ��~��t�b=��}�;~�,Nţ��H�;��"W���P�Ns�G	7����0ey+EI`��~�c���q{8Z�/�KW����:�%����'��Υ!dF���:k�-����<�'��O<m��|9�Þ�e�������R�҅�3���)�	ptb�`(�ڢĎ ¹ ��_<��,|[�Oo�u�L���И~��3�n�`��d�XN�2~��c3hL�{k"�e�bi΄Po�����o!5i{��]�[?�'�P����Փj"(��$j#����^�����|0�Zu.�/��S�YD=�\B�=�Q��}�Hd� �*�&����N{���<��%/�b����D�播nX��i��,T'������M4i�QM$�������!���D'i��s����CoS �a�>��ufn��:WY��p޼�, �f �����?o�=����	V1 ��;ļ��:F���Ѵ�ٶjR����F!.}��[�نp���\b�IK��ov�<�]۰����i��#&�n�P�z�@�3�c&��o��x �-��(��[,�0O����� �T����������OJdL��wȡ�2�
;c`g�5X� ��%G��X�?�Q�;��~�X�T?��C��s��wހ�O�.�i��R�Ly__߷�X�v��ḗ�0�F@�?�X	K�@�\7�����ΎÅe�O��W��ӄarT�|!� A�_�%H������?�П #A���^� !=�j'_mcS�
����bEoUv ݈w�����s�I3}�?e������:_�!H�ΩQ�6}��ހ��R����N�o�J� �-^���_�.�Ѫѫn�:'eV�UN*�o�H��tT����T�3T��?���I8w�r��yV����AY`O��Sh�&m�o��9�D�MX�����U|\ñ?߮����I���k�hYZe$A/������V�?��f�79�&�=��TD�8����uD��}]��K&\m�+�h�q��A\��Km�kcTɵj|̌kW�Ԩ�_gSf�bY�Bkj��L��4��f�D�Y����e��b%�I��e������]Kf��)���Һ�S�&�Ki�`oO��H�=��V�XYtd�Nv�Ϝ���h�ӘM��<�K�m%�|�?Qh!Z[�F�~��%J����{�vz`-R{c��Jf0#�@�)�H1`M �*O�$<��3E��VF�o�*�K�:���{\��ğ������%�9[���G/w����^�����.�a�/�WJ��\#� >o}�s\%f�>��8#k�T�w�#��0RZ���� 	�_]����B�;=�t�ۉ�z|]�DC��2���Yrش8�K6�&9xiP?��ˢ��,�j��]6������EEǢ�g�1q���7�$⁚~Z�ɝ\��
��ئ�k���:h�y�zg��T0���1�^f�SkC�8���C�����Ci�_�#(h6��O�Zۣr:�jH�b�U�Y��X5:J*0J�3��Nɞ.gԘ�Q�ݎ��k?�ţK`D�>���>�~I�����t��/�1ܯ�K/�<%�`����ٚ6n;��S0�s��Xg΢\IrfL%b��>�k:�߳?*�1�zO�ߝ��o	�}|��k"d 5Ҷֵ����-��I1g ��� �c���<J:��2�%�z�G���}�����z�G�*a�������u�z��-�b����� �H f����jsEv��s��`�a�8Z>s�S��
�����AK���I�|j�ww�7P��| �`j�1LI�d�<95�w1�(�i�O�O-B��!%�%�j W�����s� ^*�{�(�T�c���C+�@vGiYҲ4�VR���ް���kYnf�[Tk�E����J�Z0a�9�?'t�8y�����[��9���b����q�1D6o	�7���jD⨆���uȫ�:��d}�[�� �Ut�r�`r��G$x�{��xA��+D��\ X'L�8R���ru쎋������q����U���ky�� �`:��A�{*���\L�+� y�n�*�qMC����e6��*\�3��N��S�*��p~+���/L]�,Y����u����N�2��P�H6`��q(��ǲ��^gE\��Ċ��6�Ǵ�R��LC���ڔGlu�V}�M�5.u�94ɍ��fZ͊�@�HFh��+[��Ђ����a���R����"��m����$���ہ'V�>�**����[��H�����j0J����Y�艏�AJMms��V@'.R�ᚬ\mG�{x�֗z�����\ŃZ(����t��al��#��NOZp�¾I�i�bTZ�4��󕷆�s���Y�5�̃{���,n�\VSf�-ꑐ�
���������h��L��Cdr b�3����u�Wall~�Sw�k��Ã����SWe�}�̿�jWM��bfe�K�\'��r�,|�3w��X����5��n���c��s֫	��y"�]�N�W2��g7��1�R뜰�{��T�6G}���w�7��?�ֹ'�i��Z����,`�un��p^�_7)�?����� ��S�4B�h�Yn�$��3Dz�OBv�$hEr�r�eB�(B��Ј+{�=&R��5 f�"���=�w;N�z���.�}��l����ZE&>+��V��f��&J����TT��E
�(I��*���2l��{���o32Xrya�A��S{9l����q
FD��?˿�r�ҷ����LA�Ve���j�㖇��(��N��@�T���{z����뚘+ *7T��E��h�B+�b�ӡ@W��7�"
ܙĮ�Q�I���"+��תH�����"��#�2�"�.J:�)���,o+��iH\������6�c.�;=�\���� p-;�g#�9 �le|h��}��@p����opN!<� -q�W &�X�E�ߵ롥��+(]���:���?(���������	+���(��d,�20`rT��$(�X��t�Z�5���V���a*��.�_":`\�#�Un7�U���c�f��hio�pc��>�g0��"8qU!��e�~��kB�Ȫ�O������X�B~���O���>G�����Ҽ�����f�w����`1�57��#��?�g��(�m�-H�LT�ڝ�I�
!*����%�}�#���:����/�������҆������r��5����Ag�4[����W�?Xg���~�?hMy�4�)J�I=������c\ʆ�>�M���ׄ.�,�� 	�>�����E��_�UU]R��0ˤl�s� ����:ĵ�Z�,I3��_RԾJ�"��\&V�;�����v @K�"��6�Ikt<~���4�^���֎=��k��ZǍX�0J=�J�0����3�G�dW�Mê��a�9��A�[�
��߱����C"����L�ޜ��hOY�oi��j�}��.}r�0?c1�!��NYN�T�P{�FT�PeK/-�V,�Ği�U]�B��1&�����S�/�uD� �y���^�g�O_#hy�<�p��ɫ�
pв]��A�~��"(~bv%8h�zi��X�~L����i�jȤ�*G�?ؒHR��5�]�Q�,f�k���@[E�Eo����z�3�����=��R�'ʬ�&�냉��u��tc�KX��Kw��v|얈���.�N��$�v�y��b�q�(=��9+��1��z/t��$
t�fSn�Q�Cw�d���Lp"���r�@��u�, ����_��FP��<<ҝ��>ث2+�����:;��.L���m��t�W�LA�^��ʊ �r{8ߠ��@SAZ��ͽe����#�l�m~���K���eʋ��DؐwW@$�