��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�_���v��	�������d��i��HO�4�H`���ul]����_/�>5
uUQc�)Y��B_Z6�07ó����ج��@��(*��9X��ڐ$U����	Y��D������@j��ڤ1b|���`�czI*�=��fZ�,���[
]���`�6�/2�E��W�k���WQ�\2���[sJHoV��Caꏐ(&:w��-gL}/�S��f�pI���o$(�R��:��zM����/��KLj���55q��ƙ�S�4R�b���o�<z~ �}Qs�o-�1�j��%�Vp�I(��-G�m��>����>`��8�s��	l-�(����B)8�K,���R[���}�)�\�g����8�9Y"�@�-<�Q��b��]L��!tdS�ҋ+oE�
X�>ς�2W8�H} ǻ@��_��~���?���N�U��j�ۑ��HHW�o͋��X�͹ݯ0c�֝q�Qr���_�wN4,�uOQ���L�ur�)��L l׾���r���BKc;�e{���l����K7zFq�M(������ ��X�?(bu[@�^�0���.��>a�"�����!�>v����}�/��}N^1S�޽Vj@�9�ʬWG)li���|Ě�hN�D �O���,2�e�MBtָ��O�����L�t���z��fdEl#���3b�IUq I�:��CYLL{.E�4�>0��q�,Q�ق �
�:(�!t���J�}��;��!�m�Vf�wK��r8I�#���jwT�f�]�b1�g����)�j~�C�����²���<��__.�2dҵ�v�./�$q�u2&��v,J�kE�꼘[����
(�����UpH��ɦ�D��*+��������=�L�ox�n�K؎f���w1V	Q�^Ia��_�qJ�5�Q!_����:�����G��l�A� ��:�4^�d���gJ� i�A(E��f�܅uM?���(��!u��*��-���*Щ���߭6����l�6�'-���:4$����p�t�c�%�Ds��
[m6�w��:�+щ�Db� G�i�lam���5j��Ge�~,Y��1��i�B����t#yɸNJ�4;��U�~2ʜ�[�	$=+x� f�M�[m�]��	�����E�p9��a��LmL\h����������@�j�vj�D�S�WL�ny���&z��߸���aQ^���A�[��*�2���p�[��$�va���A�|�	��
~�2o���p˛->�J�3?�&@L��8�ڵrֱ�s:����B=4�3AU�KYи�~<j�� ��:��ӊG���8��ހ�F��Q�`�^�H!�>�&�z�u<P'�5r�P� I�hX����773�՟�P/�$	��i�V����������k�(�qN+¼�s����;ɋQ���q��.,��v����a������=�ᚼJ?E��8�48��lv^'(��(�gA�zS-��Y���S�[�ޕ�@H�]�.��Z�H�杂o:��Լ�|�5#0�#3���D:rM<zb���3�p�
�R ]��va0���8��c[V��$�B��1}Netm��T���*s  (?Ð�{K}1%I<����@i��$ˁ��� q�E�x$�!e3�2�1	�.�d�аZ�w����-@Z�m�G��`
;F�t���Ė�6
���Kß�ٿ�eN/�
�Bm���n{�Q�&�,@���}��,�E�í�Dx���9*����-A�r_�M�>L|C[l��ڥq�.�����{Nf� >�O��z��"�p'L�PN��-c�fU!D�[D(녮�����^����Dw���*��I B[���֟�	$�Q�%$����q�Y�ǬyX3��m�O�?+d%�'w"��lc��xk��q&�Yݗ�;�e�HI��Te��M��
����_�X
;���QTR�pm�E���V�ɸ;�J��r�0�o*M�Pwm�K����>���o��	Bj�/�K��fUVT����9͸�H9�>�&����~qRjE�ch���'F��	�-$D� �)D�EF���ĮY<%S�E��t/�P��KX1�9�Y���$/�`���*��T���'�e��	+3$f���w�o�8aI��Ԩ��4t$x���J|O�p�2/ t��A�����7Ba{4-�pN�߂Ѵ���\g�0E�4G��</��Y �K��(�:��ѷ�]�&𽥌�ĴPh�O�Fel8���PcC?wg%t��vH�vfi�� !�]m�4�l����?�k�<�0A��:�4* �ϖ�$l+�������]B�d����"�DM����L�����7�daU*r�r�5	BI2����C3����;�VF/ۙ�V�"A'��E`�.����:�9Ӣ���ݦ���	����F�'�I�ޖ���+K�d�ac�O3G�n�Rq�q`�����}�~�7r���� ɲJсM)꽠�?-��R�p����q(��5Q����M�g�X�E�˘!�4`��'�/OzJ����8�a�j�I��#�����7�w$_�� ߹\y����߇����R��@�k�Q�"d�� X��F�{�0m뼳I�=����;'��w!�I�F�T�\0��r\�q�yh�_�_!�6�oO����~s"����\<�v�ŢH�;/��l�t0��C�7���1P[]/㋚�;�U�_��
dh%'�Yq��#�F�/��T;����������-AP��MX����fsg�z@�����rn��\�t���^�Y˯P!ڎ�}����Y�x�r>�Ԏ��o�ā�/���"�V@zᅜG�Z��;؅�L�����yH�eψ�</���n͍(���m�_��Á@�b�>5�\;���f	!�tih�C�޺��͌*G����g���B!Hޔ�[rB%���})x�A�:��4�ӭ�q�W���@���R��GJ/���W����&��z�$����O��M��X�l�}��cj/h���4�����u�B%�zN��lPwDc�S�Q������d����YV>|���d�̵#�'�8_ur�@X��mԩWDK8$4��1�'�FmM.Ƽ�am�Bǚ������a����AN�s8[a�O��X��~h��8x�6Ԥǘ��.��E��+��l�3�"	��0  �P8����X(�k;;�k'�CLE֙�s����[>���؁1��,_A7{i8dGj- <ǣ�<Af ��^��B��7yE���e��Ft  V�7��d��-�@1L����=��-@�Xzn0��b�
On�/}�G-��E (4&`E�����͒őt�2�c(��@���ԥ�{Ŗ���|Y��a)��ˬ��`�](o$SY�qE�K*���9����X��2Ͷ���/N�F��������+��`�U,���(-L�@]HӦ���X��{�*If���ߒf��X��A�*}��~*��D�/�i��ZS��>���g��;J��Nx��v����-����@y�Ni ���;�L���~���ȥ'�����z��;AI��5��ڐ�8��EA%{�O�o�a��ꪏ�
 ;�N��� p6z��¯�ȫ�STH)��ـc�����ݙ����k�"���	��lS��#���;�<#����J5�82�ݚ�C�,��rz�)/��CT�eBǮ!/�
"��na\�s�%��iP�j��H��j��q3,9ݩ���&�"�?T���Ƃ]\��(�9F�l���j��?=�`�=��?g,�G�����w�}���QX���eI����S����`�8ډ�_jq-�_IMg�%��}�������2ؕ��1{�h�+3yE}Ӡ�>�&�A����ԣ��V-�C�<Jd��%����jL95}&���%�"�������R��%컑�J���9>�]uBG�$1L]�f]�Z!�e%k[HͶ0�@~������߸:2�����~���>섑_�;k���<zq�[�N"��3��8}�KQ&���8oBX�߂�bqʝg3����l*8�K=!�ݱ�e)�Jmˍ���3JO�#���M_J�\0�B �)����f/�~��sbԒP5���`��-N��D���%u�nIVV޴�,f�|%�Ls���s�t�����G�7`��=���KS���ɳ�T�T�t�UND�Ъ���?}�5�QM��U�¡w��>lq��T2G`��`t��^�-�U��P�EP�|�w��ª��2
he�M��ߪ\�v;l�6�E�/�˥:�\�<U���ī��-ںQ7��Ed�,� O��9��yb�lU.�
� ?W�u1���a&�8�-,7m�K	y�#zS�>�1�	�IF�����y=$W��|$�Îޟ���m�W;�� ���x�#����N��8��Si�ij��р*�;��V�|(�/�k��s�HmQ��
��Ϙ�Kz���?��Hc�qRKj%xV|���t�l~��V���Yb��������P�n��kH�	dD	w��U9Y�|�\>��=8��l,0�Y]^or�*6+a�f%9̈ȅ�Z��N�3��Ռ�<��c&L�j2B��b��"�~�����ظ�YȀ�=��Z��p�lB�n2��[L~�(�e����5�	8]��eM��2hһ����+OOm;�n�����v��"7�����-�MZ�f�'EM�W:�y�$\|-���w����\Q�������nn;L�1��P�%E|ʥ'r��O�#h4Y��N�r��	��U]<wG"^%���E�T��/�Y��G��>�1�σ�=�;ز��ʑ���z}=P��J��i�ړsAb߳Y�3�2������ܤR�E��ad^ޔ�6@4�B�@����%;��f_c@}U��&��g~М�p�dߘ����,�T�$��uZγ��S[�-�u�M����)�"�vO�Ҝj��s�3�����_D^D�ͼ����W���w����1-�B�㔠4ϽwD��U5T�r+%jB�غ�J�fDCP��6 `�����%WLcZ��L5�����,�"Af5~CB=$t%H���E���0�~����_d
7�t�����v��Jq��{�k�Q�����굪~(��
C�X���P^_��c�}�`_����	v�om�h2>��C����KvN��l�P�������I*kwb�>I��0����ҷ�#���p,��O:�+�14�ǆ��N<VZN�V�dZl��Y67i�&%i����-����G��0���,�촼�e�`A��p(���J`���,N��ƈB֛�s�tizl�V���]�p�&�SԞQ�w�烼�F�����@HGQ��o�7�E��/��f��h6���l����-���[��4�T4$�)�KU��˂��7'
a�eh�Q"sqU���.`%2��?XG#�:τ�Υग़�p�ZCb��:	݁��դF���P����s����8�o�+8%v��Q��K��Ӈ~�\���^`�����Q���H�ܳBi�.gaTfOQ\U�>M�6;��z7�ֲ�C�EYq�e��9�[�6NM�!��P��ֶ݈L
��N'_�e�jy��D석��[��J�ABk��|~פS�3��ÍEx?'�r?��d?���>�.zQ������ܦVF���@�;8�<��{&y�!;�d�ciD����X�n��'so��S�����C�2f���M�k���P6�M���,X�O����]�q��6c~��)\�hU�ŷ��
->��=�G4��߂�څf	�T�]ƱGI�ڎ�ļhMU��s��>I.гM�����m�%<n�F7�;�V��ٟ�q�_����{�����;���WjU ��� �'�]V"�f�β��,���O�q#o},�^c��N����x1�`��O6f��j�>�́�:OL��PRn*��K��̌�ߵW��x�u��SK�TF�{a(�s��=�T���M��PI�b�p+� ��c6��|������*�Z}�ᾙ����u�t��E!�`c-2}�PP'���B��������� ��#�a�]hnge�ׯ�^Ɍg�?�9�`~�ň4k;���\EMR�k[�:�s+���q)�qfѰn��92���A�Ĳ�X����#�)mG�N�Z4�ʊM��S�Cl���~�7�/��V��U���E�uV��Ғ��[�kc���>�7���R"�c_䳰�ފP{��h�>�2E���!�zhz(Ԣ3�<�����h$:�ɵ��68`�$�X�\��1�Q�)��4n��dݡ��+���.���G�|�K��]�ه��Z"��B�=�*N�I�o���z���y�<-�J�p�.��8���#��Qg��:6q���P 8;��	NMQ4�2U��%�6���u�67�:ַ$⫡q�5$����˸�G�	*��������e�%���Xl�gΆ�@�(�����z^Ǚ�B��w%�kO"��1:wgP�Z�@N��n�~�Fh��AYѶ��ι�4L�r��j��2]���0��a�Se�����T��7�l:2��}i��}i�$�2�j��ٵW7
,�|��}����5�H�CeN�>���Vw�Q�P5��fhY���gh�okq��ڗϙR ���ժ|7(k��#-*��i����\|u�[���Ԃy~��8��6}T�-N�Ȃ�-=���Je�����X�ˮ Q�~D�o�F~�XP$^T��\��&C޶xl:����#�S���-�iI+��Wqڽ�Í(�60�#��&ﮂ/!�W�:�n�x��׹��iE�^sHe�J��$�4x���P�w�����K��\a��2�G%�O�D�J�7����ȝ�!R�;E��ƂI�D?������6��1�5��C�$�uVŞֽ���/5�:�,9RsA�m�5�Mh�!T�������?;yx��B��p��Wx���>��@kr�t߶cLoW0��T�Q��U��U��A�Q����M��͑w�rʅ��^�W�lI7���N�ȩ�2�������77߬��֤��h���OO����L��w�Ʒk5���>�O�zU�~Wc�(㮈���͊�/��?�l�������B����S*3f��FT��~J������4z�D��և}?�׀�Y�T3�w�߆![z�����)J{'֪���~N���I�/��µ��>�~�� �����J��;�n���%���
uޗ_�(	$9,���4�6�q#�W�/�������,c���ZNg�2�qKO�.n}_�wO
����n�|Ӥ�~➇��N�BL�����`V���Q����l�ƀ�:L���2�j�~]�Xrg�OUU~� o����ʷ͆��R���v�bX8>�${ ˈ��HN`�R�*!��Y��::���	}k���΢o�T5��)���Ud6	nf�v6F�د� ��u�Ɋ���g�vz9@t<Hkt.�.�pLU�B,Bo�	��q���r��6���Ԓ�j�-��O�E"�G>��%���Ǡ��LH�;d�p]������Ij�[ j��ѿۮ��	/�7|\J
T��GܧxA�,�O��%S:kP��R{����*��Le��3膌�!��#R(��D϶,(���<mN$���I�n���A��K�AAt��^�H~�Y���R�M��,~ÃEHn1����������^��C����M�{Na�C�纗Z���Y�V��+WJ^�<�l�\��>���`�P7y�.�ƣm�5��T���P���pVC�{V<�
!���<�1Ol'<y���m䌫�����"�|=�&����K�π��ǠZ�<�ۗzl�?v��ck�d��gJ��.����Vy�d�'&��s5"��f}����y��ͩY#Z]�W<S���A�:��FnX]�`{,V��8К�(z�Co�Y�J-�����,#�RB9���aM�Gމ2w����܀�%��	�����X�֮(�&�k�^��KL+�Bom�S������4l�FsZ�w�,A����s�/5y��Z+��nt�!�<H,�<�\�|�:���O�i����,�R�,��`�MX8bt�	7���q�w�XQ��k���2g�����v�}�C={��;�y�r $�R��El��w���:^�P��+�Fr�c���
��B��y ;��K��E�g�B��'8�7�H�?�_�9�lض+Ŝ�H�q�������}(���4B��$�鬫rz��'o��,3�#�hRKP9L�D��IBUf>��p�*Dr���)���whܚ�:�U\��/�i'��^p)fq���O�Q��] $�rnk��f����x"p�T���N䒀d�,�tu�`a7d���F�C_����,�����\�4֢ނ�W�My����@�g�'P��iFj$�uv�BQ��*3�~�[3o��c5��v3���~4s�m� �fOD�	�v�<m���D�Կ����Ŷ6�Z��;&p0`���%6����EAK��<4���==�C���5�~�:�N�a�E5g'�hzӜ0~%��щ�� 橘h�#��p�N�ج&!�F���}�'to2��/�w��	�=m2툕2�� 8�n�W�+�`��ż ��UӉ�p�vg� �O�O�R����햖�u�Hn$�R�yӲ�`���m��*��� %a�ܱ�ބ�}�B��ɬ�m�f�j0����<��LF?����&���&C��<ð�xSV�B��<z��o�8[�M����v6�Ua�(T��WN�ܽ$x���4=�xn�^�״�HҲb���r5�hD@����;��()�� �+���f����w�A����a��C���I��1��<����.�Q��/m| ����'�֡��5x������;�2��h���ݓ�K=��k��S E�M��c6yc}�W���R	89�(����_3Z�Q�n5_6�Q����c�>@�V�-8(���)��۹˟���`E����ss����<��/�^vrK�/ӥ�|��g"���㝄�cp<pj�0V�o���>�p�� ����+ͼ����9K,]�Yo8I��D�4Կ��E�^��և��~����r�f��w���)CZ�\,+B�>�{���p��Ә���� ����v�>�����l�#�4g�$��1�K�MZ��+���n��Y	(J��G����9�<�������]���4����#$�x�Mp��
�1N�����0J5u�H���_�l�'f��
�%'k������?�k��z2��410]�Z��o��Ȇ�U���%�"׈sC�IX,u|&ۗ/<�M�6�EF�G7R���þ���i�zو`�G�P�YDGyS��I�Hm-�,EMɨ9um���w��tf>��u�2��)���:�.�RCهJac�O
�� t �i�c��%(40�0Tp������3c�o��r<�$v�K[�4��3��qN6�o���������<,2��ݽ}Ju�E��D�sc��Qpw//Y}HUٛ��s+	�Bh�����fcG؛ع(v�Ĩ�O^x*��.�Ĉ	�F���e܌)il3 ��t%��)R`y4��R8�zq-�BDN��N[s�����=�B���bQ*їv74�=M�BOzk�b���N��&��B���|^X��	z�����t�!��(����A>�֠�c���J�ew��x��u��	��� ��*����2b�w��5ʉG���U�i���1��|�.��!�2�F�uDK��n��Q8˻��Fv���r&���=bmg�DU���RմŞM�[��I�xu:�<�	n�`�X�^J���KY��A�d�����)���y��Gy5Ѡ���sEq�NoљT�^J�)]{#O����\�q��E?�׉/�󟟤��Q�{o��$ %�9y��p$H�>C��9z�j%�� xP�u����!B~�IN�l�q{�l'��gU�|LT��>��<���\E&��ռ�_��<�����גD�c����S@y-��s��֗�v4Yx�����r��[z�ݵ�Q���/�I�?:%	��ڪe+%��kr_gf8��!�9Z&YE�������Xܞ_���%�#�(w��P�X��,g��_"���G�~�$N*���u�܍[��{ E�\5���l4�F�Y��U��;o��5��/�Y��	.���0��}� 74��=5�JW>݀m�-m���$�  K�acY�N�r)at�d��M�,��˴�g7z�[_p��~��G�L�aG�7Y����rJ&�c]�qI�!w�VS���)���K*�݃<�}SA����B6����n\)�A�H%��aȣU�.���׻s��1+���;4�{�5��!{v����*C}PV�N�4 ��ɏ~DGL/(��I�'P��L���zV��jEl�)���5�����![&�4�~Փ[���8���'���"�HP��[�ͨK����OVz����(�����j���$y�wi<O�Ts�ܐ��F���ױ�k��û)&	�2��<���00���� ��R!�s��Gm�v��e�{�L��X�7�G���PU��R�V��cp�$�:_�<���+��"|��P2��#��� ]��L`4��]�Yb3��s#T��ԇ�5яl�'I�q��:'I��rn-�phu?zO��R$%�r�J�c�}�F��oC;Y���=�
;�	���sP�Y-R7 A�;^�`�ay�kP��>8
&�T�]x���AQ#_8$�?^����	�\ïy��N��}���mn&r�(5d�&B�%h�~E�!6>��	s�����V)���B�	���@]FMi&�Am�f����ݩ]I����r�ک^0�:������(�`�ঋz��3�ROr�M\�q+Im��9��׾0�V=��ͿQ7$�GN��r�@0p��\C�c��F<�u~[:��m 9�f�?(CBL��K���J�ߵ�P��g��$����O�l�;�f:�1r���ݻ���9 �����GQi]S<NML�s���y�ņ��(	+j���*���=P���p�AT��l�Gu�u�g?��T
>w�f4u�L逢�Z[PWr�k��&M1�`�e3�ʰqJ�V�:W+6���]��>1D��I����N6��*0zyϹ}~6���$�AmYQ
=W@�J,ܚ�f���i����������T���_�����fK��t��j�˞(c�� �X{�}���$rH���;/�l�b�!&�3�C��`=�X��0�O1�:H	] VK$Ip�\	$EZ>8�!�����D�s��_9.R��i%Wu�9+�m�.�X]��Fwc�[�Z	�*��f���ZJV�#�e�t�i�ƨ�L�����V�aI{Ծ�`w�-����S�X�Ŧ+�3�t�����?e��vƠ g?f�y		_#�L(2�^]s|�R�>̟zUM���J߅ZxzfG\A�_E����젣���\
-[�x{D:xq6����$z6�;�C�c�P�8d�|
�_ُ�˰lP��Մ9XcF'�=2Z��jm�#�m\@�ݚ�Y�Ľ%~�ŅK�\%���S�̀.�,
�aT/i|�?Ue��������5��A���z�7lQ�}�ԥ9ވ@��Ԓ�%O��<��t0�X{�q�+[��F�:<�����\�68�����-Ҿb���3�j�E��q�-&�������� "�g�b^�K���U<֫�B��	��t��"A�d�j��amy���,��WL`!-�3EEŸ��_-ZzA��K[Co��3{`U���}�t�Z��*H��H%���| �ac8�L$��H�t�`̝�l!���g`,���c���~Ů����}z��/&B�Ş�H_�hB�#��� ݂�V,`��s>6i����Es�S�N����-4���ܤS��ٙ����%�n�y\��;A#̐J��u�{\;��hn�Ĕ%M��R�M��� ������n�$sVw���q�*hz��D�P�Sż��:x`��f�:zFcj!�c�p�\�4W���{% z�Cj/l�٤�-U�c#���X����;U{��.�-R����q��6=�-w�>DI��eI�/�6éʲQL��;��j�w}���AS�d9�m�m|�ezKc�~��?����p��eQe��
��>�$��6��W����T�C�~N�J-���OY}NY�?h�6�V��f�����u6���x�&��ý��Ws�U�"�� ���-�5T���BC9ȿ"k-�����=)l�p^���!����T�I~7�n��|Nka6�Nm�:����BPSK�Jvr	�B/�6d�x~�
��ߏ��8��8s9��L�#+��  Gvj�*��նo3��Ψ@9B�.�1�$������%5�P>��k}V;�	��(Es�8f�3¶�3���|��Ϙ�"����:���+�C����!�m~P�e
Q�����c�Fh�W���'�'��n�Q�o���W�ff�Q(�U{��+tVs�C�aJxz��3��@�b<zw���h���:�qҲ��|�Y����Jw�p�Y�d���:4��P�l#:�Au�Y�,���� `b��/�\TUTtذ!`_J+
3��|gSH���Ռ$�~����{��#6�e8����>V�_�~k,S�"��Fvk7j�H
��4s���9�]g>���2E ԩ'a���&��0T�:�/NN$��R��~W���f�F8� ���7=���6��Jj�����$��?K��3�	�L��;�n���.)�qv$s�{�cCt	���ahlv������
X��&6��l���e������F>�Xp:���l}��t}x�;}�*[{�b�iH�ޜ'J�H��v:�VjB�3)H�I��F�W��O�#=G��G3g�V)9�����2nR����*�Z�&B�"�y_��O����Ku�[���xI��4Y�n��ѝ���!to�����Q�=MQݒdkeE���.�1��Z�L@��X��)�4in��
^,X�Y 37:N<�������YN��}�umd��)a�e�w*-2���<��!^��輒*d����(�QqbV���w.����\&5�=��������Xa�?Y�^�3��?����%.�5E�?�S� T�
9Q�B}i���8�baLjz+{��+n+�����]ި��\�}1d����Y���`��c"�����[�H���|�������uR�Cwb+�I���-��
��$�Y��z)�/��݆d�!�6f3�)������jG���u���^�9����1���d�ѱd������z��[UT��Eه��J$s	?���m?�O���%?1�ϰ��F�p�lˈ.|�a��.x"�1����]�Y���M;��&b�&F@n/!hk��FR��:c�=8��W5���0%��)֦�U ���T4�[{�#���'ܲY��M��V���Kf�j�#�Ѐ��&��o����H��"�"������1;gE�q���Q���z7`����嬭��H��4�IE`W��Vq���6-������3B�U�3�CƋA��3-<3�5/D����L��(��'���u�2�/�S�Mi����Hi�\�n��$!l�?�E���d�W��q^/ �^��X+��V�TO�44Y�w7��놅|�\�"��A�aͿ��+[?Y��%��W��#+��A��@�0���31��f�ǧ+J:��k�<Q��<>��I{�|����W,K`^�,�sF�	�,�\$٪�֒�җv��x�$DC�K�a���#��Wk����ަo ۨH�j�T�5Ϙ������]�
ZY=`w(��F�#@6��b�.y�$��lw�e�CK.+hYw�gP��cl5#g Z�E�s��j T���ѥcGzm{�>�"��+.7v���>�2N=�ߖ�Wމ!�j����1�>��~,RaNh��'7\����y�A43/��,��N��l�o`��wg��,��:`��gsVO�+Ų�:ٕ1^��n<�����g":�o�L[u���̹���_ŒͰ�Q���ҽ�y�7Uh3��(f����V��B�^�4G[��ǽu�uz�
U�`6a>�?�M�̛���Df��e,Q|�*������,�;�vRA;y�#�j�S�o���5��Gٌ���6s�W��Ku|���'�H�M���Y�?�Z���m#�?�C?i�R�q�pnѢ3#�h�@Cg�����K ��gp"�C���d0,܆��5� I-�X򣅱-�$[Coej�cDo�y:��ȹ|����h�ܢ�|��b2�cW�A�q�M���Ĕ�Q�}a8p��w�pY��:��KB���pV�3�F�zy�,Q/�%A�3����$¡�~9�M����iy�9`?��8�,��l�0~�������.yI7��@�f�R�Z$�4?��ر�Cߧ� ZD�tJ{F�g��-ɯ�,g�K�T��x>3�(���C��u�|�j̆�]�swu�0{���B�)�.MW�S#)��d��OB�������N��V��-�
Giy�=RKe-�s�Ee �~����1����S��0��Y�e��V1���M�H;<����-p>-�R����y:��f��j�����I
4��6H�t��P��td�hF�S2O���s��1��w�)y��ce�q��-���h�h��Q�rƙ�F����C-Z�
JYڿQ�nk�K� �-V�SA1P�'��. �V��6;�A;�"=t��}*$��^�B?�2� ��p�~�������V�7'8!ynǨ��Ȕc�q �C ��j�-��WJ)0����	j���8�OB 32V�봶��������w����5j��
�]��<����Qb�fe��	�F����xSp�*���T)I���Gu����AX��skS�4[#z�����Պ����g�o���|���ә�[
�2:�1c���غ̦���R�`��7g�n/�	OZ<lWY�E��jjɒᏽ�D��m��������.�S|��[�ҥ��<�9s&�*;���N �b�+����6*��Cة�,=�NcWѧ��J4�q�렽�	�e1EK��Xf�˾����w۳{���Z:-n�2k|E��Q�,e�FT?/�Ա�ų�dC-O#/z'���0��J���ZG�W]��c�������&�!��y��&���#N�)Bw�H�
�V����0ię�,:��n�T���L+Z���}Ƃ�~�f �D~��ܞ��\.p��V+'�бl�`0jjZ%xcr�q[�~1���;��u�6�)/y�%�0髥�����Z4�K�50B�y��:��֥���@�02^:adN��l�i��黠G�a�k���@o�y�B}�<@��R��TV }��"��aC�	ꦿ@X�.�)�[��8HSN���}1�8ѓS�R��_?�y�����Z9t�9�l�i�]y�{�C[X�a��7�4$��E��|���H�^J��k2�#62Cc!��������t�y���j	a$F|=��x�-*v��L�Z�$�-
(
�T��-�Q+����0@j�b+t��^�bl���SP�x���f�%�M䷾w�]��V_-��/��c��a�ډu��=�YҮ<�F�! sa W�$�g��)���������T-�L|_��Iڭ�Ǻ��~yO����?��v�L_�����{�#
i� �B�&�� L�O���=>t�	`7qouC��X��K��!v�u���,��s�d:�n|4`�׾^�gڥB�����H��2�*�[�@J{�:����bաn�-���܁pZx�n
�J��IY�s�=3�`+��
SRԣ涿(��ܬ�1�Z�:ڹ���Q��l{�E����[�۶K�z��S1^��3}o��Ds:������������qJ�˫M��F�rH6�Z��N�A^�;R�>b����.j�C��|�fe?+U�~$�պ2��&^�|�_����������c��]=g�yvي/����u'��&���D���*	K~�jޤ؞�C�C��v�(�c;-	���-�f:Wn|�LZ;�D&��&,�Z*O>��.��Ad�r��ɮ�X����ܝ���l*���d�[�,�OQX.�&���f�T�
���O�_> Ē�R�E��.F��u�6�:�'�1|��z߫�ֻ�!�jT��U�L���}�MEX-:A`$1�y�ө�C]��躩��U��}j�lݣ���A�j�<]ӄ^M��U�1����elz܊��B��W���}1�|Fb�m��̡��Y7���ۂ���S�K#I�'ﳤ/q��̧��z���O�� ��;� F|�T���)(A������0XH���z����I��%�����z>`�YR�"NO*���l-+.N�*W�⏔�͚����K͖�`a%f1T�/�T^t�����!vb�Y�W�#1�ټU,|�2*b�D��P2�ά�;�Ӹ+�1��|�MT�[HBPC��G������	��<����_k~�Ճ�L�A��O�z�`~�}w@��N�f��ݻќX�e��"+�rD����FH�����y�z��D_�i4 ���S�\Wt6k��� ����ܰL�A�_mJ.���wПr�1˞��M��'�?��Ôh��Ku[�v]\'ƲH���3�j0��S8�0�zU\
���	��pJP�:͵��7��`��_,v8�>V@���4٣C����05X��,̠�	Zi�[�i�W �p��>b75��s�u�7�Ǩ&���T#)�p?�.��GD!o���w�R���X7��9_�`�({�,�qMnZA5Ta��($�6�v�Vl3�Y,�C�q18�'sy����ʰ��-�����HPص�n�����t)g���4d�b�aǃ��l=�uǍ��%YKp����>�����N�_ (�q�S���An1aH��q�qDA[K��Φ7WV='=�*z�,�u�%<�R>���8�`��ԯ����K�k7��[,Ȥ	�֡�6�E��3��'���8�����ȾKE��:)�m�]���������"\�sS-��k���x�g�	���s���k�gqb��m��q^���o��)�`@y��3FJD�p�����!�+�>Ǵ�V1����`��
��}9k��#�}"xO�{�/-���I�� �*��=6��|h�v��i��
E�H�^���"� Oh�R��'ݚ>+��'}B���g����xb����rh6�u.o%��z�_�w(���PD������?|i�{2������3�w'��9I���M碻4�GI�%��&�\`��%��
�-qKPML�:����q:�!�R��6�=��暄dxi�~��[풒#� Z9�)?j�.j'����?�2�q�:�a�."�,�����΂�:B��{���hƨ@Β��m���&C���e�8<�a֓U�����Uq�EF��9=מǬ�)�5�S����[��2��)�	�����kE0��΂���(ޡ��#@V���<�I����qog�CV���+�����]����C7刕,��?���)R3�8�9EilH���W �zo��R�	<�����(5�i :�qLi�
)��`�"H�:�	�[�P/�}!~-�B����)զ��u�T��#|���/fѷ]R���dWE:iO����$�O�-�!G��C�)��1hg���A�K�,UI��[��7��ܱT�Mi ��1�*a�9��%9���>���"$�rV(��I�z7�t������`�fk&rg�ɩ5n��vY�z>>�Z�R�0LO5b1.{{�.=�wj0 
	$2��M������;����7��ŢH���hM��7�f40���b�3�<�N�87E��(�ʕ�v�N&s?��@��dU^ₐ���|Mߞ�H�f#��ߩ-���)�*�E�X�}v`��������(CЭ=�#�,����0��F°���Y��u�|ŧ�A��^O���<L?��	�J�i�J/g2U��6���Ң69����I1�c���Z�?�Hs�a�-'4�إY���\����p����q���B�f=KU@��*�G(����]�I�q�Fmed�0ƣI�lj�,&��[m�;;\��N�:F���S5�C�������6$X�3�'�a(�!=A*��B���e����i��QY�uhdlKcո���V��h�6�oTcO�4S�zJ�������bՇ6}�3�i��b,����=[���Ng˨H���>���D(y�5��C�gs�]�Oj��	L�HI����0�)�FfB�X�W\q9��|�T�Y�V�c��s#��<jw����v'1%j��i(�����Yȳ�����N�}~�_;ݢ�j��ȉr�����w|nuʝ�.@jL���IS��I~~&�+W꘷VՒ�����M?�s�p� Dȳ��j�Y��6�8lٶ�0�$�\G}�,��'��n�'hc��}��N��S{E���d�[peu��D�);�Iϒ��Ga��U ��Ct�݆d�p.
Se�z���oP�*;�-���EH��k��-9f�\�����{����#���7��!����0�5vY��rA��"Ԉ�������xyJ.n��U/�q��A�)褵s�ZybZ^,O�!	 ��!�ݞS�B�Dgi=�PS��a�9�t%63	��ou�2����+yԕ���q���q�i�R���,�$�������W�z��M��Ӵmj0��\n����8�Z����M�ƴ����|4z�P�ڵ$�](��뵵�V��x{ ��fq�U���\�嗮�x��k[U]�]y��cLE�^6�$/��r��gM�<����TE�k^[�n�_t?e/$�*���abA����7�[,�m��^�p����%�r3I�
kh�Rd�"�BC�$i��غ���G)\����h��~|7 P���������4���p��G��6����{g�n��'�`���Ķ��O�)�VWᵄ|-k���)1@�AǕUr,���Ύ�VS.�Z0���1~�
v�2�cf	�/�!vn�8��ø�N�I�%�4]�Qt��Gv���:w]�f17��?x���7Q�>�bqp�s{��)?��O-{��8�� ��M��L�1DU��np���0�� *n�G�+9݅I�o+ZͿ�������^f��ր�PC��j��~'�͞�T�<����oǎ��19�W��>Z7e�/���6�T���5�ҕ�j�����c�;9����;C?�.�_C�te�nk�_��5�rp�5�:٪�Hj��\�8�_��r�I���21�xx@Rl��_�Qҭ�tF;�ɳ�Ӷ�-1$I�}'����^ʃ�2@:���z~s�e��<Y���4�7�c��<*��D`�B���K�<U�=T
��������;iMK�t�p����W��HkT)�l+��Z��S���}iٌe�_��x��ͮ�u�c��w�ģ\h��+��MÜ��a�{�ԗ:��*�
�|����UM�mTY�y�TO6��M��Lm�ux�"C�W�֨WY��/�&���_�:��8!��S�IV���w�>e�6������+��}�>Un}�rEրC}|32�j5�*#r1OXH~yR](��f�8��<��m��l�j_4��bܘHi
A��ʗ� ���ȫ_���3g�ΣkB�MDtwiJ���~�Y�򧙓?7L�T�!`�`t�l�t�@� N�A����,����]{ŧ>��R�K!�1�Vn�,>[��E�`D�z�ค��V/��,�{�����S�:zR4��#o6��io(G�S}���%7�����Zqų<����%���;<ύ~�� \wڵ����#D��s]
6����f�m��'Pq�&��:��n��	h�O�z��	>�=�2��.m9���.��j�	�}�����0M�4�"��ܩY���#�r�B��Jk=OϼbY�!m|n���Va�}Ƨ�@��P7T���I����"���˖���Ӷ.f�h�7�[��K�}�"�G%�[�׌�3�
c���]�"�����w2�$�"�����.�b�V���WǣA�����\�<��)T�VT�g�]輰ǆ�q��Z��I/Qz�4�sJz�XIJ|����3�����n����:<;����%�м��jo@C�T.�@4�а�Qi��RJ�����i��1���z� �{e�q�fǝ����8�X�`�!��w��,3;�/ǥJ�%��̑�҉��B����C 4/�W��R��{oIđN��%}��׻���!o��%w_fBF��b�fx�y���'!�F�+�ɹ�6�|]6B�#ěJ̯�����3�ɕ��)!�4L@�_��0ۥ��h�����tQ�b��S{l��K����b�!3�I�s)h�7�2C*��!�b�Z�X@�rRz~z�	j�3Bk�^��Wf���]nZ���t\WtM�,R����0Qu`�׊�����v�r��~}F)���C���|���!��^�*�4��6:���y8޸��+I2�L�9�4 x5y+��ι,�w��ێZU9V�u�5�5aT�	�����<ei�J�&�/�
pPC�H�j����t�Y/����K$ܫ�ޜx@y�)��^�q�>��k*6M�P�HO� F=���T�	3��Ӧk�`�I�g�x"�T�$�W"8�o,�	�Ѷ F2$Tko�6��u��zŤ�+N�.d��)R���
]q*��Nu\�Կ�$&��`*�3�8a��p���U��.�=�c�#hlUn�Øו��d�/2dŻ2�ka�'!��$�g��7��h1���2k�	�ҁ�`U��_�V)	6�H�{h7S1�q��'j�H��1�Ղ�G I/�H�%�6�D�`��%5ó�j�;.c��'+["-�L/��Ual<
�}�]����RM��� ���#���w��?��V�i��J+����f(������U���ħ8ė7�e6#�<+� �Ԩp��u�A%����{����8_���\9y����e<��3�$�;���!���:<f5�]����s>�{PW�Xb�o8�E���8��0�8�XZ
W�b2c��u��'ᮕ5�B�t	�񘠣a��jW�}ob[����}0�%Z��s�e�f��ji�y<U_B�!��ao����?�.�J���9�e�˂��'dZ�^J�?���D!��dmY��j�pOD?Y?&b��N��UvO�e>�XO[KPg^�o-����&9/��`�YY�&�xC�����
������5��F���k�[�9 $9� K0������Q�����(Pe0���Z�p�K3���4}V�A��I0�`��i�_Bk��H�`�c��u(�U���N���ƛF�����1��K���Er\�w������h�5 '��'��U
�l�/F�8F 2�(K�W��RRV-�q����|:���;
�u�{�pi�q� @G-Zn]����
_p����-[rm�̳�׻{�o��u��}W��J��b�^�|wz]�E��.��h�.j�{W�Z���P�8ox×δ��ּ4	��b�1��k�����*��)n������{m�/����0���p/����c)T��bDn��Ϊ��S`Z'ڏ[�8�cGᆬ�����Il��܏�#q�@�̟�ʫ�))��.�8���v�� �����<�w�4��{�����W��g��y&�H%4p���ݴ��Ro ����za��=�la�ɺ��ʣ���.�a��u8�C�W���el�9o�ũ�}s$-{��j�|���
>�yv'�v�N���`�Hs:���j5�ZT�Oe���Ԏ
�S����ɉ�l�̨f\�����Y�9��E<򀗀��v9�'Ny)Aj[�@WD�_Ndb]���P�s �����J�,����A3�˹���<M����r��Y��57�o̒C�e;���u�<��C�'��m��o͂<R:�I�H15��q0��-\=�JF�-2��:h�\��|(�CS-G(�8��xv'@�#V�Z�X�L�M����l���F�5�.3�Lʿt����=��l^����L��R��_�S�������E�3j#�^Z�0���pg0
�l���&6���D�[ <w��	���2$)c��rk{�S.�f��7���k���h��-�/Z�xS�s�(��&E~ez(b��p�lL	����YI����׺����Ś+����0ޑ��7ԩ���a���7�����ǟ�,$r:�_H&��Y��P%���xA����Dݿ�;�C(��sr�ihP����L&�q�ј�Q³�A�;UA��,��p�ɗȆ`�U&�+��iqDy�\8fC��J�;M%�����Q>����գ�g1x�v�O��I�p� 6���榬�3���ߥ�q�ɞ�A�%�oH���u=b�#�N���(�s��p���Q���0l!�1ߠ���.!���]NG
����+�E�`Gcya���HS�ψR�{k����yMn��s��OAh�;߾�\�/�,QT����|`��ϱN�b�Ԕ;��e��W>�(]N?/p3��J-���{�^Ǫ7+��`��3�3�MzQ�͜� �C�4k��$_��MAu��js3N6������'^�`_�N�"[8������~)�k�C��YR?~AZC�0�Df8m�2� �=�O��{�(��(#�g�QB�NI՞+�jtƩ"g�ٗͫ�V.��|,�F��^�)��̏n��h8���]�N"ːK#.ޑ��v�?��WR�T!wZa�D���C[�F�n��������O��b�-�,5���[�/O�ę�G�6�/\"Y�rF}x�&�ge�����/��1Z{��-r����1n��X�FnV7�U~l�_�F2�_d�Ǝ�:��aG��/������-v%ã��AӀ�=p� �d����&!l�0����j;�\~Ψ�|b�����9�4Q �����s��Ot�QtF�N|����X�n�A�gm��z�:��tƌ͌�e��k15���$[w`�/������ʃ9�f�$�ѯU��<h(o�@��w�,�c1OJ���#B"}L�T�&�E)�q�*�h-b���T���Q��Dtzw"�+,	���F��6��प�%����n��P|)�N�:��2����tY�4�"߳WL
sY���֞o�ms��'��A�w��Z��e2M������!�W��ҩ��o��1n'~�P'�܇�.+�K
���䮗#�>&����5w .8rz�M���m5�)`1S�u�?���/-b�+n�7)�Of5Ci��D�<�{��鳮�LiI�W~�o��@ll(
L��e�'���:c1-$�tղX��ܗ������p--+sKU~f<�d)׺�7\��y{ֳ$0>���8��ӹ��=����Z+Si\Fn�14{�街G������Y���h�y�?C���U L[���Z}wǪY�������v!Ъx����FY=~]��~����蚷>b�e���hw���g���՝tv�]d��n�-{\�^�h�	^�!/\c�ONZѮ#"����1��fI�G���6v�������Qz����i)�,�5:����l/������i���+�=p֕��T���U�d|��|"���܃༙�'�Ѥ������a���XArK6Ay���J����R�KDjV������J�zJ��K��u�m���:a���x�N{����0�
|t�"����k�e�O��^����cū��`��{���k�|�}�o}�8�yp����.f�{�O��y���v�����7T� ��@?�w���=�j�E��.ϡCk=6!�AU�MY��A�j~�=q�<%emHKVU��Ig������#�X{i�+��J�b��ƮB�j��SАr��/��-�������	V\�@�c�����u��?��~�ӸT�0:�a\M^�ʥ��#8��es��H�݃jsfb�|PZ~��2C�t�[�MqPE2"����l߶0j��G~}�%�`t�xY�$JkT1��u&[�A<�D��@�$���[(f�oF�=��*Mo_�rm
�Єϼ[Ln��7�i�A|$v z/������FId8���-w-���k>�;�l�w�?�����J��&e�,��&��_Ԇ*��$4M+;�ք(�)-ܺ��D�ù�[ZS ?4�E �S���d�|�g�N�d4��