��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���:����~׳�jB%����|�nmsK�����v�ϸ�m`�p"���O(�)��������X;|Bf:N<����Q�����qI�9I�>�������Q���~l��e����u����h�y��_Id7#K( �N�PXD��݁���^E��m�e��������z���GjEI`�4#�Bܼ�-[wT�)�?a��~�'��.;�=J=Q�P
�����	�����s8��F�'�Ķp|8)�H�^[� )����������������)ᤰM�b�w�v7�+�>p�����z�⽡���<̕�?o3�s7����cUÚ6��YɫpW���um�<(����#�Α6��{���A����+�d���LO�嗬-��ᒒT���,�d��9���D'�"z汲�q������5mx򔫭���pNC���ʅ�-�r�剗J)YW<M�����j@��ȇ#�K���%��F���^q���s> ���T�VQ�t�ɦ�M������q)���������gT�%����m��5}� ����׺�q�`���,�(�:VF�_Ʒ;vP�Qb`O���XpVR �-�5 O�Mj��9 L&s��`}��w����`�8�"p�V�_V�F��yYb�����O�`Z\V�/{��F�1�Z���m`2���`�P�wh8�v!t�Ѯ~� �S������(p��'W.�!����p��;m<����@�s4"�)�I7+�Ґ����;;f���$��ƭY��b���N�%��V��.�\��թC����<�9}����f|��1�=ӇIw��ٟX��jGw�O����aɤ����fՓ�L�"�\�$��S�'f������ S��a����}��]�3i��)���ݣ��:d�*
�љ��|���.,3���p|��z��p4->TX�Gƻ�۔;�ĝ��X�R$-(�W�\����P'�O\=���u������d9|Ԙ��s�|�<�3TyL�6o�4���SDfeTȑ�_�-=�p������?��y5)�����!�0��X��\\�o��/ʱ��w�"��˶�!��b�Ci7ZU�AЌ'�:�ΰ����aAZ��c�.?��5#�_����,��D��6v�5OY1T��`Pu,%� ?�2x���f��F>Ǽ�;�W�vgU�@����o�R݅�Mz� �@����%ݜF\�jr�'�#^���|���~�P�!Wt��h�v��2��n�[C�#�����Z swF�G��n��C��8�Ӹ+�8]�6qP��%;�
^�YM���.�8}�	���j�&�l�8�'�[:ٚ2 ��&fg�7��y7C~L�&X2r�q�%Ӣ	Ob�w^=Y���Qp^��W����o?Eŷ�NXci��N��&�G�iv����t��w�3�/-F���O�M��P�1qp��r�8�k�	�Ɣ9����P4b�k���&�"I�Q_Ai7��I���Z.sd��`ζ�۸��)\��B�ͫ�c�ta͖aR� x&CbU5���"=�u�j�������L�Y�H�>X4Y0�[j�]8����{�m�&����cgd����*��Q����%�j��XM�-|-���8~9�����a��P�Z�++Aj�f����Mؙb��MIL�e��D8�.q�ֺ�[�S��g�m����[�k��7t�s(��]1T��l�{�y�Հ;�݅?���q�y���j	R�/�Q4�(a��t�	m�Ύ�
��쏈}.�XB��񓋖��{�	�w����:a��Z������d]2:�=:3S��X�H����W�Tȓ���\J�b�(�XOM��4��qқ/�DX�S{�&�&�@�S��"��ٯ��N����~��ڒ7=Հ���l��˪��X�F3R��s^�X��HLj��i9�Y��
�1j��6��D�x9����\G����s�>��:�#��/nm�v*�;�7/�k8�:B�j�;��I""�ZW�s�"�F����҆�× �����+�)�!dCE� �n�oM]0��_��[v"�B6�m���&��EK���4f�ؽ(k�S	��0Ō����p�����ƣ
���5js���M���)˹��3��|;��	�Ti�g�X-�7�v�ĵ^�Q�c$8�>*�&���G�p�EI� �1+/w�y�|,�����׮�R�C+�z�a�	،��ʟ���B�:�����0v�6��K�ŞӃ5*Q��]��?��g0���_;8w���W���#Ώ5��@��u�8�{6م7��	�1�,t�R��@QU��I��n�d��sUa!h�R=�Sc��+�~�~�3�lI�.{��#t�)�*����/���u���?���$��Z7��Ir����cC�>��ZU*���5��7M����ϊPM�{��[�
�&�(T`�z�����AQs��ii�=������i(f����3���a�Y�!�*j�^�4�k60��n�Ͱ�{��K>����^C����tW⦓��� ��7��l��H�K_V�?bq�|����C�����,X���2�3�J��9b�.�i��ӱ������!��R߁�5�=���I N�x9ԉ��4y�s7��Ő=��gr���ӐeCc��(�ZT2�c��'w'�H��3�,� D��X��q7��3��m�楷w��FK?���4�ی������iڤ,���A{ b�h��ZFK�ٚn��1��
ܼF����F$��s�)�E�F���5�4OdS~�0�(�o����y$��I��>i�צ��כ�.�������lM�>W�Pk�~�̦�='P���f_K�~��ݩ�4k7��ڑ�q��[�0t��T��q`5H1�� ?��QoP��l1����ב��S}�c���;
P�cWt^d��t��4��eª�
�lj�!{��~q5�X�Ŝ�jP���y�3�aGY����6�->��t��������;�������j<P*ӄ_0���la�R�������� KÓ��v׋��wUx%9�Z���e�pK�n��݆�5�2�1F���c�����sE���&+#b�.R�#9V_`�T��b��׋��䂛EH��K�s6K�=���0`SM�'
%f3��4E�y�EQ�g�t`wNG�U��~��N~�K��F�K|R�*ΞU���<�����al��+�&���=A�b�Z������d�z�h,"��#�s(g,+��^)�8
����.�%_*|E=;�{� $%L����O���L������*
��Ñ��+B�{1��o@��� $�WW�3-����ݧxd����8Mv��ZĒ�����O�d���-`������w�!��Q�Ŗ\�Q��7���^��yr�\�C��i�y��"�K���q�m����+4a7l�6��n��%���K@�]��"�n��e����Ne ز�u��&��Ͻ1Ub`[�Ws	Ɋ�&������B֮��VQ祿��ZpY/�"[�>p�)U��RS�e>����@��_?�н�fyVr�g��-F;��3�bm���n͙�D@�W�v�S]�TЏ�&
��5ă���:N��R�w��i�|����Q޼x���%F�|ŕ>]�9��#6E0�~j�cv՛��P�]�^��C�6��EO�~��Hyu���J���Zp�2#Gg����sO�ۤE!f$2�2�����Ӵ��<Ʈқ��Q�p��������R{�O�2  ��v&������!8]��
��9o�����7��웒jߗ���2���L�g��h8��,�`�a� �&��f������[��0���۪���I<��ʪ3/x�$։l76�fS�:B��곮σSQ�wB�/�#� ����DȢq��ݙ:l��ʔ�f��&������l�/u��l��2#�8 =L.��X�9:�g�4V�U��+�幑/�&�)��LT�lWE��1>t�@@�'l΃F�M�x.��ZZ�$ӄ��c�+,ڠ+�$N� ��sik%��<�^���r9�tzc
���wFS@A)��n5�C�%bx�g�OC_VS�"֨�}fZ����S9�7��EC��k���9�\�ٞC���hO.����G��\������9��"�{Q���Oiv�����vĚD3�L���Ƿ�ǐ �/�	���v�I�q��乊�h�'f{-4�����&�+2���g�[�Z�3��W���:�!��ʖ����x�:�Ӿ��(ԍ���G�jFT�D�����zί�Ml�����X� �[�IYV*� ���3��v'e�0�ٖX�TBle��w SH���]���f!��(p�!u�����@�A@�+2W�R�tyA�%o�/�5E��3Z��y���iŪ���[s������p���3Q�RT���60��W���t��ѰqS����Zc��l��o̤��-S݈�B�+<	W�pĴ,�y�ī�889c?��Y_@����P�T���
�h��x�߂)�%�U�����F�]��uzq��05�T���p�lU��عq���0������E��M��~@��g`2`|���j ��D����)�q�xZE�PQ�J(���]�7�}�8~E���/哦|}�-m�W�}Wu�����j_r}����4�amQ�ДO��$͈{��)@d�0rC9�"�?r�);�����*�+,���~�����D�`S|����;���/�΅<�^v^�)fw��(�>��J%[��UNP�
�F�s=��w�'^�5U�����&��6z������&�/���rם�g��i� #Il�����������7{�����__h��u�J�u���G��
�g�NK�0Y�}Gu��h�\���-zm���g|Gh�$�<��0�5� vo ��<A�)������^�մ��/a�L�0op#6IEfJ�ŋ9�#��'6���!<�I��20k��k%g��=_$��BC��jh��X������cK\ ��qu���?�3k?�H6�h{�Ǌ�n2I���g���ފ���e��r�Wy������4"��C^�c$�����H���� a��j`Ƒ�� �F0����(&S90���Odo	3���(�b1x�]�|�ߌH<���"C��y�����a_w����|�`���a�&�4׃��Y��U� ��\=���|�#�z��&�h*S�$n�f����H0C8�k�O�E�Jv�8mw��i��:�v�iiG���o)�w���t�#�Rː��(#[�!�n���N^wEg.�%:Q|�k�H��_Oj8���f�A(۩(��r��2t��!K(�0-����`��H�&��z�=?�_�y8�Z�	i��<���iv�O8_�l+�+�j�YG'M�T��Fg��N�4p�0K���2M�=���$Ce���feiu�S�C����,���!b����ѰP�M�%�k+���jd�<̄��W����X��Aja����Q��A"�y �'9,��D��Q��ҙ�9��:� �R͒��4!=�N :C�׹a&�Em�0�Gy��[(,�O"��c�)Z�Y	e68U�|��L����qr�kQ,�j29��$y	r�?�G1�M8�{\i��~�'��7'wϯ����P���Fo*�kV�5��ۑ{5Ş<yH���<��.J.:"�s.��-��KVj�+7o���~4^`�����ED�cY`���C�@@qaJ���+�EА֖֑@���R��l������_4��*�pk��Fp�u��a���4{�I�m���"�4��;WDgW��y�@N���}�8Y�E0�v���5Mr��/��r�s�]M���kG����?�ˠ<���"v�������P���s�B�� �0�՛��-qr�+���q��cS�m�U\��H�Qf�'��L�D�m͓�i�����)�RB�O0�P�ff�&����0l`�们��͛$�p-��U������km�]݃�?�k��=�/رf�w�h�
+5k��9S�����S�*�}4ktG�#[�i+]�����}OI�I[(|�Z���kSij*#_$Ƒ�0?QXD�m@ȳ�!sie�)�"��C
�X.�:�-�7���C�L��w��|!߷�i ����e9��R��n�D/��I_6��C.��j|���͵�]������םB3�������:\f�>wՇ��+�8�Q����z^xv΃�˸(2����5�!r�Y�r�[8��?\rG�.��w��1��ZZ��O++�#���నB�b��f¡2=mt;�"��nY�+�9ܲ���]����6��A��rL�p��{��εB܇���W���_���[��vB��o"9�`�P6FbPJ�C���Ǘ�V�7=��^l�ve<�����!l�d�AN�-�������d�E3�8���*��;|�L�U�j��;v�`� ��`?W�R��9���g!|Q�Eq.!�+�
6�'7��Nr��$dFE�*ϹY�0;M�
�n� �?�s�����j訳���d7.;����U��X����_�xAh���+�����Y��r�Ċ��-�6����0}��.C-�R2|u
*��v۸G��ѹ���1���Z�p�͘j�P�1c�\M}��+
�|`=�%�vX����ճ�Q�.���a?�j��D7��H���&�>˜�*���Т�w�&���39|�YCO~�@u!���w� ���R�b�Z�s�(`�d�=��o��4�ǜ��ja��xL�fǫ�����<Թ<��W*��3q]T0�K#�R�̈x�[�c�_���S$�.��ur���!�W�����}�x�F!����7�KȳYhyM�ff�_Hm��2���F�)+�[�AP��� �k�f��������ܾ�NS#��٧՜O�?��#[�$vt�^����w��u3�J�?9�Kn�-������q#�vA(�"��}b�:�������*��"�%?%y;E��"\;�vUK�A��.�)�6W���3����t3��5q�a2�h��%�v����
;��e��N%�Z��bu��-s;�p�w]s#�d�*���ag����cb�f�B���Uϙ=�Oǫ��H��O�4և¥���$�����S��~R�UAʧshk��C�~�t�
8$�Јu! �T�X%?tēB�'5����SKr��V	-�����X��Ų�tH[z2ͨ��6^כ��ܟ�����yX+�S;�.�m+��gE����}䪍��R��uAf~����]G�(�࡭��`Ij8��'j���
Aoxs�ز^���tߖ�gw�B<O\�8Zv��ڹ~��o!��ciWh�8�d�+;.Q%O�w�[S*+��0�)9���J~4M1�c�r�N�$��S�C"�j�h��۷���P�`��f�����N���*?C���K�K���'�]���T��A١��� q��RR¾��Q�9�ܖYm��௷v`���4F.��RaGy]N��,��Q�'YAf�!<)��J�Dl����cP�'\�$-n���4&�>ʒ��Fm�>��]�׮�r��FR/ď)z����#�'���K�Fފ�_�Ǟ�M=;l��sv���	�|B�ǫo�dsp_���4��'�L������С1�]�r������4I*��ӳ�~*4��BH*�鲳��Ы�[�T5>7
��c��t����^Գ/V��4�m��'>]w����Q�d��'b$;"JH�i �zZ? _�Z7b���\��[a���g ����STyߍe6�G��RT��qژ�*2JJ�oo���B������I+:��e��agM�	�d�;��A��}D<h�S�
�&��[��R�F?��`֢C�����=��8r�K�G�(�i�N��^�jM�v��$bܒ�E��vy=�ǹd������-����s	������c�*i��.�Σ������~����r˟�8+�l�/�e��7��O|r���F�b%��h`A���-u5�N��p:vLH���
-����f�������'lf��C�hq��wNJ���M�hW�>��q՗�;0P� t�SF~���P���R>�bS{����q/���Gf�Ƭ#�����!�0�\�(ň��@(t��$��S�#<�fd�gn���n%��F�֨T��`u�3���A>;N��@�������z'��=�W�5ڄ��M�����������JZ>�	%�����:����G>�� ��n8��0�Ł��Z;�#"�O�IV|@ӫ[�f�eq�hJc0@��QO�WJk?A��`s
ż��` �{�+K�ʾ&w���|TF86e$����]eX�M2�y �w|��N}�J�5�}m;��?+%�J�w~7`��~��sQ�ͱ�[a�-��Ho��v��X��U�786��\Z�GOB�K_\+PC�l3���	�3y)���Q����x�y��f���B7|]z&�P͒���]EWQ�Vױ32��4L��CrA$�W����D�`�d[�.�ϋq����ѿ��?S�8� a�A�]�jz	b:��І#i~�s1:$��:�����jx0�g�4dM�2��0m��w�{��Ԙm*����_�m �2~��:xԳr8@%վ:8���3R��YV�)�(��F�7�*��1�b�{���^+�:����S̸㫁��VVx���|�9e[���,,
3��k�:`�z��Iu�஦z^_EU�ْV����ǜ7�Ȏ�h��95��ɇ�`E'Lv�F��z�.�ͱ�`�r�a]Y+j��(\�ZZL]t����R��	��e6�u����	;�\Wg 	*K�b�9�i
:�����S�������"�([=�toz4���x>m�e,@*��6�I������������V�$��w*�y{�5�\?�mR�����hqE��J�$���#DY���}H~���C���j%ِ�������zՀ;���[li��s�$�C=  d"��[��y�_�7SMF��C����J�X���4��'�q}��[�E��[�7E��'�w�\�w��"mf ��ƞ������ͬ�ƭ�c5��s����\�kPץ}:B�Ҷ�+�MT�Ժ�:��@�B��E��[�v�_@��G1B�sn�;L@���GtBw[��:g�F�/������ӜǮf|C$i��$�F�A�Gb|�^�j��Jh&Z,����7���8η�^�e�E�ٖjjU�
��`fL�����$�*_��H�<�ex'�A��t�9�i�o�U���l���=�U�@�������v��!�:{�'
L����Nr���v���D��wo}&9Rh�5�&ע�|RP$���ٱ\n��(!��˪�L�q��2�gFۀ!Y�sA�$7���S��k�۵�<]i���m� .�4٣VnKE��vzϦ;h�Sb���9��|�2���ߔ� ���'?�]��1g:F�׫���M�&鉬*5�v�G{c\[΄�l�P!��o�K���|�3�=)?c�#���{Z؈���Z�L�L�'�P?	)��*E�����!��w��߂�G�p���q�I�W%L��NA�4q!�`��4Ʀ#��2���|sLq��O	�sV��<A:�cF�j�V���B�f�죁0�c/n@p?�9`^��?��T� �F��?�;y}�tL�7�,��T����,�V�����`�\3R�X��U}�\�����O�Q���l�C�A���kV1+=�8�c&��-�\��
�����D�#�OO`����j��q�I��,1��D�Mo���8�Z���&Q�<L�v���-�/ɛ���o�(��:��_��*�A�����'�A`�2(P�7U�ی�j��n�J���a��o����[e����a��S|K��٥<��˿*�a��7��J�����`f��Y&s�;��<�R'8�L�F��[��
�A�{���1��R��ˈ��G�h��ԋr(-m�210�Re��Ԫy�	'�H�Ƣ}���i�H�Dp�:U�kah���7dǤ�UW5U;��I-����N]F�=Lݱ.)V/��E#���i�g����,�+'[���;�`|䟹Eq/Q���$�B��Zi�H��{��<Ѭyٚd�'I|���a�_�f��#�;��϶�݄�U��
@�a��𬐾���+wW�&�o�)В���b=Pz�g�8�9�Ja(�ߤA-�$�m���%o��q�fsԇ���9���'R�L��p�_�N���	�[q� ���0>N�{��kZ��X�kד $Do��f$خ\��>E��Sp�Z{�)��8�h/}�ז�m�'q�|e,:]⌳��Q��^�U�-a�����en��mu���}c��X�IP�)�I�b� Gs~���9O(�+����n�<ݲ`%��)	���-��
f�l�=a)F�` 	�6��a������C�g��QBhl*�
��I�e-(ou���[��y����G�z�V�G{���$�:5�����B�(��p�v�eH�X� ��J;��<T^�h�����g!�R��ۏ��|6���lv�c:y
�v����I���x����� ���3��;��6��;yI�,)�f�X���ix<���o �S��R��+��HNcH���w_)����=�*��O��ѝ
Ւ��p����_�
f�}n3z�ǽ�^%^"�#�f�p�	����34�=ǡ�o P��Vt�ؔ�x������'j�t#�˄�˹��Z��W&�Q�&��Ʒ��߯���������S�͡i0����62KX֪����hŚ�:�si� .������Q���5�%K (�>oIOl=�*����� ��?��V�'zr�h�.�<dm2`^�iza�#���v+恡P�F�} ������S��͝��R	UǓ/�3��)�람x��k�Z�	jw�a�P�6�ṫ7�J��U���{��(�>b��Åd։v����Q���n�K���DjG������N?Vf$k��e%6+^<:^Qd��X�P�}�1�����:��5j���@m�t�yg@_?Ё܃f�����{����Lh�)M��Fl&P~�#?<���`���Y�|��"Jlc�ڪp���Fy]�����j��o)ϣ�f�x��3n���%3�>���#�
��i;�R�t�AG���>���Kͮ�������f�dJ�3����`J���wU�t!D�f���x[@��h8[�h��`Fcf*�����_��_�Kʎ_"}�=_����[3���-?}$��D{��%�ճ���yHG�{��r}�ݝ����M7$&��$���VS�M��1�t�%��e^�t��ݱL4 x��+1��+��_�$I����D:��#)���T������;�j�J�EOɄ'_d����kl9=�MK�맾#��ox�����<Yj �+��A���s/�a;eLݘ�3GMae��9S !*Ig�=���ӞL��j��ח��F���W#V�Kz�Dc�K�C�!�<�V|�Ao���`�`x�� ���%x�@�X����vk赾I��(��d�#�`h�)��>1νno�_Y$��1�í�\�2�qĠ��4Z�wWM�����c��Z�o״uI[>~@F#Q�JU.����Ri�ئJ�y����0��BT')p"�)λ�	��L/��T,D.�D�jcUm�O	��2��΃5���#����B]m��
UF/	v/D�H�++�j}*
��iY|`�c�~���A!{v5ނ������7�V�H�5�d�V��_��{BC�ۂ	�^�����o� ��*����`�#��E~D�/p�s��Zn���Ͷ*�5���NMeKd�sǹЩ�&�I��O:�
������
v#,�C��9���_�饃<��\@Q�7aS��P��*g'�g���q8�#�s
N�Hǯ��Ŀ�@��ʐ��=������3t��Z�\�� >���c;�NP���qHf�S�%nA�z4�x���b�Ez��Se9��Fl��6FW��`��5�����oM�%�5c\�x�q�A��BT�kc��1�������/�E�d�V�����^:o�F�DX:��쐰h���'o�l�=l�K\����s�#�k����*J<X�b<���J�"1����b|��[u��|����^[w�Q��5�|:P�ts]X�Z�Vp_��m'���FM̧�`R��S0`�:�آ�����<�{u/�v-��"�]����������)lCP����7M
c�.S����EY�����t~����=$��*p��D�m
�==~"�`%C����p�R.k�����"��0~���h��k� ut"�W���9Ks��Y\�P�=&ZX����v�?�9�Y�\��I� j>�_ʪ�J������s���(r�R��q��.��"����+�V9:,�M\�V���#cb��
ֻ��3ЬD��Q�yB��G%7��6Qҏ�4�Qu�a4������:Jz/u`���ֈd�4soV�p�_ӈ|��V��6H(N�
"Qe[�gB(���H�'����K���+�����)˱n��;2�
�qX�����L��[��,��c�ImȀr���+�G�'�:�����~:/��� �Q��,Y�+*ޢ ����IA1��c����X0� ��K�mK�Y;����H��g{���n^S���Ġ��1���dt�����_
>)��xĔ/B���F�we��ΰ��q�ۛu�B�\�r\��>�9���[p�G׊I��l��m��%�d�Sy�h? u �;?64��K���(����sq��cࡒ�I��-�G3�_�?+�ޗ-mV��f��yp�l��P����oW��~����%�}�2����Fu!b`��d�F'�\̾/aqY�\�P��t�vS�/���2{���b7�q�f]���"���(�r ߇�G�KI�D�X�!�F}#�����(�h��P��������q%vs�P�/�L࿩�K��s@�0�sT��W�]YS��qN 5�i�[n2z�j;�� �zd����Y��<���c2ir�n�1e�
���7a�5���P>�<- ��&P��U(fs�5P��ŭ���v',�'"�J�xM��(6���%6$66��0���q��1���-xΎ����F�������[%`fE"
3`��h�q���*H0���l���?F�%�$���+G�d�S��M�dtS�y��<�-�8�������wO?�ś'�P�SSC�
!į�Źj�4�).���̫h����Id�#0CMy4��#ܛ�� ��8���Z���pLbv�ʊ�Pb+in���x{h�K�}���xI�?N��_/BX30�4�VA9kw�9F���e@I&y>	9W�p����B,`W�^=v/��Q׀���]O�	gȌ0��!��l�#҂b��Ӈ:��1��E�h�/I��5�gm-���:�y�໯���K�?Z�҄��S�C���>�\ܴo�{�_0�<�'�X�@�.��v�s�,MgE���Rd6��{��zIj:nQh�����]����}�n`FǾ�ǋCCKª�I���O{�x��L_]�GHF�����eU�H�X�"K��=ȕ̜C,�Ka�}�]�C�t��K��M�Q�3��Ǵ���Y+}:'�j�	��Rh�juȼ���'�5Ğ��`Ρr�f4Fj�X�b��c��qGn�-Y��úC��'Qz��lĨ�eqn�����>S���n��8"L;5jd�����s�Y��o�֟}r���� j<	y���͑J����i�`@nd����h�v�x[��<0f��F�j�&�!��D$V�PN��9ƒ��wO�i�B���K政�ؤ(6�U����m?�?�y|-�m�vN���.��j�<���P�0�d.�x�0x�IZ�B�7$��Y�D�������1��W"C&�N��?�_�k�|5��tp/��q �2�Ǐ���~}2���7����{�EQ��q�|��1R�H��K_3���j��(%�]m�jOٴ*S=&&&���ނK��5���b����j��X0��N�ܡ��8����j��=s lhC�71S4&�ݗj��ݕ4��WPpڜFjn&oTG7�*���j�,A�k��Z|�"B����G+�񪓅��BT���-��[aK|��μ#�(Тt�z��M\G��!��l̫~�o_�ƾl�9Ԭ��tŰ��R��������s߯J����)m�%;�TH��s�����I)��˗�靻�#b�x�j�`��d+a��Fĉ((_�䱧��oK�GM}����l�wk���K`R	~�9�����x��.��U����\v�� ܛ��v��@;�?	�`O� �|pC􋔟�UD�!��yj�C`�"�����m�m��\.�r" �Ԫ�׊Ͳ1�)�����I*m��6(r�a��L�8�E�L��\�
���a�^�I�`a���UZ_[�t��w����}^6�E�����?|٧���/O��m�����H���Fx(.L="���ktU�P�Wғ���"�����}~�q��c����5ի�i���rcP��Akg���x��٬�1B����s��4O9�j��@_{�9x�j�5����,`h��N�ˡ����g��W
��
f�kX����dd�h���y��5�p�Iw�|�gX]Rv�
k�?n�y���I		
4��ֆ�z��f�g�:]A�0E���I��Ў誽k��v+w���ܜ7[��sUת	ٸf�bd�<� ̡"��xf�+⷇{�.��杛�U�zpDQ�U)_���I�Z����kj1�Gd&��j[
�]�K����'rK��`ng��3!:U��)�PΒ�y�#�̟HV�9?��h�����l@��D�5~R�X��&�@꾋��Hl`��|�;�="}9�h��^��x�H 6�)ɗ��?�~= �0oF; v������\�J
&�^�S~-�_���`�V�!�E�=T.3Q�FhN^�@s��w�\��*����U�>�{ڤɇ���S�{8:i�$���J�夤�|C��15I��&��\��42�3�n;1Sg��IY&�Aʑ�}�$UG��U�X1�=5��3��g^za,�/�T�͝@�@���tx���2�dl4����P@i]OP�|��n��r_� �i��\��u���>���C@doc�%&��{fq����p��}Cv�6�l{ 9S���a]�v?շ�ת����Z^��@=�y�$���Ɂ�3�*������P�2�i��oD{p"�Tn����R�fO١�f>�}�\��_t�g��5���ZHv_�t�'I���!u�J����7��K�
o/
�Th����*Ȁ�d<�� ���S���G#�{um�p^A��uL
Ѡ.e���	/�p�qS|��|f4K���\s�p?���b�2��xC&66QV��j���ŉ�0�K����ɛ2v@w���)R�6���}�^7m���L���J���߫�����49�@���^{��:D�'K�	?e�U��+0����	��My�Ä�b���>�����`)7��N�:�(ja�̎ ,Z�w��I/�n�@?��
y(���W}ē��\+��<}�t���3ۯtO�3c���E}船�mwJ�ڧrB�����5�w�c��|A�r9�����q��8I��ȣ�B�V��H:H�⼳1�n/����J����?]�^Tb|Tf���fN�G�9��.e]�Rw�X���9�Z�T�#�|6y�j�{Q�?�Ͼ`w���ߕy0�k��>F���IڝٙYb�"�k�k�g�rgtFр����h�km���[i�ogo]�R�,b���+�URթ�D�~X�R�	>��i#���@	�	Ù]�%�sK����I3;3烲IM����)Ps�q�p��_X�euE>s�š��ڱT�É�Ϫ1hd�ȯ
;����ɭ�4��E����NP���)/Ӣ]��H��E�:����[1�Z��j�&�uO�ܸ��������F�Ӵ��Bq�v���0�ȉ�O��üͶ���r������r���Ɏ���!o9��u�:C�z�Gi��1�	��>�}�W��4���E"l'#2��1�#
 �	���̝*aڏn�H����SŻ��1��\gU�v4򪷍����
\�F!`�|��G9�*��i���>(�@~}>�=!�Ӛ�}�'���z/Z�Y��%`��p��5�MĚ��B�vp��~��5�x�����Gx�E�C�x���w/�������@��,qٿ
�aq�M��s;Ű��Qxq��MJ�K��eu�+����k~~k�W}rS6�n�$�aP���"Ύ��O)���Z_/�V��`�k���*����pٙ���D�M^l�N����da�D�啸�*��c�~~��e��H?�b�I��e�il�,
��=[��7N��E�M�sD+�����Y@��&e��ZKV7&�J�g�9��R#'{��V�3�/�-E�#}�R�B�GuM�a{J������p�u�J�ԑ���j��y�m�x����S�",��[4��g��"��iNx���2N�tg�SatA$x=>�tcٖ(�
�tZ��	�o�F�W�oǖ�MS�>
Q��G�~ 9��3t�˪C|NO ����],�r��U�6���e��4��@¾�j���m"���/IE��G_��\��="a��V�)1�^x�ƻ7-*�����I�nE*z�=�X�w�Ϟ�fT��}H��;��^\(b��|՜�I)O�����s�K�p\�Y�h���v0�m��gr�c^�ϸ���p��:T��z��Y��'�G$�w4�����������9����5@s�Uu�N�eF?���7��^�JT�3��sH;BC��o�|*@��I�{�"n�(F	�����1*᾵d`��_�����JL�HX�s�����ήXxz�T,Ň��%<����ԣ�����&�܉��H��=Cf)[���tF�q~Xo�:�ן�HA�ZTth,W\`����
E-E�b�����2S���v�k>�e��8�a8� ?�����oh	q8�bqy���f#�*���7�Z	��hf�,"y�f%�j�d�ӈck�)EP��F�V�$��Q/�;��]��2K�!t�,���vx��z�tx	M�����a��tH�����Zqj@��U&���GG���3\����^��5����"{7w.:��+������Q�����a搗����ݮ�p�?��vM"i�w���b�B�'^�
�8�E�؝_���\����o����7��O�V�d3�V�h��F�?<O��0�gjE�_!���V��j�zr�s;�o�EK�OT����x����ȥ�r�j�NÊ
���r�H%S�9�+uT�j+d��JPe�G-�(飝��d�|�xc�����j�>W^lصJ��1�s=��+���<M�:�( �,~`�]ԁ!R�c2UX�yz2gBDt5���ػ]�q��e/��<��1����l��'�?��*w�>b�y �_̆/Q2��a�l��0���?]���=Kɏ��t�����jI�&�,�I�n���}@& ϵn�).�4�H���q9�(�3���G�i����Ĩ5�R������|���A���
�e>+ޞ'��(���/�K�i�����`��U�� �ޮ�,���_�y$���}R���R�Ӣ�q(Ѿ�(��,�nB�A+���Ͽ�m�S�2��_��/����N�	�2�?Fv�5�l��;p��b}���&l-�����R!*��%ѵ�!�,m��݊�N�k
/�}�� �Y!���4��h9��m
J-G��=[����'��A�_�DC�?�U��(�Q.o�\��.��*ZN��}b��1�$��f �e�J���3�9d�������^���Y���NQq�r��*, >l�`q�f5PG����3�QOX>���Exy�p,Mq�QŊ_�P���G���Z9I���I~�tj��z����zl�jt�ٚ<�N��o�Wm�|��,��H�c��������U���梁�*Jx�7�>���F&�	\7�u��܆%%B������$��yuP�4�lx*r���ȿb����O�ŕ� d��*	6� K]^���:at�w����~��Mg�Q	Y�}u��v���t+�/fy+S�W��DL�X�L㺄���V�����ݾ=D<ȩ) �]�]����$:g�/:}�d�R֬�D�Z�iE/'<\��w#tl�[;b\}2�������w>�MQ�x��OV����] ���7�S�!?D���u�I���֠fp�����4���w@�N���.�4jπ1��w�����U.§�-�H���f�y���>�u#�������'�p�Q��gg���9*~�?����_�P
kо��H�<.z}�(ى�=eo��aE]L�u8tb����L�n�)N@��7Vʺr�!P��D�OE(SU=��D��?��Am�:��b��~ ݙ�P+����'��~�b�-�bL��T��� ���8eЄX�c�*Y�N �-QEv�
ݶ��2+	��.�CV�ʠ��e���;f�r���c���Q��S��Xݪc���s��4F2-OY��?*xm��gc�aOqqfy�^i`x�vj���K�z�:��@�"����Y�w
�zA��^gl���G��햟.O-���a�t{ʾh��ަ�N�	���!d-���dV�f������Qo��*�����0����v?�q�ɿޑt��;�K��2u��
4ID�$��k|bd;��lexw��#~����%#�i�����e��mh\#��p��ү�"��<,X�P��D�OH��Q@�kt��S;D~l�e�4�m��'>�ĜY�$W���9��7$W3>ը���q��;sTG	�wJ2���.V���2�X��\�1�Ɣ���;u�V6��F��Z���s`�����(����]�@Y�v�=o���q��\�~�����xU�A6�|/ʐ�GKZ�{���d I���UXjA�<����!�k "�z�|��$C4;z+v-����.����x2��u�l�'D�{���U�Q:��¸�'lZ������%;������<b2R��Ȉ��TR�-3�LΉ+n�Mx��=_�y���e�*7Y���@<����WI!�(ȋw�WF�f���OC��CL~��"�C��@�r���$��tn2<�+A��8� ���cJ>��Y�f�K�[dʣ�tw����RCϪ�ɑŭ�%��=���-M՘`�Jd1 �5U��-�!��Vifz q�uЬ�fA@�y#�"ӃQ��[��gI�h��z�3N)c���Ga��y���Hp�%}�Ԙʪ����o����t���P�����E�u��޷5�R Oa�d;R�U�v����V�L�,���
�y��]ڹ�� ��M�1��w���5��)A�:�����o���x�e?�E�x����+MD!G�gϩ�Vl�$$����G���4�W�I6�jV�I�<�5t�@�nK�u��u��wZ�N嚌AM���.H�t�Kԥ��k����W�b��Qk�H_E]������`�L��=�↊�3�ۨ�"�^g/g�J �0�w-�������_q��o�0��Tسל-w�`۪O�:��M��Qrޮ) ,u~O�M%�m��ݕ�>�%=9��Ḱn���,t�!' w�2���W^��-�e���N�l�	5+���<��8	��bM@7A���OLm(�*�!�gK�δ֟�l�&0x���n(=�q�Pt���~���j��6W����7m���T�Y&����Xx�~���҈�T�L2�tv4����Z��� y+O��ϥ_J�[KZ��_��<
�p���m���
`6H#j��P[��4�j�����o��pp��|�1�UK�`�:.�yt�m��^��Pܛ��qc+0��"�w���n.'���ы�b=�d�kL�h�)�yūs2u��n�8���ÒsnT�܌�o��)�r�������FJD��?�ٲ0%v�X-m/�q������3㰢.��������9�锳 �U��L��Ik�ֱ�����w�G���8�1w����{a�o�l���E���.�Uء��!�N���(���sb�gD���c��(��p ����a8�t ��F�� �ϳ���fK�r�}��w혎���������iQ<,�<����B~����*��:]!�߹�u
7�t�<G�j�������D�Y@Q%�L�:j��SӖ��(}���������ެC� �����3!�����,��[���*a�>.W�G�zO� j�ܯc\;N�nF�� ��y0iYcų�W+��^��t��f6.x����P�Wϻpm6�y+�|��7�a��\X�"��y�_�?[�S�7���?����u�N���F�b��D���#[>m�������@���ӿ���t�=���M�2i�m2A�茠�o}�����G�a����8��`�,)j5�^׳�W�V��^�Pʳ���5S5�1���!�?a�0���0�g\�_�;P#�L��w�Z���`Vn�N1z�E�T�������(��3w���o�vمil�'�h!dY���W�vp	^���óYp�J�z�*���'�87�fhT����{zwho���Gפ6�e#W*�h.^h9��G'�s@j�DT9EߢP�a!�&��:�1z�pw�;��!����<���=o{D֍�h ���0/�d5�R-�m-���<�bQ�����������\�YM� �_ݳ�v��G>6�/��<�x�P�����?��}%�h������"����L�o�D�j��}k|,l$���b�J�J9���]R���m�p�M�J�@�����z���72�k���v�O7�u�ŃS���#�(_�v�y�Lk�uW7[q��$���(G����� ��n�o��9B�_�[_oj����	�_�����曔�;�5�b����A��к�a�)�g��"���Tj6��Δ�#�V�O�z��y$�tU�@ I45D�Wt�w��O��1I]��(�C ��z׆s:&�ڮ���?-h=Hsp�ք=�n�H��i���h�Q�/���/�@����{Y���>��[�Nc�3�`��oL�*�O���[ �:����$|h&�6&*k�aj�{�1ק���t��E��9�^��"��	,�K�����f�����Ǧ���'��d#�<��т��=0��+�́K�#u6����rTd���)�Ը�|k�l�߻�Vά&s}����#�%���o������&X���Wҭ����S���-T[]e�?N���r4ƿ��_$N���#���	OD�x�Uޭ~�+eA��,�e_Ĳ����{��-,n\�B��B���]�N�y��R?pu���>!�B�q�3�5/B!@)|r �b�}h̩���{}ؐg�t�6>�d����[A&P�=)�� �un�意U����9>���9W�q���9.̳r
er
?��pYg�ef��A��yRΰ�d��6d��
7�IBH�A� F��[�>w*��  ���� �q\g����dba�.���ޏl��AK�R|�� c�O��[��j�˓9l��և%d<.>�c��+J&��&���4���ַ���I��CTY�*i=�SM��)�Ek�F�laC��֪�����[���g��}`���N�h�Y��o�c�{e����~K���ٛϊ�$[~^D&�;�[b�.j�y�Ecf~�](����1(�	_���s��G���ږah*��~��1�j�B2�/T�O�YW���i)�wr՗�t�4 5�MD����	��o#j��9�9��w?�?O��.���$��F�=O �15�f��cH��1�&$B� �H���L�܍��3�و�fٕ*�>x���n~M���t�Û°+��3�8��(n�1���l���y'����fư2��ʙ_D�W&�!���z��;.��c�G�"^�˩�܌
T������X3*����(��I��{� �ـ�o��s�
��yD�\�Jώ��n}����	�/5��x5��~��~/������)v����H��Ht���p,C�9��T�E�H���Y������@385l���+<��}��Bn�zҎA�=�/ز~�`���g��*~&���ޣ�w��ȩ`�ґ�A�e��f1�W�|�!OK���ϣ�F����.�,�|�<��HvV8x>��' ƿ��w�����]�6� ��<��*<��f�a�:�3b}���p���WU+[��'��"��LI+��ց���x��hm��W����p�g?K��)8S�a.x�}���ʳ��xWt�hw�0�\�r?	`:=�������o8�X	Q�9$7��C�cAy�][P�T��ၠ�1<�lT�J����O%,\��s�)p
�+=ЌH�or�f�;��)*�Owei���N
-�����F�_*��W�����9=,�2��\i�~zth��>y�u������O-�HX���~��4�)�_#�?�¡-JD�������%&�J�d�3Cӌ	��Zu���_���*x��
f݉l��S�qU�5��	�z���"s��(��x솵�i[�.;p,�i>�m�bY��4�������%5:����g �JY4��B���y�x��`�e���д���G$��/EO��\ڹV����ڊg�K#/>FoF��g;���H:s>��禺R�x<ؘ�T3��j��211@6� tc�805x;�i�w������cɞ�"#gs�FbOu�?oa䗑��e!,7�Y�����*��=8�p'@W� ���+�8K�G)�:�ʫy�

�ŦZ��;y�h
���[��	 ����ò��-�I��u��
2�����K%ڻ�}M���Cz���K�����iu�/+CSӭ9�TK�� x;�c��+l��?~05I�}��:^�IHV+��=�k:Ўw#2�;?ԦeW�U~$����� #�C������E�r�۶uR��*��(�YO��)&0#}
�~wz ����I^N!�3�M�A����R8}s߈�mϪe�&�z���D�67������/5uja���{MU��r�c��s;�ʏ!}�����V�-�U2�)7o�\zʒ��Sb�Xt�_I:�� ��F"�������f}�2��`˽�Ev�=�$^C%��s�EsE?�d`��W��/�E����rAk��?*@e�F��d�U[�v�3��^y�i�N�'s�K�z>OV�uS�lu�^�4�RRi/k,�M�A��l%�����	�a��x�P�Q
K��bN�g@R�{p���>[LY�N;�zM|�*!�)��\Ι�����A|��S`����*M4/��K���t�����xIS���(}�A(�ΐJ�FՏ*O��hl�?ύ��H���s�X��R�=��ќ,������<�p�8w�5�UHa��h�ۅ]�8.Ch�)e������\�ͺ{������OL�޵���ީ�~��ȹ@d�Iߞ	��Dwy�V�&9G��O�t��b.=-��$I!�6>~cp��G��6��;���O�=~�G1�"Sj�Y ������K��U����d���9��@ߎH��������)��b���4�����d7�/� �M��B���n�J��S|��-�k>yfb0/6=���\��w��^�P���e�d;�� �����j��r�������vLFF�iP~��,��M�n��Մ�)y,Z�RQC�J(o5�����u�q�+Hy�����>���H��/|_����݇�dm�lqh���V��W?T�~R��@h��	�Z�ΰ��0w�}	����5�$Ĉ�k���|q��ѵ�"�h�<������>���̤�����]��y�����j��g���$�3�C�8-����͍�Q\�e���c<���Ը��c�a��6��?'ߔS\�
/L���k�+��n�-�P�W�K��g����^>�q���=��d\}x=xC�'�+��22�"as�B�T.���O#��t���,����1��������%d�U���^�ᮩ���u���O��	��6v	�dn��4"���8�;t`�ܡ�!�NG�Ax���qp��2���Q��VJMޡL����E��@Mڇگ�ֆ�BWM���c0=4W%�<\����O��$���!l�|����ĔVi/�cd�ng��8��q�J(J,�*Z�o�n%J�Js�v�P��}F�=��+��0H0$�6cJ5S�)�bZ�d$�~x�K�F�46霩�T������p��`��{r߂f���]�_�Oۏ&�<CP��#C��<* ##������|1�:V�[� �3����C���wͱ2��g5�4/.��D��ﯲ#˻�2����Bkњ��}
B�yY����#�}^�e44�w%p�S[��8`Ve�4G��vEw�B�5	��_&>�C�$/~w.�����X��+������(P�]� b�tvwh�|
֓|"u���o��0��	�li�g.�w[K����4<=�g��"mZ����6|m�=S����l������yk�J�b%A�p�r��q|�,	�$r��a@������V,'se	��+��E*KɊ�r�Eh@�Տ�$_�������^��&�xg11�EC;�w��=&=x��?�֬]�cBC{5�<�iY���N�6�>ؓ0��#����V�{d�+��C��C��+�T����Hh8%�(bN%@r$?mG��ˣao�K�nԕJ�m�~.�ϓþ����W�Tn�,\��"�e�ǅ�\L(#u�>�7- ���0'��Wj�$��2�U�F������0A=� s����p"�ƃD���th�'���-����A�������,�"鷘�x[����z����*PSBk���ŀ"��~�&��!ѣ4�� ����B�A_�Y2��:�z���fqlk�E��_(�HPO���r�j
#h���jXȖ_w�M��SI��8Q8(p6�\�ӳ,\d�kk��w�n��Ȁ�`�p)�w*�T\�$�f��=� +D��,�uB]�cC���R��-�Z�e�i�d��/��t=+ [��Ǟ���Ƚ�ӵ��wr�b���~�	�$]�j�]�j�T��
3�9�8K���/۰=G�ɠ6^ ͓��َ|�]��G�#W�	���м�k���FF��� wY�Ͽ���w�nw'���T!�Ekb���=NY�4�2�+�k �32��'�A�f�;��[�c���自|��C�V�mYD�x#��n.V{$���d]F��
WV���9>�q�c�9�F?�V+Mo��j���e�p[]���gi��N:'xu�z����ϳ-���WW(P��]R���'kvZP��L�]?l��9�Q\������5���4S�ȁ`Vu6�1>ӻ�����ڛ����g�7�4˼[	�9�be {������c\�]�!��)��`T��w=����<ɐ�ؾ�7i9?�!�����Z�~y�~��άvA�����B�%|����k�T�dJ��&�5�f���U��I���Pf슇�l�1�E�WgP��H���c���Ð���g�L��~ι���*������7{+�����u�w:E�^�E?�!�S?� ��LJ�y�vc҈1e�R��p7�%z�U�����*��k�k�܍#\6���2�y�8�6�sr#���}1fu��3�����E[P�E�(��6|�	+�xa��gw4����qjJ'�~3çnC.?U��V���!/ h] lQ�ޭ�����I��s��U�o�F����x&��]w��3�=*�b7QEp(#Ud^-��EP�SC���錊�/Tr���ѐ�F��o��8D��S���2�іq�!�z�C��sfM�G�y��do�a�����!}�,�K�O�����ޘ&��[��uMe�]��������'�����q5,�*��U�'N��{$D2(��eϋ*k�}dG�j�g����sƲ��G�
S85������.W-a	�_�fc�ˏx������R�&75G]�>&�\�~�(���/m�>��4ɻ�3I0��H(��ٹ��®�L8�]_.���]��o��_֪�u��zD��S5Z$�Fb�8e�s���A�$D��hs+V����ɤ��I���1��P�K�i,��x��w�Ys)z���֦���c���D@�QLZ2����*�3�,&�[�\R�I��y�Ng��%����Ǡ䪓Z�,hF�-��g�A�k�>���GzQ1���`�(�v��n���ۄ{u�(�a����X�j��3vGN)j����Nn��K�^�I���	c�:����ԁ��qQj&�^Tm���SR�8@���!�\l���z$st=C8�W�j�����f�T��Sr��&X�_��)���5�O�ۏ��,��4顑+ G~��Ta�3�b-������Oo�@�K�qqY���D0GHR��+}Jt�lzi_�L5�)Ģ�x5�Muf���@}���R%�.�9�si��ܰ�2���yq�V~�RP�y��C'�z�������
l^�r1���-��:�)�1f�Z�gWe)��%9�����X��Yo���YX��`?��Q����m���!Vɞ����ʯ✽#ݞu��0ܩ�������U�P"��Y�@:趸&+�y#��w�?�nŠ��{t���S7i˟;�3��m�C��]S��@b�����tI�f���6w��1��1A�3�5�p���9^���[����vl���{�PgO�<h741{�*mSo+�f��v�	ѹD�oj�<g⚑˦^z6.oh3��$X/��8m �ЙO�ԋ�_��sh� �/"�+GsS
 �����.��СfT�����*�]F�� d'(������K���uU*:u���PK^"w�KA���`��+m��ɁZP��ufl{��F����P�@�mi�S�H�IW�y|�O�eW�vc�W�������J(РS�h�5����n�B���>b'V��a垴4UP&���ak!�FM���9�����[���0�b1�tٯ*�C�yk<��o'�;~%ˤ�œ�Lw@�v�0�������bgo���$���~�y��X�
����#�Ҧq7L�wF
�3����������� �k3�]��������;G��!~ϡ���3��J��&���-��L�cIH��bN��u�q��%�hbS�6�{��]�-4�r���D��� �s����./���̀Km<mo ��Z �g�N��pU�T���J4��m����L�+�;��^zǐn����,q(�gv�5"l/�Sm�?/ �A
y�%3�oVA:/ā��G	/�F$�BWЕ��G�_y����� 9�S�e�g��9L��"a��9��(SIZ����[4��W�����C���0K? �m�a�`�1̀$d(��]���ҕ�ʢ�&C#��]���A�0�eg�c�]-���E���.C9i�-��|��͢��%5�M��ڟ�O�̱4hc`�Hj�&	��&ys-�N6I���̲:��Hm7�5�^�bW���m:�RC�f�ٗ�WSx,U�[}�q	 ��!SJ�4��c�|>Ė(�(�����t��_5�=�U�n�����'�M@�V���u��](,��l杻w�ܾ�fEGh��ȱ��}�C0��"�7�LG�
v�MA�J[�y�n ��@�c�U����^Z�	�y�d�Fec���8��qQ�"S��e�*���\����iX���9�M�Q����t��Io�"|�FbgzY	�w�--.�pzD�Y�s*AW>�X�Ou�Z�+�/�������4��6��U�aL�mB����>𢡄4�̲".����.��M	��-�/����l��?{}��E�ZtmE�4�j5X�oB��CrֺM`9��	���b`6)T !.*�bo�� =�M�v2f��v^��~��o�g?��:��O��g�a�K˸����@5���� ����Ȣ�������l��B�`�0<'����V���B5�h�T�b�v�:`�m�}�����/o=A7b�T�ǫ�<\d6� D%h��6�Qr��GUm<n��Ϙ�A�����O�����B�َ�8����x���VEv�ɀMx���ޅ�E����#:sR���i{gIkH������<$�REj�͆�� )RaMgT�a�'40P'���X��UL��Y�&��-G7-ypx3K��|~�UN��ˉC�=�/0!Tt�s���Wb�̉�Ʒ,����$��X*0;�32�R�(I�;Z�'/��iU�jaT�^N���2�H���tئlͅ�/~�����([��tyIݏ���˕�N��t��Kp8� 7izπ)�  ?n5x#�e%DY�@3p) WHhNNt�"\KS��~Z=ӉY���_�|?� �wyǀ[�_)͚�����P�6�Z�^z\M?i���>'��L1��'��i�濆6�w�Hǩb�@��?�~�Z�O�|z���Zr�fƕWN�� �2z
���c*�5@���̅U�V)�ۿ������e�/�⨀�\���InӞi�%Hb(�=�</%�2@������`�P\A�-A�&�A�ꏥq�
�%��f#|�_�ؘ(a��.&�;;>P���	7�78�g	���`��U����s�P�nv�67X�]F�������9�L;^=�2��b�:���?X�7���<�)��Ĝ�6�j��x4_���.���*1n�7�����v�`Cl�����w���B�D��E��غE��mG��Z7���󂐪`�++}�2Ze;��mO�w~���?�mm|��\�G6i���^���ū����)@F477�(��zB]�!Ô��6AlP	�(H9y�<�s�(kl9i��^�# �� ��I􋺛%��1Tlf�9��y�n��P+�/�:��F����¿t��Oʛ�]������y�$���Lx�'bTI���l

��\�R&h��݃�i0A��
;\)P��)L�Dʊ[�o"5hɇ�l�ݵ�����AS���\�$qA]K̍�.]������wy�Q�z@����&6�����H]?n���RwDRkl�2����jhMꛨ`��X�����0�~Y���k��,��ش0HP0`>�96lpU�a�t��jI ���H�r��h�3͞O�7xO�<ͱ�i"Mn�+k�_B�1��*�E�Q��s�=b�<�^���?�FrD�Ldd�&~G�����עj��F�	�i2<�(?�wɐ�һ��oզ���\��퀲aeRT�6m����_ܨ�!��m�J��Ą�^��-��C��^����Ywqi9P�RX���76ٶ�7�Q�*wN���pr*����'A�e��(�V,�Mv�uҍ�C��[�e�*���]s�5��<�ܟ&��ό�'���_ɲ��cg��v������u�����f�$+I���8�f]����?��E��h�ڋ����c����e�"���<[zɑ�,ʓ�	Е�����9��Yy�U0�*pk%�!�,�KsI�b)]�,~�?��:��떟ڔh�<�^�h�eQ{x�_�U�%�~�� �ä�y�S|}�ȱ�0D@
gɓ�l�C�C���I�Ф��W7S�3z�P���9�)+���%$����7��9�v�2�9���jg"�]$��es�`���gw����j"h'b]�K'���9��}!y�:	c�~�_��+P'��M=�C����������lJW�ue2N���1�0+�̌a�2�sɕN���2$��O^%x���z�R�-�u�Z�A�r��z�����6��Q�i�q�N\�A���jы���;��ۑz�W�P�5@Q�����7�H�9p\	٨Q� �/��{��� J���Fyj���;����=9Y�ǔ��Ȁ�xw j��L.x�]�����, ��(�%��x������Lf�c�A�lfjG^�=��k��Xt���k���.���Hi K����~#N��|ì���Y����6��Ԕ�;e]��*�FF�Lt(���V`K���=+�fⳭ�p���\�#7��3E�������][Tľ�2����i�A�!3�����R�r�1�C+��Bpcv�t��Y|3�$��P9�xg�Oﻑ���Ǖ�)�i�ݳ�͓�w��k[ثae!,=�7妟�������O{	�q}����ˇ]�
ah�����:�Y\��M<(��ks<!�$����W�P ���*1|dp|��7.ʖ*�)���ڭ-��S�x����E;�T%H�YӉ�(ҵ0.���J0��y$�a���[$18�%�d��ڭ��`O]4����,�<X��+���0�0�ID�[��om%�G�g�MíL��?o7u��
�|�w��_�fiUB���c���6���7�:�Wq^'��d�e#��0v���X������O���M��5���q,�k.;B~�_�'��(w���Q���N/�N��u�9l�\�/��ވ�>���K��u�ѸA���e���Ͽ3%Au�â����F�.'-6	\Ҹ���~;[֝*�M��S�,U�v��'n�� U���0��Q�@�_2�1K�A
��Ǚ}3��EH>��c��-Cm}g�j��*�-��'nQ��`ܙ��4� �b�� P�%J�@%$�j�R���wj�l���=K����.=ۧ3!L'�1�!�5�'�����M��� �8=�CT�2��u��� ��/\ƺ!A��o>�h�&_u��[s�b;Y�!�`�cğ2��dF���T����]���<�=A��?�йЁ�Mpũ���u�����	P��D+Ђ�7�	sX��N�����/k�|Ñ�V���x�j�`������I�)��×M_z�]�$atX{߂m��Һښ�Gc���䷫`��ׁ�y�y"�K�G����
�����]�./��jp���=;,���'"���P�3�3�1	� ��"f5�i�	���s�s�!#��L�Vs��f\u��c�/+���Ċ�P��j��=zI�Q�⑻ �?����7+;�E�wDC��"2x,辜!���lY��|r�i�f��(��QMتba�[UZ.fm��X�pD.;w��-i�hn�E��7A'����Z����l����:\�m�[�����=���L��60$�R
W��\���o��FC�P�O���Gs�Py.��ܓ��n�]u��u'����Mx�Ĺ�Lh �W�1߭��-�e�o��;���j��:0�
�H��H��ƺ�
 �</.5�V5���;�f_r�g�U���ܙ�	k|x�j��}-#w��\VqlIĺI�����c�z�y�����?7�<ܜb� �,��.m0�4��r�ߊ� �ܴ�5 ��<Xm��N�%�rZ�8�l�1��[ې4�k���{Gç�R���.���O~Bu�SM�b�lT��FIa��d?t�&��h: ok�J����!�4�Ϲ����k��\N-ݾ|��!D���K[��	LPkxJ��f�}�� 6�:� �Aϻ�֞lL��� �S�$	]���<ZNV����y��^3x� ��}�Q�Ճ����]��H�v�T���*�ߟ��(�&v������h~{;�;�����>P���+#o��[��L�`��)[����z秈Xl�}�t����=�-�Q���V�n���R6;aFx�