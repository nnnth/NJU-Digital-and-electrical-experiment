��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t�3����+S�-k�Y�C&���t���$Cy�u�4�>w����7&⇀I���$B����;p�ꗕw��h������2f�lw�ex��զg���}�	q��3�u}(�C�j?^���=� s�r/^B�[�Ĥ� w?� �����['}T�X�~l�{��A�����sb�,����F��g�F�����qZ���,ag�XFHˊM������(@�9�O�
�� ��BE����1v1�obS����&c��$w-��撴D:R�Hۡ�Ǜ��(�BxL�r�Nb%�f�ۯߟ�_�i�=l��pCSub���u��d���x`����Wɋ�Y�gX`��|c�é��Tl\�y�ÇX����`�'�7�Rw�He��p@���m�0�7!�! u�{#���zco�tƋ	ZG��s����#\3�>^�XԐs��c߭t�5w�^���	��ڪ���i�S@*�0�ޓ����'+�*�r{6�<m��-����?V=�S)R�޸��T�����\Z{	�,�t�-�M���(�|�"�0�O���'�����WcBfM�,z�Iء��:\���;�k�«tN�n�?��������^�V������n��E<�,�c�krE{�'��Q�e�2�	��(���mM����4FI�?A�{'�z5��7a�G\�V��fEkE���|�t<��P���E�ãv��&�Q�r��{��v�A"~|�X�����}�ډ{Je��� ���e=�V;�u����5j*K�" �Wd>�_ͬ�/��+���B���7.��v~k�_Vd���n��'��Z�򋢟K�*e�(�rX��o������B�d�]I����D����*oI�{_#�J� �������.'v��щ�uܥ:����&����8(%e6���N���M��<L%@�^�Ʃ��N�`�d�7�96u�q��l��+����oC˻#���[-��ȱ�rJu���a�����6�0L�k�
�(?���0�2��\dύa��L8���y^n���F�&�gw���G�YgQ2.�J	��֏�@GE5��N#O�]2$���+Z�z�l����"�<����M��<=�)��<[�⼭!FTE�:��V�̢�"�aMt���Y�R秓U!��rD�+n~3bǷ}�vn��l�Ɨ`�@s0��s�]��_�:�p�r՟�OS
�D�
J�S[��v�N@<)�6YDW*+9)B�>iHl�PyhG]^�d���=&x\�/���sw�^��P�r��ZB�� C��C[�������eF��iP�Y�,��/3�o�
>hg�e�lg��0�#m��Z�W ��ת�B��(�9D嵃���m�-�2M��Z���#8}=,�dx˜xa<��)َ^��KM8�9;�E$�EM�I��BhD�6|}�i�I�pI׹zw{�� '��<f�}�����o��뼔��}ZV�h�8T̫���+nmɷR�T�y���y�u��f#�l�O�j=�J���	< b�±K�}�z�k4��.&��P�����)?��ֶBS>�Y~O��j+���ջ�c`0H,���!vS2���� ˢ�p�]Nv���Y�����m�����/o�aU�E��c(�b�(��h�3F���0���y�u1��}W{�,j�JMb��d��b�7�L�������lM�$ ���ɵ�!�
x�� h��M=k�"��E�A��#�� @�EOE Q
�b��v%b5�unH�h/zm�훭.������H�M�vd�%�h&J肧p�������ۨBX{p^s� sc��E�p;�&���ͦ&�W�9����4�5��X�MC�VZ@�Mϳ)����w����=Z�}��)8㮋\�imK��G����ց�<#�ZQܥF-�����o�@'���}ψIMֽ��O�!)N1��d���v�1b�$����e�ܶ=�ٗ��=Zc��R��?�U{6�J���&����NM"5!f��W|wq�@H��t}��`?�a�8�	��ɰ\b�ծ�І~��ڟ���v��t`�u����qݓ@�ưuy{��[��
�hg�Y�*_�gT��������D�Y`�0v�΅K_��2��B��C�gV��}Ng����J�;�/X�WL3��յJc0�"}3y��"f�F%(�-����K�'�L����b)�E4q�,��5��2E�5{+��h/M���Q���F�����tTp�o�h�;A�\������4�K.��hG�l>Z��]�9z�╁̂2��2�;t,y����9<�q��a�	�'��H�*�G6��B�+��n&�|V���k���+���9²l��/�M���;���#�U���u�eq ��W�8�5t�'��v��R�}"��#����0f[Z�y0�e�h�-7O:��.��͒�z�}{�i��������g\�"�䄣Lɟn��x%b[ V�p�(���{A'=�?�Eb��dk�f��s}؜E���R�<���q��U�t����2Z�Ae��ޟ�6��]@~���o��t*��BQ>�i�<&$�d]ݣ�p�2z��w�>��H.o�.�/1��p>�(�ICra�~&��G�Q���.�o�>0�.~�m���������ģ��nn�y����G�_4�_"1X��Ԟ)H��oT��V�8T�{��9��ՂgJ�F���Ӛ�����]�7G^q����S�0%;I��AB��g�a5J� �J�E�\��w�C	m��{�H��$��d�!a�R���?�xy'}�8���`FiG��ҕ�ɴ㿫�g��w*ǯx�y .@{�Gi������P���1ߑm����=��vו@��&?�9�v��\B?^�D�SYY�$GE�h�0R�`C�����o��헟6��l�'��s�y?�0'��Ch�}y -�}5*;:�΍��2­���� ��>��}�%p��F�Ñ���0��@��I�ILq��l������$�1s�ZHR��}k��xcl����AKI�-��QI�o�թ�7�Esќ��ΘW/��:E�N�^Zk�`f�����M
�~p=��j^�c�dwҿ˷op-�fx�ۤ+�☑l}+X�F�;l����:���Mr���m_��9~��~�����K�P�*ؒk��IY� ��Z�'EDhV.�&��0=�_E�{$l0�*����L�#1��꺺@�5ڼ���,�6���`���(�:_�F�Ѡ�D\��_��l������̔&mϸ�L��ɴb��I��@�t��ӅK.L��V��ю�b����!~�)�I��:9Lx傐�NKB��M��?������\PyW) �ĥ��8�Rc�8����x-R?��5�?NiV7�Y�rů�LUs��ν��`��(����ۚh۝b�?�����^`L��x��n�	w�L�A�� �L�v��KvG�vxl����gNDܾ�`��=<�o���u��>�Z&�'��@�m�:.AIF 0�Fq?��r�8���Ϧ;%<]�޳5)u�(W�a�-�$�@wĦ/R�%�2��VB�?#��dƁ��,M'\;�5�FFF��` ʄ���1�>�!���q/��_�P<�v���:4Vc�0�0Eh��l�>?1�7�N���"j�}5Yt�G�*���O�B��C�/}N�A,���`A�1�6���/ϙC��q��
�
8<y���T�и��l\Ub������[;���I�nؙ6�!�ek A��&J��/xq�1�E6HV��B��B��a���ø.�i2F)b^��,��Q^!HJP�B�Z�ܼ\�N��e�4�qiط�va^y�?-�|��m��RF)����Ӱ&�y�@���	CJxu�H�����Q ���;�@2�_b}�g2�͡
�����+�`HW,4� ��a.nkb�@�ۍ�;	f���թʞnĝ`�u/�*��U:.n���N�����?z e�xc�(�����$�hM^�7Y !�5&���'��R�z95�%qB���lJ�A�Ze�Y�7�p���f1��<C��AZU
͞��'�Og�*�]�����Q+�*<��G}0�ݘ^���N#ȼ�!*�^c���`B�#>�˛
�vL�^^�su�K�fR�v��K���V�,-�����H�єd:�8Z��-"�/�S�D��|+����{�����e�#��\�*玊�8��#�}�b=���y]"w,ڟ�B�wp��w2���*ؤ�PEr�ZK�	7����O�|t�	�G�f:G���6w�{����P|��⾝g��+. �`�(�ЄWAáɚ����@4���4�C����4�+L/0`��=Չ͂;'�.���L��]�L����p�dݙ.�&�,l,�GJߝ�B?K�΄9/s�����Yr��ȅ ��:���x(q?����f~�j|Lм���A��K�Ƌe%m�9�R���q��sj�w��ܒʥe�o�����Hp��w}>^O�?��mH=�Ԃ�{����6׶��*��G�
�j���z�G��,$��4��{����0Tff+
j�Ctմt���ߩ��]G��o"~����k ����
*9�1�~��"aG���_�-�;��t+��M�s��uU\��=�VȤ��d�^��¬�b �+	hƂ���QqUQ�	�c	�@x	�Y��4�4
G������V%�� Y��k���F�=J6�͗z���N
�2	�&�KV+��D����願0uv�>7a�p�$��	�:Yt� �k� �&?���Μ��ph���@�VC_�z�R��☄B�hA.=�DT-ﻠ����y����,�bh��m�`�ዘ%#=ڍ��׸�^^�|��I�u�����z>��/85�7�?���S���2�"p��P�m�2b�_aQ�����t��_̌p�2%"FX�4I�<����5�W���-�?�:�Ҿ/J�vG��<��O����Ӑ�z������$.aqnV��u��OVz����ʣY �o�cl}!2d9���{�x��@���3Z�Z��
�<\8�L�U��Eҡ���[-3�=a�y�1��h���V:hO��g $��;�o׿�P��m��/D�wj2�9����Rק\�&���d�ن����H�^�?�>�ǚ:k�nF�[��q~Q�w�(��L&J5C_�cY�j�Ft�G�N�	��9K��v��������Z�����4/խ�Zf�����E&�z�j0����m'5�򸓦�I.���t�S\��,�j[W4
i��G.�x��>���u1L)3d_�M���w%��ZU�[���Y%M��jХ����:5y�{AT����~:O���2 �\\�:��O�p���<h{�v'	���SfK$�?7��x�KOK`?1\����Gq���W�=���iv2fꄚG#��R:cKc��J��eu�*Z���6��@���4>j�����+�G�b�9lYül�ES�"�q�B3�Bre�8�fa�%:U�u����On]|�W�
%�����I=�L�D/�rS[��#X����hAJ}5tS[��ޮ6�{�Rr����6CC�v����U��5dJ�u��k�Ʒ#�`���`+֑���Yc$m�_��^�?�.�����din��QS�Tq��4b{_U�����m�h�P�L>z[ݧ�\����cŁ��S2%1�aGX��
c&y4�0y�٦(;�;ȥ�F*�E��:�h��7i٫N^��TpNVcXW�j��K' ^����Ż��ϖ�{56r�IƤ�t>]a�j��g�C���Je��l��Y��Mx/����V���Ѭ�׬ow�0��<�4+�S�͙e���;_�_.��$|�2�#��D&M�3�պ�8����H����p�:�֐�V�P�l����G���(����+����oDC�~Y���ߺi��?l���dy,۟���C
��t*Ŵ� ��k���(<�Z�ѵ�_�x�yg���$o�s���|w-?co���Y�:�3V�`@�����oo�bV�Z�m@��RYC)��|�I��פ�U���@l2��| �C�l5R��P�1,��M�n�'�V���9���f�15ˏ�xT��^�l[��l�`܉��Mz�/��Q���98cS#1��Ec;?ҝ5����_�I�y��@Ld�$�0��h8���� &~Q��ԳB��	�ǌ'G�j�,����Zo���J����?�]�@�Zˉ7$�^"�͒��%�:�`Gt�9�5p0����]�6�/�@Q�E�O��m�\//�Nx���3(�E���Sź%����@��I�St�����b���0��)�/�[�]!�Yv�P�$��ʏ{P��ۯ)�_X9��A�+$����_H�1����A\q����j�Nm��1����?WIwG��Dg=���%G����-�,���Փ����ت �`��؁9�yFÀ&��� D�GV�oޘʳ����Ov��%�G�ϫ�.缝}�tUR�c&���(I]�!�lr*� ��AH%��߇�%�����*���k�ϖ�Z����^^Ѥ���n���5�����yB�%�u����<$N���ˎ��/*�fl �-&[���s�_�㶽k���$ҳ�%�@�M�m�ō��v�VBlj]4U%�nms}_ȠM
^e��M!{�J!!6h�i��9���{N������rމ��,� ����A��J���H�h�W����f润��(��{��7�8?r=w� 0��gG��v�D��Q5,���S	�թh�i�d�];�&�8��UKn܍+��4�O1ZţE���a�	�=X��:�x�
��Ѧ����k��_9��לʧ%;�3��ɞ�J���E�4d�+��XЏfd���'Ê6����uh	}��Y\�U����b�0�A��\�e����rh�y��)��iq����O�ȡ��5�Ff����C�5��K(�Ď�^���JǄ?g�B���6�o�x{�L�ʳ�~Ƌ�<�E܍#��(p�F@�������')�$�������eW��}L�A\�8�H���z�o�w��?�:s��Q����F�^+[!=!�6��)f�P(A�&��t'�D���ـ�z��`.	�`3�r�4����=�fU�'/}챤��0\194�ٰ����+k�6�oKҲbL��������d���8�*U�"��6�OD��I��7�e�\��n���^k�{���$���l?�����s[� -闖�evw�P+��N��2b["p!��$��y��?y�6o��+�R{y��a�Ё�`���\_WxK����c���=�ݞv� �]��f�ʛu�7������PqI�9m�Rv�z�잡n������0�8`a���kF�R�;�j��h�3 �~���A��sّ9^M�9�Y��yn�V�3�hi���+�©�Ȍ`pI:4�M�T�������p�!ȋhw�=%)_h!����pL����{8�Y	A�H���2,~��h����$
�&v!�E�%о���l��F�"��[�Wp1����W��d��\�.��ki�Vp�1�S~��9��fQ��f�g�.7�bH�pQ�&h�J���"bj�&�E���U�wWVV��$�����/�&n����DY�d���T�ڗ���������A��\�b�@qحF\�,f1;�Kz�g�l$�-0nt����'�(���������"�Qᮠ�7������+�-KnBtөP���p�7+;���O�$m�袚�X/���U��k n��$��ϓ�VY����6e#�B���c�r;���r��}N�<.R�����s�
��|q�"͡�=|_�تK���I�����~�tK�+xԨ��c�p�Q�������V]����q��"�wjf�Tj�� �c�zΣ}N�0%.��f�z��͇���f�������1&��9�(�0����2T�p�s����/Q��Cl�HG����4U��-�ɱ$�W��1�e]���~���O��-rQ����fwkǸ�@]<�p�!Ǎ�P{9u0��iGG�.����`�t[Rq��."�H�@�8����`����ʉ����6�P�rV��Hh���C#R:HyT1l��k��x6ўNX�����^u��,jy��N?t��/�-A)�XI�̘��]�洃��-Q�Mi�����J�7�
Q'��s��f�����2����eu�n��K����YI��c�[���5��աC�v�kO2=<�ߴ'���|�]
6�t+��������	���j���3�v>��WE�-ֹ���n�eK��o�p��Tx����dꆸoL�M���^$��I(�����㇃].�^	�K���Y�}�s3��
K��@뉳c� ��,��ez�i+zt���^��0N�#$ra #ꆭn���~��:�p�(�_��!��=����	��F<
O�����ߓ�����1�}�
�L����b��$��a�Y��7�YSS�8��k�Q����(�GHF��J�ZC�rN���#�vm�.P3�������8�C^Xxn�� ���Ų���e��@�~B@��!�n؄˪K�W�����.����c�a	B�P��[����*�{�����ad��yԚF��|4ߊ��} �qJ�2dҾ���{9���pK�H|ش�hm4I��a�A��r3�
^�4>w�z8M��=X\��S+��"�!phg`�Ǡ�߉���J�,�1Mq��4���\@�I����i,�S�EE>=�`��N��_#�v�p<<�pQP�$���sf��o���52t^8�?�s��Aʭ���3�0�.H[֐��X���})��D,�3f��mr��7�w�&$�5a��>�0nL�]�~��M�%�T�.��pس=����2߬��l.��>��h[D	��{kJ5��R,�f2C�a�U��ftƦ�H��7�]ސ�8o�"�������!4V���f�T��e�)�]7މk9d�:&��[ۋK?��E�~�����6�X���*#iL�jC���qL��M��RJޣHvl�W��I�̣�id����لG�j����]��fF�8<R�	�9��� q&:��M<�6�nC���\śSw��������(�8���!��I<��^��S~
��@�sF?n����k�u�`&\~]ǜf�����������Z��/���ڌ)�Ȯ��b0�_��P���}��i���~>�{vam�X#�5�S>!�[+d~K�R�P8
����u��KC"�CD*�o��h>��Gu���N]
gh|�k=� � ���:^ǿ��V���]�����M�̿��º�>o��a?h�K@H��啃ZIw@Y�x�����$o�����!&N�3���Zf��,?�����}���р���/:�w-vX6���W?9�DO�!��U�K���)���_�ˁ�RT�����3ϑh��/����������!	�UIL���q�2KpI1�1�d�t�!�y���s��`�߭���'@��UA��2�B�CvD�E���[�6o?�rF#��I�Yr��C��*b�AtH�4#�����|���&B���'Z�V�L'���<�~H\��Z��3���E3K�s)̃'L���#���g����X5��N�+:`��Wu��v������%�Z^n��"�?ླྀ�n8��s��9��n'"��l1��`����϶�v9"��m.�^�-%>uC����P�7����-��@�'�9�kr0����HF��Dl���$���\�F��<{���v@��/���z�)��@ݹ�E	�F�Kf�=����w��LoG��̺��'�n-J���(���tU���ؔ�d�I�~�X���Dj*����!�<+e���I���q�k0��ʗ�F>����7� �]$����j��C���E�F�z�4���kI�g��咛[הh�m�����	mx���0���귻��޻C��2c��Pd�d���\�G��G�P���0f���hyE�6�l[��T)�;IpH�^���Ϗ�.9(Q0�x�~v�<f�?���_���Osk��f�AL�(�@�7V����S��?���-���*nA��9�����'�����}��;[��4�A�os��fι yYR_������`��A+�<�
��p�*�@����^�+zg�R��hs̗^���:8^�f9zB1�ƨ�/P���%.w���.��ι~��3��"��W�������\E��MK����Q8�w�1�p|�[�WS�,M�#��#'��q�mR�t�?�ᮟ.0l�͒����!i���Gg��Ǉ��t;L`��dVF�.9k`�\�K�8�ҫ�WȊOhծ���'=��TD�QE5l