��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t>g;G���m��7����z��z�[0�� �Z��PͰ�Z[GaO�p�SD�����s�|�,?�|YrW��϶�h$0�&��r!��Eٜ�勶XT�����'eJc�������;���Pu13�O�GRy�$��vH� �Fv�A�ң���]ϛ�*R7���nF8F?�7��+�Z�̜/�;���,�<H�|!���>ѹc����Y��p��y���u�'��4Y���>�l(��OO�!.�!��1�S
�N;D#�ɱ�H��D�h�7@�2�a�sm�9|�F���
����� \��?�
jЍ���a��\��n�*��VON}Qi��[
W�O�Ӧj�Y�~�1��ׄ����)rx;����T鹽1�%58��0�����v�D~��v�@-���H�vv�H�3xWa�Y�*8h�| ^l��;�GႯ��*�,'��1��d	k&Y7�Ƃ@] IN�V[� [�d�瀣7p52/�ra+p@�ݹ:	���3�(Qًzɪ����E���	�v�b�v�������g�~�	׵k8�e��Ȓ����K�u�������Q��K�����D���~��(7T�?�2�&'
���t@�)<G\J}������橜����l�A���}'�I>���&Z���zJ������K��l?�T��so�XȇH�aT���jݗ&_=`�୸��׳���j�Y�C��-�h߀�e�q�D8Y"t����U��u�զ��G�U'gA�a�]���,d�lm���i����NA�Vt��8�����W���!�g��|2d�{�w �3e���t��2�#N�*��,����"�˸h���� W� �*��Ši���&�;�`��y��D�l-�iňp,�0����ǽwڸ���'x¬��.�����Ɋ/����=s����c�/Վ?p�hl�)Q�����k`��AQp�QOd�'����0��@���;���Wttj�>�Yn�d0_�j��ƀfYݩ�p����s�	Yv�k��������%���K �������&��i�a��,x~jl>u����>���^���nB2 ZN�<��O�kԬ��𙫡"��Y$��y�*��8�'���j���	����GW6���J��rב�q$��$� v��7O����yk�#s$�F���P��. F|6��Y^�5�*u{�Fy����؞w������Kj#�H[
�q��H�� �8N��3�a��ު��bY\$���at�TוRnlR��]��Jp=q���dP���n��g�z�8��9��4(�bu��aE�S N�`��y�&��C�2WTԌ>(���/�6u;aK=��?v���y�95%ly��c�7����Ce����$E�y���V9=�!IFq�vӵ�?�y}'Y�@�Y����K�'��C�O: ���g�LtK<�L󪜮�o�{$;��ww��J9u��@��hYB�7�)9����!��4���*�uj�b`�-q8�M9�Q���3���VBAfR���k�5�6z��1[�|\_���s-w�2�+2I$�J�z�ɺJ��8���T�r�w�����F�!��g�M[���|� �e�4D��K��c����x�!�yT���'Z4������L:�Ww]'l�y�A6�4~�.�-iH#��fv��&.J3Ԭ���*#�C�H�P?�O��j���]�*���㍼��&[b_�S�L��N��]FnE����5_X���Bl7K�.ځ91�Q�ӥ�4�U	�Qs��n�����0t?�,Njn�n��+.����*�yP^#QWV�J���9U�!k�/Q�R��ΐ���t�nX���ؙR�>���}��]�7O���A�aL��/��mr���*��$��2脝��^����&c��7/�h%��(��'�����QD����&��HW�-���~���n�4�4vwq��C� "	-�<���SEHƥ�+�I���9B,��_��z(��������w��HƳ�����K~s���N�^	��$}��9r�z����\*�4���]u_+���n�V�Z��Av��z�	ߊXM�9�m��#��t�ϳ�M�A�2� PPڋ'a��y~�PнVW'����P|��Ao'��Zg�7mmĢM��W���z��;k�/Hw_L����^�.=a���
���نt���'1)��0"��q3��W�I������=���n�q#��G��G`��D��+ؖ�?��9uُ����1>V�um�������ؒH����Xho3�^�����u��łr�g�{c�%٪�z����\�@#4���>��z��y_���T�~?���rC��� ��S�?��ë�s#�� &����9��b>�m�=\����	@%�ι�����ؠ+@��ؒ ��nZmI�AŴs��A�ܭCa�x搿�}qH�׃邻?S΋`SP���~l����NKF@-�4�'!L��9�D�Wt�5C�/��Ǿ�=��ҋR�9t�:�P��o�CZ����8����fk��M�EM��l(�7�L:���Q$(�k����MG��j=���f 1p��6���6�E��*31��)��G�k���Ń� _�q�N�k�s
��ԡU�8�vi󮇈%�W4��c�+�"�6t�|@7�CHy���1�P*ó׋C֘^����t�AX�,G���q�����_�~�j6є�l��L)Ti��v_�t�������)�크�&��o@�ӱ���f�������u��H�K]����ԥp+�e`����)3���FƬ=�g���f���/��ŎvI��֛�LO���Nt&L�8Uny�f�N���
�[�����"s�v�"%$�)g�uS��әC����:_7�,;�~���G�ОѢ
NL�J�E�v7��w8u5�k�)��L��a���܀�n�0�8~R0�bvzCTё�N�C�gߘ8�I���U����^54��w�/Z�=��g�y�/�O[���l��٧��K����y9�N�߃�`�L�D��o<��S�_$/�%�&K9������i�wvD�0]�ռ��������˝=�Y��6��b ��w#�O���0�}4A�Uʟ������[���	�D$vP^���nR�2v [��bc�R����'u�h~Roh�ʤ���#XpqH�Q�1��δxH�z'P�S� ��ȱ�n�Y�;�+��	�\V�����c�(�� WK2b��.95־̓��۬��/�&��s��C���A��s�"�2k��1b�^�T�p�z��ٴ}�|sy4fU���sv�RY���Ug`؆W1*�L?O��c��
'3w�ZO�d��0��q�����#f�q����n�T:���[d�]��5)%�?��.���!ͧ����!'/p������� V�{�d�f��a���|?����b�'
�t��86��'�So/*�����C��X���x��ZI�~������ _��w�BH�D����p)11��&`��X��d:�!�-��z��ܫ�Xcp��$o�6Eℑ(�~�����.wpx�H�s���c����VE�ڥ��t���_�dI�����P��[��RW0~�fo�{���l�ϱ��k1�=s�D�)��璣B��7��mq�X`��h�2`C�sq�� �*��qP~�ܺ=�`.YR+�`]u���U��+� 2*�z(�w�l-�4�0��;_����f�3`�W�vOVzBܱW�⻘�������H9����{�����t���SֳH�5J����!%U	�iEV�K�yaM�/_��5�����x ��ŘbO 5�	�.���9�B���j&lZ�Х�|�t�bdҹ/^p8�[7D���i:�l&�QD�`�.�C�$�JG#X��+V��RV��a�{Z��+?߯h���uύ4*?ه��顡�
ʊ�ש�M�i�����c�u�H���k-֩��n�3��\�밠ũ�:g'R�vj5�7x�̐����G!-���t�%�1�Vɻ(O�cM0cI+Y����߃ӄ�\B���K�)�d���y�S�P�ǵ��Kh�������3d,FtX,���hH.χ���$t^�U���O�V�db���Mj��L� �'G6[�K�*^���ܹ��x.S�,'\{N��ҹO�bM�:
�!1$o,�h�q��U\����S�|LeNV��{BAh��G���;���-s�촣o����+Xf�C����QR���>a�iD#B��A�ȊT��T��i'gN7�G@?jS��g���uK���Im�nϖw�.cL�Lܜ����|�*o!�]!�	�a.�svz��$8��ǳʕW��/�e*�|�����:<T��vF<�.9c��.]p�=��o�k@�j�91��,Nh�ǽ�/x��k̵�LI�����I�}�-�+׳�Q�-�F�?���0.X�G&�5�J宏5�bSicT�j�/"7@3�`X��B4�����9<�k�^"=����ߒ6�y�=eR^�������a�p6�h>H��v<��[���m�����-�/J�>�����=�������MՓ��>��姣w8��y&\�� ,W���hY/�C�1R����}�7֍�v���F���QBח�9K6�a��^ތ�@��Zl�m�*���WH"NEN�>D�L����y-��_�K��<ԖY�>��Q�9���q(�D��^	��δ�e�����*�U� v��3����%:GEz��k�Y[F���nR�v:��%J�n��g��"�Ik��"t/��1~�ۓ-��rʄ頻v��}F���n��{��Bmc�J�^HM��,���	����k����.y��@��nR�w�l�x�wڋSz���#�0�A�?���*	֭�*����T���ڄ5�v7۰3�SlP1U���}��p����U�)����G|X��g���r�8@L}��Q��> �3�a�TB_,�4t(������N��(�(�3�1��ʑ�\�0�A�y��VjcI(�� ��U��u`�������v��
:���� C��c�)�M��_��0uQ����lj่M
za�u_db�aA�M�2<���:=��6�*����t5����`���2�� ����?�1�"���<LP|܄��m�ٿg�M�D 6Q� #"ǵ� B��{��9���G�9�rn$���z���������Q0��f6�}�#띄U��+D�hI�.%��ɿ�%2�y-�;F�n�=���$�}d��v�,*���EG�8��.�RA�����*����A� �g�#��5X����q\N�P+�kI��Af<�k���Y���\:��K����-ܺ����t��X�(�I�%��i�ꋭ>g�3�6\9'�ʼN�ã;��!��K�'q*$�+=��4�FT�4�9�GL�>���k;�˲q��5P�	-sV���۸t/��ɸc�HS��D�� \ObN�k�,	nuQ���n`��#�F�w%�9!�tq6ߜ�E� �H˯���|����6���vb_��! ;������/-#$�Ywmݶ�#>��6Rc������SnɽG&�w��T~`i̠+��+�A;��s�"�p�{���|��0=Fb�U��S���av�Q������u#G�A�����c�ß������bY�w�;aS�u:݇�*� TJ#q�B��|x�l�F�$#|vI��;�J����G�l�N�`ϭ�r��n"	ز�r�ʲX��BW�J��&��<ŧ��f�t��/Py%�g(���K�η"��Lh�e!�3�f����HN~d�C.Z�g�΂�=0�4ԥ�8tk0�n�E���pc?-����1̍�D�X�=DÆ~��4�@�����'wR�{=�{��M�1��GW᲏ǔ��Sv�Ǚ�X'&D�j�\
o.��NH �Io;AG��J��P��g��VK#���]oB�����\m�pw �ȑ:�r��%9����XE�E� ���-�^���s' +��f�I U���$AV�|l=ɰ)�d�U�u^v��ۿ��h!�9v�:Bq0K��>u�ҎB����tf�1�b=�����~��-���"�[0@��/�V"��%B]�h��$�$�?���
���PPΒG�\�qn�KϠ!m������;���AB����N3=J��X��;i�2r]ѱ�c^�,m]��z�y�Y�F�,Cu�	7��(�R(���r�'Pbz��3>n�{ל���)�����ŝ��i>dPJ2e���
 }�p��_l�Ճ+[q��i�	1�)��S1{�'�YZ��I����2��B�<9���������T7�C�:��
�@՛s�-���?;{+n��D�g\�s�[4��^d����}����茷����Z����\HJ�w�� ��E�?`�]'"������ؑRo�>~�&?�[�fVy�_��(����D%�'
;m ����A%<����5���9���У�7�/~�@����{|7Y���������l�S����������a�t{�_��IB;�v������̸Xv`�l�o�{�`|��-QNO�,A\����Q��t��k���*��\��կ�-�#�2u鈋�56~��@�W�:Pc����w0a"�d�)O�$s:"4SUD K1Z��������P�w!���p��
/�պr��g���"�8a#�����4�JWt��k����6|���!4���,��(�ƨU�[||���qsM��&�,����~(��#�sɌ4�#<�*ޟ�ZgC(�{�2&�{�RO.�f�w�;�օ)�r�d��m�,��|V�y�2U� �(:�fXBwD�ߕ�=6g��kzw�Ҡ�P�3q?������-��8L)Y3˰Fa�����,N�څ��i��;�}5��wڛU�[f g��1�;���!��Jػ���7����0�������o�,�����;��D��f	p��r�5��`�D";�����vrC�jşg��,_��������g��T���zf"��H���+�m��
����W�ˢ�JŨ/\Ȩ�ڔ���_���������r�5���X�c�o���Zn���'����g`3�?K�ߖO�7UI,��0�MfY�OU����'%H㴺≔��p��΅��խ�p�ps�u��X���Qd�R
�H��2vѸrަ��K1N"�R�)�Šo�M�a�T�w��$y�@y����&~Zz�5�ӆ�g���3|�����r�	�`����y��>?�6�?����sRaC8#f�I�j�n��ͤ�jù��P'O�(W�2�Z�b�KO�SP۪m]��Y(�8��*IItXά�6W!��v�>�ㅭ�dXr̊02hUG��+���\ Ac�*fMA|�$���p(>Rf�A������Q���V���	�'�$�m�7�'e'����6�߅6�<`�/�Q����0���u�_�yb���G��я>�}�@:����s�q�XǷ'�e��隤��j�έ�ă��C����]�h������Z�Cȫ�4"�,� 	���
'������S���B�?�q����*�D�D�����Y�D�L�n:����������W�DPd��g!<6/ �8o��OJ�7s�0����1ǣ�$�J֚����$GKY$FM�v�0e"�&����K	uV�� �3�{��>c�dJ�����lɾ���r�+�lK�R^~��=`]'���Ht�tEb'M�'Q���3D�@�zm����@ܕ�#$%/�MS��D�[�ϢXP�2�tt�
�vp�B�׽T��&�/�7@!���'�JR ��	T���������/��֑��ɰpn\�����5�Q*Z�o1j��.<x0��I���G�	�W
3�E�}FF,L�����pVSdp��Nfs�a��Ug�V߾���o�^��b�2����ն�ڦ�x=�/ϵ �ϭж���b�����b4_
���]�1�j��1;/��3Z���%�`�K/$�I�Z'5��P�-��GxI�1]ᴧV�d��(s�����B����W��K�8~�T_�K4��u��4��P��É�>H���*0�
(*�K]ss�5�`Rk���i3�����	���{�CT��Fq�L(<!�ct�����@��H������|�S#����T���X������s	�G8��V/��-�D Kۭ}�}]M�����M��袼Q���H�%��G�w�f�X���BΥx�j�p��9!�~R�C�� @�gR&l/�I�G�B�]怍�0䦣��kn���ˬVL<���C�ԙ{FS��Qk��^����г������ygCCw|H!��h����)��!ģ�ѻ��ӆ��� ��)[@�D�K'��m���m�^�� ��:����z�&�`WXf�}J��M ���)͟�`�Mf`LL;���V�#�5ɂ~_�ۥ6e"�+bभ���Χ��3���[3Sd����)���2:�p�}�>H��V����:r0��w1���0J�w�x�����]8(����ޚ�J��u1�4��V�75��%�#�0Z��Ǒ^e���ԩEj<oc+�):L9
��_4�8"t�S�Q����9��dܤ��7�T}���ʍ�{�X��9ض����\�p��Ï�,���1�˼BG~��ZV��x��lI�3�֛�T-���Z��<��Sڦ'������R@�
���K�Ry,�]��x&��D�7ғ�Z'�G*�W�v���Qפ���j��T ��������V��;-�u�_p�\�����5ڴ��	���#bn��WB�6|S�v�ZrλP,���y�eȽ�|�ldI����{�00r*{��}������tN��lq�\������,Z8$�q{�����=7��9�=��2�pX�0]4e@���'Vd�F�G���:i��ds?*�9����@��#�z��� 	��K�Ev��Q3Q!��Z�*��1?���7��l�I�^��P�,T��5e��5��M�TpP���f�����0�P���.N��4�����a:��W>�o�UO]������ɾ�x�m�Эݣ ����ѣhP	a����r��H�z�(�Z��MCku�"%|?Aq$z���i�`��39ܼc)�-��W5�Ooa�o?/5�0X>��k��Z�Bzf!�G*����֍	���P �U+}t_R�s�n�QEd5���H,�X7q�ɶ���'�S�6��O��6�����-�ٸ/ߪk�~��fF'�d�U��B��8fMS#�: Y�������?���Q\�*_�<� y���(K��k%��|�4�3�EL��~�S�Q11���;��Al\�G���Qp�P�9�o���đ��� H;p���������ғP��5��p�}�D4�!��6��5�wh��{Bg���C�û>$�E��!M�"h���ҫv˕���bZ�/���X�70�� ����,$'C&�,���T���٤):K��^gGv�`lV2��/&+�a?����+���(=�����Hd��CqQ�
�KCp�5;�˭��.�!�oN�Y���3���\f�H4�V����c���s[SW) z�Ӧ=�����8�������Eݣ��H�2'܂��Ajг�BV^�Qx��6���=H�-2>���ұT�kN����E����<� �6��d�څ��4�������c�Tn�x(���}N�(��6��*�p�YFזAg�2�����22���Ec&�-wV�N�m�HQ�Qȹ8�ZP����>o8��艇���*�r�#aY�>DA�~�|Z6�f���0e�ټN��G��o���I�*����e�lz�$>�Rb�J86��1=���}I�zч�;1SOp�<�j'W�K�	��U7	�Q;a;�@�L���ԐƵ.�Fm����2Q��%�@d���}�1��&�jX�^Ұ�����í6���_h�����8�7E+����s��z�e)�8W@�]�����2�g�ؚQ/��^�{��E4H5`ؘ�t�w�o���+(@�z5����#H����{��I�Ao:2p��9g��.Ƌ]�Z�|�v�M+�	#��#�� ����e��܈�=&;�2�$
A ۼ���+"�EQ_iݺC!�a�R�0.�B�I�`I4�f��㇌� �I��J�j����.�]�.�g3��;��Ӆ�\Y���+��c��\fZ�;����L|Q	��y)(�� �"��5�Nbڴb�9��[c��_�}��r'�43]� ��9`�<��*�~?{�h�0$�=�]��Y�N�-b���A}t,Y{��R�P�������n�I��>���R�l57��C肉��-��K��4�T��SQ��t������q��P�b{:.*&P��k(���RHKˇ_��X%O�����H}�Tn �\7�y�(v
s�~�R��!npqh]]E��EV�Z����ⓒz��t�'����r-�$r��nA�C/) �����zV�;�X�׍�:���;K(�8���`�gT���>�UR����~�rNr;zԦqA}�FA3��ȔL3ky�+,��)Q�hX5!�rk�<�3��2��*w�(i�45���H�d���O*�^�s:v�`�n����Y� �J���G�!��cpB���
�{<މ�ޠpOgcd���mM�����,��h�����ݛ���!�|�w#�<β�hn=Q�dU��ګl�@�6��ѿ��	��S&q~~�Z���t/�B;�$��W��qjέ?qY�Zg�"ÿ����,��z�����`��Oj7^q2#�rߟH�.��Cm��m%��w3z�r:�AG��
?����	A��L��Їfb���|V���<��z����~���l�!��#]�)��=��l:�@۩�����O͂�y��>m��&���_e4鏡�i4յӔ�x*>z�[���YPmD�0�����PKC<vb[�+�9��ݳ�W�].6N;���-uK�Y�P����f��U�J���5&ߚ]`�1KA#?��^5w��.�/B,�ļߖ�s $d���Y��X�k"\V9����&EP`&���KZ�o�I��κ'��\�(*�2�nA������&s�R��5�ؖS 1����(l2{��FŃ�	R��]�.Hnq_������oŦ�I6�e���jk�ꮇ;K�&97([�ɱ�Ov7��RvV2�����;UKXgeiqO��taA%,�R%���H4���t���0w�h`�}�*5e�F��9Հ��)����a�S�g�.�t=\΁�:� ����n�PZy�XY�AH�tQX��!5=D��E�2�*���T8�Ȳ�*�ޥC�鮶����:���m���?��u�w4����Y����p9x�.�j4h(�x6v�=��_��z�O��-�
G#t�޼R��mA��j�[�"��hC����"6���AoN�g1^�W��N}c~lH���Y�����R��F{1S���2�b�s�6����t�s�yDl�IEd9Qst����ԥ�kt���zP������XT�[v7Ԗ�|#|�Z�EЋo�f���>�6���~sY�Y��2A��	��F�h6�I�K%`���j�vz��=. �V���=�Y���E��2/h�+��rMԄ?�d�k�=+��S,�'Q�R��,�h�_���5�:�s����/)�֞�޶���`é�С��4IN�ʨG �s=�%�P����&�{/���~�C��̉{�$e�0)���,ӯk�S���w��\��>;Ե?���l�����n|`P=&�|�o�7���i!���\=�剟���Tb]���ˑ<Bz�r�.���8�P1���%��j���\~V[95�c�AD��\w.�#hk��(�o�<*b����b���oI���GT5^ܖ�U�����	�H��ؖ�e�2�w֞��E�:�N֔�DTM���!ݸMH�ő���F(d;��5]?��m��8���Լ���5W��;����-Iʃ�~��f����E�Ց�m�dR���*�����H��`t<�����M���Nۢ�oþH�`ũ�"2�ˊ�ki�	x�H���D�B�|�`(t�
!6?�^���T���OѬ�#�BvG���
q7_��0|��lL��=
��7�*����sx1�GЇ�X����=��{����������@�-"�W���IP�� K�D�!G6�ߧ��:�G�V`����@_?���5�����S�]�X��X+���>6g�
�p�- R�o=yhX�Z�ju�U�CY\$ F�{%�.T.u>z����>cXWy���m��� -L8�O+?]���y�RR�%6��T=rTV|��8l��_�9;$����	MNg{	���4PÈ<eiی�ELD�4�����q"�����s��?\�dx�R5�[����o�5Y��������=**��{
��4���ƺN��R;�?�@������/܏�[Wڬ�-R���2�|�z��������!9�[��$��:���[��<	�o�r&���NS��F���Â}wB�����h��y������[jǟ����A�������W��'Z9�@~����m�VK/�����A���i�y�����>��H�v�V��jo/�J�"Q}�H��<�꓅+��'��(D��
A������Vˑ'<sb�4�B����P��}@&�3�6?�7�Z�7&øv���Ƕ�/��וxT���|������LE|G匰����~^{p���yI=&��8�dE;B=������P�뎼���n)�d���~D��J,����ְ�N��{��>�6�˰[cNd/��a�U���aa�5����a|�t��(W��0{=~SS�8��g�?�UփN��]v� �����B���G2;]�����.v@�0LEV:;x����f(��N|��s\�\�H��P\[3���m �pi��YkF����_�I�f7���|�i��)�?����-@-j��AvT/��Ҿ�0�
��%����H��m��*_#�n�*G�X$�m���	�*.^+-�vF0��M2 Jl��~*,�pfl��8d�i�5B�4x�ZA�D�?B��W*��N��4��<M�#�t]����e���U����3�y�ףM�4}4q�I p��Z��d��H��m�̾�i�nQ-D��Z<~�1Az��	ng�G�z�R>^5�q!��p#Z1��e*@��6+�k�@��=JL�[�������L#Q��AJ�P�F����&�AQl)�3�����'kg9�w�(�uI�U ���F�#b��C;�|����������H�� PP��y��ij��o���b��,�����+�2Y�0�7�����i�O݂���Qy�y��Mr�1Ю���$!dqp �_���F��L�x�������bā(�vE	 t�����\�ǅf�q�ó[����'G���%U�Y?�Xn�^�ds/�P�f`׹��`��S卝'���f��~�C=�i�UM=<��B�L?����� �J���t�F��ŕ�L�'��ں<Z������J7LNZue�$���  ��V�����w��HI��6@��~lY��"q}v��܊�~W��y�`���������~%���{�b��u�"L	Öp�@�!� uȁM7R<|�Q�Τ�M�1%"ה=��S�<B��e���Æ�����ϖ�O�>�]�m&s��dL誨�)7>�Y�~t�i(.,P*{J��!��,d����)��-.�*P�=�(D�M�kM�|���Ek��}�+���74�7�D9J�&�ٽ��D]��y �s{ΫՌ����H��ĄCj�R����?5݄׌*n�1m}[�6�)y>�����/�w�ja@6a
d!�a��t0:�"b���nk���Ed]���`"#����#�_�xʻk<����"S�RY�/��Y��(�"�q��#�ܿLõ�WP^cdD���D�X),� �`��g�+���('�0%d-��_`؟|	�.�&g�m<an���f��}��d�}A)������1}�5G�,ܦ�p��i]>��Pz��c�\�`e�/@��J3��~G��P�[�������,�dX������tZ��zn1L��{�Cϯ�׵� D��L᪉E4@��0(��7�ڸ�g���oǽ�|��O3�6�ٴ��e���2ȫ���* ��n���:��ҵ����!-�jzˎ�l�����.����	������q��e�1��,G$��Ѱ,�R�^��A5�_�[�hު�>s��tZe��1AW���HҲ��.��~�n��F&K��-ݥVæd+�A�1_zRq��`O�q�ơ��<Y���E��ی�kjz�*hz��5�a�sE��� ��h��I=���rF�S%�ý��;�cs���dR��r�����$���w���Sk�׺:����������
ʺ�e�H�-ƴ\���3��I��a�:$��p��l�)����Q[�A4�
���w"l��n*1�N?]��P�ɨ��bu~�?v���-�V>�%�$߹�|R�&(�P�}X$[[Ŗ�M)'�ڄ "�ف|-�k�)z���KNz\�s-J�76�rl}Cj�"f�r�k+U�����~+nY�rĪai*��D��f@>l��-7e���m�b3��r���Q����z�:��Iס �_9�77���g�o��C��aӗ�!�o�� =�hmS�A��*�ֈ�;L��� ��$�Dj�Eu�5Eu�M#a₸1���D�u�6M�����k`�>�`��\4h'�
��m��L��!	.�V�Ǻ����-���u\�c�ͬ|:�_>a�y�gW$��BG�>R_.A��uQ�qW��HЈJ@���V^9X9n'��(�'���OQ���9�98�[�aȢ�N��3u��I��J��lQ�H��SQ?/�k�9��%�r_4XAh�Щ�3kS3�����~?0�zl�'�Q��}g�I��8���j�x~e߾�=;-�l��p<$og��Z�J/jG(����*Qn���b����l�;�����@��Uf���>�W��3�>&uaAwQ�� �:n����1�J��h(�UQs��V{�"�W�ǩ�J(��P��S�W�v�'P�����$�ۚ_�R۳�d����&���8��%�A�A�����w�5)��s���Z{4W4c�V� ���O���/mA�E�ՐIN��%���gr�2��V� ���c��Z��7-�)_���[MU�Z��P_��	ڲ��{����g:���;�7-^A=��Q<�$��ienB��8,8'��|�Q��)�E�JF!�Oc��,�A�r��s�kؖ���M����5�Y�;��z5"l|�)Hҙ��sb:��S�����N�}3�w���H�E�b%���0`�f���ul����@�����F�����v�%b�{���m�hUn(�r���ׄ�"(��1K�>���-c,���r]^"� �[�N۷1y{}1��2cv�3�@��>�G���OK�z���G�(�a@4�j	�XHָ� �"�:��'���U���n�������0���E�#�dh��}�����aeQ�%�ywBz�;v��9/5��y����9�yQ2`Q����9��`0���l�xk��~�^B�P}d�6��0Kt� ��
�x�Hd��F�9��a��iO	lѯ�8���CD�v�	-��p��0C뮇�0�ݵ�\sot�S5����K�	��<V�,*x' �<J�� ��p��ˣ�bJ�jlK3;�s���?%����[��n�+`�����+�3ej�8O`��H�mY�%�X喿SI���:VA���d�j����u*f0Tg��S;��v�����FUl�#y�R��1���'sg��[2��b)��.�l�� cD�W�p4	�#6��	`ws�![^3�1s���}1�������\�I#QL���RO�����}���&Q����d
���M��" �d� �;��l�������
�E�PwC;g�a��8�� �zxq����O8�Q�&%�&��N~�����/ȝ�K�A�:f�ϋ�)��c�+Ail�Ǎb�nv�F@�M�#�PS_wjI�^<t(e�~zE��n��Kl�5��te���g���<��;�'6Ѷd�3қ���<?���O���V��D�и�Ƭ����E/����:�-e�weۓ��d��Y��fX���!�$��'�rZ�?s7��'b����Lq+Q���!�{_�����Jʲղ���%0�u����2�4�
Mb� C'C��KΙ �+���
p�*�B�V�(CR���mm���.O)��C�Պ̽x��T�e���=B���6�r��1��ء��^b�3�Lp���7�>?�t���1�{9xИ��;s���<BmLbQ?�q��V�����?	�o<Vq�N�	�YC	�5%�����a��V��V*|�+�9�<}* H��Xo+���0f����\׾�V�L��[E7.������YA5&nM�������{g2��?$Lh��*��&gӮv�����o\%7�)Z��o�H��U?�N���BH����!Gv��B��ӥץ�e[�A_!�U���EU���dmw���D~�޴剄A��5�]ֹ���������ľ��^�{����Tf�w���U�HT`�� B[4�Q�\�S�|���d�M?[�A��b�p��d�)�;P�����c�k���Å���g/h��H;-^rC-����eAʹ��(M6~B�L�>kDP�e�0��NJ v�����]~�d$��|��,�X��)C��Z@Kx�DK%Ec������`�P��j�?�z�=�؇<�$������~�A�^���� "P_o��A]�����N�4�'�[��M��(z������:�@w�5햠l��5�u���'���'�=��>=��_h�A�4ؽ���Ȩ+H�lW��yن�� %�թN=��E. �P� ���p�[���h̉t�՗]F�^�^Fa����o2�d\0Α,��ly�h�YΒ8�법24]+����f�N����Y� ����>�X�˨�^ڬ¡mB�>BK��mAS�S�qc�G�-]k�(��5����D�z��G��@݁��E�)�.hy�'���8	����O\��<~&D��qZ=��	��n~	�a<p�e�v�s'��E�@��F�n�Y	�M�NjG�����4r_H�����P�vi	nU��%�]�� �w�����U�����x
�Zm�YXł֎��ldb ����o�Ch0�5�ܔ�\��BU���ď@+�/��@�F�4���Ԛ��s#
Bn*L;����TDi�,���h�<�8`�g9�f��s�������xy{d�[�������(�k]!)C�lQ�:����C5�$[GK�͓g����BmuٵS���m�����ɬ+����uh����W���y�{�g��S�H~�-C���$����ö�F�@�� QN���H-��@@v���mLK���:�?(��y�K�+!��䁪�>�9ԧH���$ �Pw��779MD�������T�xk{|�[k}�eq@g!*^Zp�,���W�i�d�,!ߍ�J��{�&F�p�ݚ��mǕ��5�LS����i��B��c��Ϙ����RS�ޠ�g���A�����h~��LŮ�=�p㗵�@q�smK�٣�l�W����'��,�0L�8��Q(XL��T�s�E���f���D۳�CsK\�o$��#�y��s��E.�?q����J��9&�\����|��_����M�$��ఎn�J�@oJ׬�0�|������O�#�?/rH����0uI"�@+�����O[��J����o��'U�V��[w��8��'�����:�$�٠Wk8@-Ɇ���B��[t(��E,�˳y�aVv�6�JV��_�� P��``�S��o-� �5�2���S�� ���$R�	��ą����H�^p��#�i��@��ܤ0��`�̆u���y�ڣ◖)����V�_v�=��r�F��q�R\\;SLC
���~^N���ԯ��78� �H��犷��"Ɠjq����oP[!��޶�S�u�v��Ӧ�"��Q��L��p�UN�O���}k���+5.*�O����ū_e���#0�,hH����"��9��28R�sF���)y���3..��-�K{�:8fly$�Ͼ�!x��`�����6*p
��☫� dG�f��B1aNb+eM4���Bɩ��5�f#l��̐��K�l(Q��ۈ��\�.�C��|.����L*����2��;�#�=���-֧���$�tm��=타��5��R+�8*@=���#O(��^����vh A*S��I��������)vS05�dm�4~�>C�~��A�<�!���ust}H^�-8
�GH�\#*&��c�ػ )"`�����!�ɥ1��`��T|�ܹ-DF��'�h�ń�����s_Ub�V�_�-�y@Q��p'r(��O�����Znx����R|����<�\}y��	���\9��q@�vTT'D��T�s)��a�|͟�sڠؖ 5,bQ�{>GQ��{��5��W���`�Zm3�X��Ȑu!z����y#c�= ���*���Ϭr"�yyu�YK���IU6�Fy{�.9/�A-~�43!�SX���Xҗ�@) a�I�=����I�����j{����n��D�t�Ѽ�k'Q�!���A5d(����J��wy��ʂ��Pb����d����b����A���@7"�|vz���(�+���p�=Y#lYYn'_��&���f�p�":S�d����(��h���A�J��p�;�ͽ�3@��s��1�9�Vl��?���N��,]���x%��4ו� �9�<�|-,�i����0 ��5��)�˾%G�����ԁ���D��`�ۅ)d.��r��m)�{�x])^�ƲJ�e\��T��TԱݔ�T7((�b�啕�O6�Pƛ��J�`�~�x���t+�0X<e��%���P���_2ZŧW��|W���m1��(���Q�Ԥ���|c�)�{&�f�1�ii��F�����,��tA���Y��_�}>*��X��gP�qg��7W~�jV}�θ���-'t`��.ٕ�&�ל�(�䢷�\H�q%IF�g�d�0��	���m�a�E�J������qNM�_���yw�QPt�
�	�p˻����'���bTiSi��D�Z��&��!H��ۘ-6|�5�+ʮ�M��+Yx����݌�OܲT���k�Gr�Gi�ќ���%Kf���h�k~θ���`��Vo{�4Xħ|<��lqU>��n(�F��hD<_��{���y?üY#����Q�a_@{���I���><��{WF�]��8��̣YC8�ő$y�<�C��!+�}p��hޕ}�?-z�F2x�E�r�j��k q��G�+���}7g�u>�����\�"D�,��&(TY��;�j_
T�x<Hw����Q���g��F��u�H{׻&
��:�tdB^���΂�(��u�f��rȴ���b�۶�cM)fD�ɥM�Г�yO�^v�>����]�Ư7�Y�_O��gb�g���Qq�h���A�l��27�gh|U���Ar�`4vG�ZW��aT�e��!?B��I����P��c��.�sԣPz#s0��=�b):�glb������^
E�xډ�iP=ID6�"u6_�v�4`��3�b��i+�8Ԥ���k��4w��Øo�i����ڗ�V�ʰ<Z��]���ൢ���疬�W��f)F"���R	����Kh�W'�J���)�R���	�}/(��v������a?��y��`��G<h�&��b�>���~�c�W3����R�GD�G��}J{�,�:����|�C*�
	��%��{��WB�M�j[�OH������%b UKnG�M<"�u�/b��V	�-�������/ܹQ��T���V1e�Ѣb;0�C�����	o�EJ����M��2�ʚM�L��zVB��Z�^��Q �5����������n��K�����1�r�����=YuI2�/���2�/Ȝ��7�l0��17��8l��(!냠�8�n@B�~��\�խA��%ȧ�~�C��ѺPg���w^`��3�wf��L �����
����M�1UAM@/�_��1��k$CN��댆IUԚ��1��5Ct��S��뿺��)b�ȝ�TFM�s�g-Q�O��x ,RBx�=��Yv�������$��Ys��[�&�J����I��Z/�8��_�쪺n;�b�����~�-�q�%�'WEm������dQ!��36z�p��f���	@�;�m�j�bɍwD��8p`�B�CʕB�Q�1�c$��e7�<703)�O�Ȩ�J�UD�j�*n��d6�C�5W��Ջ�Bn{��n�|����{��¬�\&6�I�A��$-wZ%����V�]���g��c��'�lTΖ�ؼЯō��VMl����=^K����b7iI���>� h	�aI�s���mS��v�.	;VX����� 1K���{��;%��[Y��bd�;��|�*�WH��c�4	\�\�O��w�q��Xе�	Y:���`g��қ�J#h���1��l�^s'����c�u�J�;Ȁ8WNp���,�;��:J�qx� �V<Fq⟯�l,ME(�|��B�t/*�Ҳ �	f�KV6�,@�C�Ow�k���EV��緯��8�Ew����
cA��FoQ�>�b��X�&����Uh ��(Te�#���QaE8WRd3�@�GU�L,z�� ��+�j�(�0�ߕ�t��[]V�n�|d������10����5bX�Ӕ/c����Psz�,��^|C�kl��&|b�$��1���K�q�׏'n��Hx@�=O"�4K����n���Ŏ|��,4w�_ڱl�R�	뻳3�ZE����lz,��K_yN���pAꖭlIs��B�'��i5lbg��8���P�	u���=y����hPZ�ۖ��ε��>��x�s��;���-?�9xia�r��p���N��i���I��2���C��`TviݟRSO�Qfpip	h\�γ�i���^���%A��Q�'&���W�|'��44��Ct���o�i+u����(Sܧ�I�3^�%�
�Z��A[l	��9vA�A5 A� ��w�	��9��h���rT�ِ�rԭ=	W��5�hH�7��l��E���clz�B@�πd�[�3�8=;x��)Cj�^� C���m�?/�ᩉQ'g+D�Ш�|�ĲKո�eZ[��~*5F���PU�tt'�Eo���l3��Jњ����N��N�wCT.��/K�U��w˭�'�.�&�oЂ0�/(�i��w
��������*nBX�=0�����3Y�O��B����do�S�*Șɉo����T�XD�{h���-u��u"��}�bQ��M��j%<V��E����T+�\����R�����`]��~�t�-�n�]��Y
�u�)�OT�H��Ec�<��j�俧���~U3ՠ��[�ȷ�j-�� 0�w�H䃛����/f{̰�m�"O �� ʹ��R|9�rC:^Ю�Y���E��F/�qz-��̺���
U
E���ue�jL̥I���k�4����ߺ��e���>*#� ��{� �l�h~���>�c�K.)�B�����6�J��b#P
���AI��>QyO�.�9;�4�V��qI�?(�I��b{5|zm���!w#?��A z,0e��J�Bj	���A�Cf2���+]�%>��P�r73��jϖ���f���=$���g�4dy�
\<������O?я�'<���
���_�.�(;@��O���xDJ���.q�t4V���(y����B�m=��Z�Ī,%ղ�R+"J�ý�m���"B���d� �\�� ��->�����k�:�k�L.���i`�ѡ|���:����;��8Ɠ,x�@%�]��ЕX�[��%�ǔ�^��1��4�;)X��ι�zz�7�{Ҵ�t)�g��9`MZ;���Y�k=h�K�"��H~����]��W�k#b ��r_/酩�=���c?��2���x��C� ꝑ�,e�L"�>�ȟo�e�fyĚ�7�g-m凜�#M�ncD\�(R�۩��-'��yL���#����������.7�}��j���$��#Bh��I��eBG.�x#A��鯑�]a��5ȦC�5gj����7�r�Tt���;�^hwi�^Al�(A��+	cZ�J�����%�O�aG�|���ru��(��
4�B�@b��6FʸBN��~�5q4�K�c d��P�8����xҡ���nx��/�Y�gF&�N<L0�u*��M����z�Q���r��	�/���4="��b+�(u�����u$�����M���6@�س������[7Y��UI�5���.:���ǁ����wi���ڃܩ`G����~�[C�y�sJsq�:3�;�b�k�G��23�1���T����N�X��(�2�4���J�#2�G3��w��q�!%g.e�̋�PPh N�tAv-n�sf}�F���?�0�5����')���p�,��������z*d�
U�k�V�жS���<��ziSP�ZAS �y]5�����Κ3�V������̄O�Q�?�䆮ԓ���OP-Z���\O')���q�TflB��v&6������[��H���>" ���1�*'MQ}�j�e}v���b�@�'C�i����c	�--\�Mnfa�#�g!�r���Ρ��^�b�j�������ǜ�}|�y�j���0P�����;TE�=�x��p'�����t�]��]��yя;u+JKQH�I:.��͗�Є��\K7������4[�����k)=�L��t�����\��̊��5����p�+��o;����3�|�����Y�U���Ŵ	�fn�d3O{ۛ.ݞ#]��3Ѐc2���5�r[���}h�`�=��?��	P�l����%��Q��,lk�u��O٠���Խ/6�R* �����E3�u�B#?v0b��VȪ�b_m="��S�����Q���s�}���$�O)�����}@����{@���$�7�s��_�y�7{+�]�r�~B���{�5�B7�:�.���d�|y|J��.�(��eJ�iJ�L񮈋�2��/��� %ׯ�Џ�5�*#5�}5}��=X�q{�M��SҤa��Ϙ��$^� \�0��0��38\/�x�C�&��v�����T�(����/��Vu:�TF��q��9PE*��?X�]�j�k ��_�()A8G�\ ��C*(Vڑ��	�#�7�(�Rs?����E�?�@J�!�WU��;~�}�<ylU`?�ӭo<̕�M,�3>�]��H\��h���g+�G��z� 옞���Ś���	)I%�[}�����Ff�$�[�5�W>`""}ա�D�|,� ��dYl���������*U�J�G���'�!�W���s����KNՈb�z��W� �zmx8���9�$�
^�������:���X��n8՛�H�n������.ko�= ]H6	�;`�sR
���-����BW2���*Oٻ�Q���,�8��͆���������q�E�����&���p��u}���eXEe ��r)����;IQ�.��!	.@G�`�]��S���#� ��Gi��S�t."�P4;��5�u[ο���2�V�>���RMiS��V�M�l��6�58�^���Q�{��b��P�N�}]t�<=�+=Y.w��<�3�Jv��q��b=��B�g؏I.d���7����6�[C�]�[x��O`��7F��
U�	Q�eK�A��77�~�Ý9M�w�i.��8Ɂ���`�D��6�㗾h�1��D�yZ���`LQ�F�?���$��U�;��{8�g��fTe���yp��H�9'jFIB��-e���l�7�qo�6���	_��A��T���U�*0F��9�؊�DS`�2{��o����[y��x3t����j��ƾ#��/�\�����:��w�t � �K.�RK-�5�t$M��j��E�Ă���m;�d�N;W��ݲ���©j|N!���b�%�[��ie��`~�H���	R=�=���>M����)�2��d�H9�<��J[8l��T���FOp�w�y��,�a�/����>ۂV�Jԍ���w��G�Im׏��)$EKR���D�Ͽ�Q`Ҝ� P����F�<�x6�~��\�2�6-]�/&�&��/OS���CU֊���!�ԓ��Ѱ=Q����`���`q*FBh(�u�D�_~	d������L�0"ta��@�m2��`/d2��q��m!~�Kn
G�]��Ix.�9hjD��l#^j�F�<I�Gx 3G��}?���+�7�� 5TE8&����Y����~*񈶆SK,Z!�2�e�Cp`S�9v2��C�G��v��D2$�6��r+�|d�%�F쐗�_�`���9�N@a�M<�����T�p34��}�����x2��w[y����ı��l���s3�����$���<�x��Σ�k���j�k��6�����0>x���gm��a>w�{޿�Wb��RZ3�79d��0#�.,��i{�/'~ �
��zA7ZJ�'?�d��,x����;p��2c�A��/���z� �T���B&)�o��yA�B���|�,�@�ݎ��eiDѹQZA.�B�2S���:�1��c~����r�ܜm[�Q�j����U��2^�[�ȝ>�Z�ܟ]�hQR��N�%3��Yt`y�%�r�	����W�o_�W� �����&���x74�E�W��P�:�4_C�"�<�-�n�8��P雒�YYm�T=�A��S�P����D��t곛4M^��o�Ա�g�9�>���B��
�,0E���d�|}j��n	��_^���bB�*�>��c���<D9�Y8&u#<N9Υ���i�V`�W��!]��|�q4��*�2v8ݚu�č�$2*n�cs?�DK(��%n�"7{Z-����>-5tu�t����oCh#���a�P3�P�Φ�x�U�_�"s|����8�	���!qQ݃��R5I���K�С�׺y�Cp�8�,�XS��/���M
!��ӭ]dJO��%�}���8�/�'ʑ����3��'* 	�STG�u��@� ���Nݭ ���N1#�y��q�n����~�0�G�r�A�&�����bFqhb0?7(oe>�iW��k]�Q�������]��|����i���Q:%[��u~����W��.�&fӝ��[r�ˉ���@�J�v@l��SZ����Q#)����?$N������Q���A�a�-�z']5��丹|���o#d�tOx$t�¬�����A�|l'��C����Ǡ������r<������ui�w�{w⤍��3��(rI05_-2჌�o聾Ǌ� ߣ�f[������
��' ����$��>x�=A�K��-�gg����}5�`{���5�7�lڢК�!���|u����ٛ�E�^�uk�z/��>(v��%9��_�K��X�D���p��)��8�9[��?��~z�h�
�gl���-y�CVFY�Mf�-$L���ؗ0xNq�;ַCih�_G���n�de-�.2ɶ�}�>RuH�	*��b@���|w�d�c����\�_�}�@QS�;�=�r��0@�TH S��4� �.����޾c#�e)������57Ġ���I8p&�y�FR�+�\��m]SJ��]�{���71�+���	}q2@���8��p�6ٌ1�[p/�2�Vu\��i ��������`�NI�ʩ���ų��G���&�Azԩ�`K��p�ٟ�2�S�������-3���}���
�"B��ʑ� ��#==������E���^���t�C�L�����ew�Y�_��H�7KDiǎ#�5���͹O	,��Irh|�n���n�@�Nf�x�D/H4KYO1�}oqz �J�,ǐPf�`�My!^�Nr��m�w�Z�Qծ��a�&���杂29.C���1�v�>�n>���m3b3o�B�yN���=v�F��F��'���>�n����x	>_�xMm����GJ����n��p��p��A���Y/���6:��I�ZY�F-�@*�YY��qݥ �3Hk6�+��1�� �[��#��a8���\5:�Η3�V���K��P��6�ZQ�t�8-�ה@��zҍ$K����c�ҢAπѾV��}>:
��r=@��uc��T�M�2=�����%��u#�7��E�,/qP M2#W�R��Y��D�ԑ�:��](����r���z��(�1(!��&k�b����		��:'s�2Q�����
g��M�`Q��4pD}5LQ%+ï�_dq#}("x�r=�	Y�E�Ь���7�����Ĵ; u�Y�I����&��T��E��)k��}+`����������_���TԀZˮ�D
U
:�ŪJ�^m�Ǒ@�)����Y������~��},|�3��?�a�Q�q�ao�+N��KTfmB����&�����~�?�@��Z#���$y�ە0��SRh�o��^n.o��й�[���D&�[�io�=�Y��D��v�[��"��e����"��=�(�4��x���D�|��ܐ6�ml�"�g����ecD�~[�',UK�oM�u.m#i���S�E�ʵ��vX����A��=����4H�}t֜�k� h���
6}p�Jh�eq��A��/6�^!��ވ��� �t�P�cH'�[Ȼ��G�`�Eq����&`X8b�T8D��CKP�B�G��xn�>!����W�#˧�]t�
��O�l��m�d,��q�??c�1��FPV>s�$�۽k���B��&D�~T�͝��ف}�"U��h�V��! D�N���S��h�����Z�x9�0��|��1+����}��ْ����57b�a/���j܁����>*�3}+J%��q��O|!Ȝ�b�W�87}�7*���G��}\��~�gWI�T��Ӵ��s%Le�bF��0Uޗ�8�c�0��Z<�d#;��>�]��ۦ�r�^uj��Z�A�-a?�s�{'�Uxo����J܀���U�s�ԫ�Z
���m�����=�$�٪C�Lc��\Z�N��6{��:bk���U��!�keTP�yVmXA�&�����{�">B���_%�^Z�DgV�,��PL*���2���³zL��;l���0g]J����i�X���b�/�8�X�Z��׵.V�SɦS��φ��[0ͼ�����9;����{��l*��Đ�-�1	A��e�?]ǧ5r��r�/#YU�1���ݪ��Rl�� �=�`D�9�Xbl��HIU��u�.���e�@�S��ѵ;� ɍ"�gg{�$�8wFٍt[�g/���Wz�:0@(.��JU���F��6C)��z3�z�t0˨�:�0=L�wV����r��ElU}T��!���Y�Uoҹ �Ŝ ��vb�-������;C�2cT\*f�a�,�oԼ�UR��s³ے_]^U�4u�2��7՟�w&�n���$U���8�w��,���L"�=���P��@�����铗5a���{�]�+ М}�?���v_�scΥ�	��jCK����i���ҽ��+5<sr����嗕{n0�����0�Wݵ�����n�;���{]�_��:���61�i4���f�
������v>Ԩ.5#�x�`h �^���ؽP�7&�}e����_�����Gn\�W�7�
���^��ڛ�&t]:�q9"c���D��3\JAϸmL��aj�g8�Z�Շ}}!�ݺ��1�8�H���Ni+\IZ���ޕzH��@&�7�j�����
���u5�j��!�F�oB������y�.zv�(9��Gv2=��O���������R���^U���5a|�&<����c8��1��|r\%�22���͟7��M=��k�B���<��IE��ή��E���:X��
d��S	Q&�[H>��t�Z�;��?|���eņuiW�V�d7�3%�/��E��>�~x�%5�|[�_zHU,����U���%�;N]��?)�`�D�t	�0_�~�w�|k�JZY��b��0�X�St�Gf�
E�raec*��|�	�P8���Ue�j<!�׊���󋔠%�Çn�iѝ����9������t6����&i�wh��%���'&�sY6�-o�����D#��x~�_��Fm�Zu����L�O��Yk�9��pV�:}�@�:{���~��4�8m���A�Z.�zB�)$R�f�&>�I�LD�t�7fޖ&�<�z����a�h�8̦RL�ۢ�e>��_�$k���Gy]�f���	e���H����_�����~���M��9Ar�|<>}����/�eC��W���F���=-�K�d�L�Z��*�WS[6��2�B ��t���F�%Ɓv[޺��z�B���|hh������x<0`S�C8*��o�¬� �.N�WY�sB�=���G(�=��5�z�g����{�v� 5Q��� ��@(�Z%��+�GJ��ܠ�I��l�nO��C������U!��(d�ֹx�R��H���`��orK��>\��ƒvJw��1
��
e��}���I�+���zK����e16hM`�s$ҳ&,$0ny���Ͷ�{�;Fa�,l{Kj�Fef�������4`�lr
�"���a��M�Uq��.ӷr�r�C3 �vf@�i�$6��ʋ��,B^��кHf �E2e~���T����SՃ�e�a'l�|H���]&�|> B��r�����������L ����LIr՚��|1����Q�1WH���O���%�3BWW�L�x>3g0�Ub�/0�CZ�)���CI�s{y����'Gm����h���2����G�y.�稴��_��K�L-ˏ�m|��>��(����$�dR�r�RV*��֥�w�]��q�2ާ�����Km&�NV���o޴�K��������ȡ6?0��J��K����?z��R�B�
�8��"-���\AjۼuI[y��񏊀���ʣ��q;%�E5�{���-�	(ZA�8��hi���o�|hƶ�۟�B� ������a�A��&R��eT"l������N#s��-���-,̋
>�B<���gb���'��Jk]-�HR�Dbt[ ����F2�㴚��〄��	i�_|��(Ѣ/��A|�����qgL�n�C�S��7��	��'C�`zM^�`Od���|�Z�N�㚔�0�o�΋o�ya�;�m��/+k����.��F�~�A��`0���e�Eέ C����TSHr��H�Q5Ow��u\�2 ��Lz߷�K��H�)꾲Ф&�Dpc��9��o���C��$%\� ǿ�F=!��d]Zv�n�^����PL��',Vl�t�ȀSg��;����CV�j��[�C~�N�]��5@�
����7	svb���7_����u(�� �n*����8D�}r��߃6*�S���l||�0��������'y�\$e^�@��\�ؕ��;y��b��u��J�>vpUtF?��8��U��GG������f�7�\T�����$,^�b�4(3֦��6����8y�о8�����KN:�.�9~��U�k�V��	�_r���>�������G��D�v�r;�!�����{i����>Q�i�ZTp�0vt��}�*��8���T,�5�����KK�w���!���M{q ��x�����G��̐/�F�u��E-Ys. ��Q�����l�t $J�X����V'T���E���8�4��)9 ��0��R��`bjb~x<�͒fy5�KJx�Qd�1$��s�U���xF����Ts+��O={�5�|w�Y�[��K��?�[e³�fO���6&?�����\ %X�	Zj	����UF�`�:5eqn"�d���iǅ-�E�{�/�$����78*Fn����]�FI���ܝ�� �H�8���kG
������d�f������6�w�t�OA;Ϙ�2�j�{ePWIp´D/�l�j6Tǟ�����7���Q�^�4<3��A���p��70b��r=���,\����-w�h~g��4�jc�T4���5Im�Ш��b7��AR���mI��-���+m����`�{aǙ�@����p<�G�:_�qצ�j�S�:�ܘ�5���7��##[n��zc浲&�i�?)�)a��<�S�|C�P�o+?V�>J��+�/�޾�0}�ig��X[p!9.����n���`W�h�M����	��:�F��6���' |���=Q f���p���u����G��H�u��G����	 b�f�m�t��h;n��.���ԁ�Cԅ7�w%hD��4R�3^d���Hߔ���j<����i3�_@ު^�`�9z^��6jzy�V��.,;�oC%܀%��pqѶ�5�C����P�����K5�
����T$	R6UV�b�M1\v$t=�Q2b���sr�MQ���Yr`�]3b�g�xQ.�GU�/!�Ֆ|	�NuJG1R���I�ń/%	�J?�6S0V�.{��Ƌ��%��gd���;@89����g�p%��VG�LS&�i\�$#Z�b�2ȯ臷�(pm�E�1�W��WhE�096�ܮ�I~�`8D��,Nt�'[+�-�B��'�u	�#�=렻P����Vj[iq6h������ ̨�GS�����1�0N[��KihdYZ�R�n���-c�5ws����#���9ޡ#\�1/-�\\}�ZD����<�~��c�2�����>���V[_�͏���ˑ@���j��?��v��=��\̋�ޝ��;G���E�6��um�B���N�8d%R�;[{�Rlh���/����$(��"srj`5�I< vlS��.�a.� �I��v=�#y�_8�kl����!5��=>��U�7�B���O�RYy��1氚��AG��h�R�wM��¢z��� �+���ܠ����vKO�-�9uZ!Aw߇��v�m�d�ڟl����+��,��.y�7m����wP�c��c��%A�`N�8Aƈ�a�J�0�7yJLK+'���Jw�)�! ��I
J�'�m���^�%-�j�Irq�4�̉�g�J�����-�Dː�V4gY8}�}�w�lb�H��������@�I���[���v������]�#��(ϔv�%�!�hc:a�����V����(	M��E�nlv�h��~T;��6�7�m4��s.�����Lj�|�4���6slh�����%+\�\���Q�F?�݁�7FiҤ��ŝ�ׄu������;vS=�E���M���;�V�W�*H}�^�Gi`iTK���z���|��Њ�Jm�SPP��.��H�;B� ���������Kggyzl
��(e����������N�� 8F��.�2]w��)��H9����� +�t��~	"��s�8��^���__$�-u����ٙ��\	C�A��qo�������j��ܢ�[;X�4��>��`K+��%k[lF��GupI��@fa�D�1�9����h���3�K~\�\9��=c�­%$m�(2�����M�s�A�:p25��Q�[(�qq!ZVq?{:�ӴE5(֡�s9�� r��I�[M�K�圈h�A�w ��� :���?�@���<�#�d�T�)*m#� ���`j� GMs�4�!\�JH�c6�ޑiU���й�},��e)̺��
�V�}N�9��9�!|�1��b������%o�d���&������P!������R�-�l&�Qǣ�)�߽���_qL�����܈����4�-�{E8��l��r�ڞ�Ҫf��G�;b�F��޸yp
VC
�C��Z??���
 ��R���=M���]�o#�.��X'TX_L���_��?�*w��Y�k8 �^��Ԑx�V	Hg��)�A�y�$����yg���E��WC����4�~/�̾�<�ro�)�i��o]mk��D���mb�u�2�m�k%��Wn��k���,���/�X6<<{�������$>��h��x��ď�Z���Β�G�i�$�wgB,-��������c�����*�빩}�d������i����"bF�4�8 �(,�dkO\��!�m��0ҏ�PAV
�O�M����^�`l�(�VQ�����q���-�A1.oV7�K�ԢP]g�a�3�y��u!���t�l7���~w��M(�{j��	Sv�5�����D�{��B=̉��j����4:�e��*���G�B��y��u��u^��n��/�h�a�*ß­�1�F/ّF��
������i��E��u�����L�[Lӕ
��9�rAwџ7��,�����<�h"�w7�%Hm�K!��0�z���0c��W�wj��<W�Q�a�1�/L������W�q���W�z?�AP:yjr�ks���ꖓ��8xN�#8������@*��ӇFNE�)SH�N�T�����	B�[uH����U#��S�m�S�ܓ��OP�y�'Y��^�{f���h���ܔ��4���$rۈJ"�C|��:�����IF�xj�p-�O� ��a�����Ӽ׺��|��䠋S�[��N�s}g&~58Az���Sw��1.���A{��6EA�WyL��Q�D�9���K:���6�;���3�^�;�O64m�51:,P����.�q�a0'd�⸂^����0���*��\�%b�?Tݐ@?�)�Az�JK�2�#0��x�w�*=�7�Ĝ12�b���}��P~{��}����d믵�qkҷ�I�L�D��F���G^x}�����%�������7+$�+���^���+�P
��4C6�>��(����t���>&��u1�i���$��0i��4�o4�8�"���[���V5���Ch��~�(:�H��Xח����O�W<��g�F�P��=����U O�=I����\�w :�"����U�;����X6+���@-�q�t+t�m'IϜ�:8d�D1��,�ܸ^t��y�$D���~�biʱ��A�B�1>��v�r��y�P����E/�~�Ly�U�NĐ&�H����9 ����6Z����Q�������5�f���~������"��?��0��z&�C_�i[0��rZ��F�k�y����Y+�w�Ҵ�4�^a��bf�5g]�_�	�k���s������"����d��1Gy�yY�@��+ $d
Ǒ �L9rv.A����0c�T�����6�a?r��m �Y����W�ɩcJ���'����lJ��,.�tôZ|���꿲�)'MڸJ!�ˡ,�, }��Gn���ϻ��ٳ�'N�ֵ̼C��5�!�"
/C��V�i
.,���E���de!�EĬ�\x���D^�buz�Z����¥�I�?&�q�NA���N*��d�=*�|�@�.Q�WV��E7��(<Q6����.rK�#�]�y+�*oi��ƞew��!5��������1�`�=ʛ�A?/Ω�4�2\~�'I�oȴ� �9���q8d��$���3͊��~�b��cud����aT�U̖����`��-����o���_Q����Y�S6Ŷ���i��K��׺
����sO��D%����_�� �!%��iu��zh$\��� �@�%���~6W�,��{��k� ���z�|�l7)�0-���I��ۇ��,Icv!"(c�����MR�j���-���X݇�%ҝb{s�8��Ӗĥ%#؍i,oC��ן��{I������O@�)B�n.!T��eD9��Qצ����)���VS�$��n�
.}�� ������_7C	D�tV�t.��P JͿsV�w��\�!��0);�?d|�j��%44����w�͡S�]R�RP���@8�l2X����邮e�0T�핗`�\"���XW���k�_u6�� a�#����	t�R��5r8�C���h�������ϔ	�IS�+ޫz��[�E�f����D�S9Kׂ�|���`��VF�|��R�+��(,���(g�5��մ�;����ipo�����럊%�w�u|��\Z�M�J�m���Xq�1�r)���!�����̰Y�53����sWh��S8���N�i����Jd�V����q'��u�(�Ce<+�+���7a������!�� ��e{�&�P��;:	�����Cah��[�cn����},�w��Kda�|�h��MB.�����=�'���{��Fh�Ac������@��c����SbߍM҆�@t��R�i\`&t_2,@��`�%��h��H�x'1��
��}Ed�9�����.RP�hEqgt�b��;�����7�,�6�H@��b�Q�"������VvT/~��Ӥ��+��RQ���_ْ\�"r�g;���rf����7��i�&Q4a�R� M��L��_��G�8��[J^RZ���1�)���ȼ9M�54����[R�O> ��=��AE� �Q;s�"�N+U�P���}(V{K7�[�R[qG�@�&��{�6e�V���hMlv5�qFH
tCyܫ�%72|x/=
t*�J_\ ����"��L�'�Nd=�+[��<�������M�Ȭ������7��36?Bb-���$�%�pq���Xƾ LՆh7�~��z����Q��hF��̧w�E��=*.sOR/H�������Б֮���G�B���-ȮV����<B�IЊ��c���4���l�t�����[s���:CՅ�hЙ�t����D3]�A�5!�	T.�?�*UDu��Rժ�� [&��'yn����ͭ>{�O���{�?fM�z�A��5M�<�v*�8�\�G&V��8j��Y&�+~8�� QH� �@������p�צ�L��X�8��^��f�;�}������ʤ�G�)(CyһNw�D�լ�����^�n�T��:�	Ƙu(O�2L���9������#�
󅛂?�&6�,1-{�F�\��c�k���l�U��S|
���J'�)�5���)�ac�-"I�Tm<U1J}'���s��q��O�ݔs����m�DcҗF���#��,�H�s˕�t�;hB���b ��7}A��8a<���'?R������� H]���?��K��AH{l��7ۮo����g�f?��guݺ�w�\�v�6�������p��vXV@� ���{k�mt��� w�1z@<ٟ�<�L0Ѱ���X����h���;ׯ܉/b��h������?ߙm�+�� f�5��yn�LwP�<`�Y��������tE���s}Ĕ�u[�WU�d���*"��2��)6#<�ct&��'Vbz�łm{�aMgƃթ�yg��x�>X��
BAʮz �&r����0,Na�rwK�`��l�\/�EJ�UE��g~XM��	S�{n�wC{�/T�ݒ���b����Fg��j~����Fڵ��G�s�"��9��,���N<���'��_�(��I�5���h�Z���xؽ�=�
��U%�L�q�P���_r�S��2���{jh�d:��̹���t(H����s>뱧2UzG��l�'��|>oA)#|dc-Fn����h���/�o�=��,���]^�r�'&�����7��m����J�tY#�֣������h
{~�[`�*Q���`��W�W�e�bq���pg)��`
 �yׂ
�}�
��a@LǄ�]�e�T�/��!�q�����\,�ێ�i�	��OE� ��i���y[�L&R"��f?9�`��uG���Ǖ2�_�x&�-�hhe8���}��1�<u �O��� \��Z�ٿx�vQ����>;3��zE������s6�[��:��#��˽q.�#�)%N	Z���<�������R�'�`r��u��b�}�[�jX�[�G���Ӟ�>�u�6W����|Tu,X���ʔ8yK�.�dĦȀm/��q��i��u�H	؇Қ@�f�u�1���Oo����'�v-������$�s�M�c��Y{D!�-A�9K:�P;A�!+A�4��n������+�}%��b�|�	6A/tڶ�Z���ᛞ�h�Db�~��
��DY�FUe[j1D��d��������3�x�-C��(�0�=H�Q_�d@Nz�7�Ѽ�Љ;o#�i�qP�r��>iL��5=��'y�	x����Y6�I�2W7��0��r #�i�bk$H���t�N�B�qBˑݣ�^�cQ���c��X�'i�4ɦ#'�	dy�;�N6-Z�G�^Ps��$ qX��S=�1�<ߕd֪/>^B^m�Eݚ���ix�?�] J���\�/-�/`i���j~���ס��}�_��I�Hb�~\Z�^�3�DX�E��%ѿF����DK��L����
�������O����-J^f|!�L~�aY��\>A{�j��NS�pCj�0W�Q�Ȓh(��:F!^�A���&(C@�
��O�F�.H��/��J43��5EVqw'撅���7-Y	-��xp`;�5�����J�MǊ�[jr���3o�R`�����ڢ��=@��E�V���B@Y��7��N��*_a�OH�D����OL��4�x��(�3]�@v���4K�5����,��krA@�ʯ��~��zWG�YrC-��g��f-Vms\�Q{ 2�Q:����Y��8d}+�m&�ů��>h����0�Xϴ��9�ݒ��f�a�U����z��%����'�}c�\n��� �O���D����(,kMBG����$��W�3ك�	Yl� ª;��9�z�s�gS���|��A'{�OM�nmQYOnbͱ�8]|΅p"l�3�+lQ$w��PP$O3^�Ќ�5؝� 9-缴o�YH;M��DRn��J��J�~jN��҅3��&k���+Kjɾ�'����W���c�[o���Ɵ���p�!���]����d1NsÙ��N��xo,�"� �/�h�'��X����^��Ⱦ���[��q<g����?�0��K˝�ԅ�1�Pĺ����baБ'�.o�8��.��(,�_y!��Y �Ao����U���W�gА���e��R\����n��!k+��dxi���#JrD��@Qe����C����X������8�Wk�c�. \�%S�\�ƞ���z΃�`w�~T�F뾥@i��ӥ��O:��j���c�`��l���+����͚{2�I1�_}?�}F�+:`��ŏeC@/�Fß�$,���_�3t��sj�ˑ���Փ�Y9(�{�`j��W ᢖ�h�P.	{	{3�|���1� ���ڜؔ�c���1�\�J:{`��?��E���hKe��6-ev�K�ys��R"����K:Q�\���n��Sg��td^KZna5������7/]++uc��Ѥ�o[��%���ʂ�=wťh�&CxN�<K��f�U�tRk#��{���v�)'�����t��!t5���]&��[��E!Q�;�;�]�����uz��>���opŖk��#."��4��T������>��tS��S�Q���8����[��	|s���<�˵��޳O�;+���'�A�񵵾	��I���X����+�*w\�ʥ�6v�F�	��Ql��N���)r�_���C� ��W�2�(�s��s��:_O��'_�ZR���k��j�Z,Z��w���R"�*����ݛp���E�X�H~\0A��/���9X�;?�z�z�0��cZ���q���z������u�d&�XP!Nw��XLDv~q�<��L?[�?�N��U�'�4q�r�Dan�Q	3j �1�
)C`D�:"��<��ZQ�Y�,/�l��[�n�o�^3���)�~ր�~�k��b��VSp�|�m�����tR�|����뤮�ե��x�ɓZ���1�#?�����]}�0t���YNG-1_��d���+H� ���*�9��p0b#�H��G����V�UO��X�W���B9�����Ze�j��19'UMҖ�3�gՖ���t>Ș.�E�C��~��`���LuӋo'6:T>�NT{P�_'�3o ��!#��`��U�ԓ�}��*��T�V�Ҳ��D�!@�Y�b�s�퉒��������5o�-��5uiqEn���&�M�lG�K��"g�By8>UVA�07k�����a�MH����2������ͭ�,?<���u��'��b<
�I��"��sP���D�����s��2B�KWS����!��'I`V䆎v�����q	�Z��׿���|����Ή��(�(R-Ǆ�x'"�
ʹ���H����yn0�X��ia�G��R*�7Z*l�ݎ�]�uk|�h�����aZ�V)]�S���iR3(��XVV'Q>8�v�����7��t�r���hv�rTP7�9 .~�l��mK����v`Upg��͢�r��)b�Ͼ,�o�m���'P�vU���	�>��Ħq�z/��#R{`���h,.@�z���G=�h��B��f�xh��^%���>��1�Pf�x���ev�k����RLBL���u�h
�����J�Vr��cLs��Z�`�u)��^d�Pxc���JU�cxE澻4�E�t�6Xi�H�����q�4�%�
�6n���S�lWUԊ^��(�nF�U��7c:����p���̎Y�I_T�~��>��"�8�f�^�=�+D%�����J���Y�q���gM9�G��v������A��>'Q��\�hNI_j��;�K���h�6��2�^fG�`KK�)�F�jI��bW���Ҡ'�S��`tΫ�Q�'���*��;��YZU�k�'���tW�|6�h��<����x-^���ɣ�	7h&�>u��}gԱ~�����9�g�3R0��r�.��niSŚ;\k���U�&�E�3|�=E
pm���v���|h�^)��oo�����E�қ�������u�*���{�|���H[-!ȳ�bĴӒ'S}�I���u���+��@����0	�Yj%8O?;3,�f��q�9-�5 zdƒ{�i�r׹��U��������e�xZ�φ���$Ǒ��m^���T^�"y:el�����_�I}�)�K�sm����ԯ&�N�iȳB,j�:����v�Q;�4��J���M�S����Jsd��=HIQ|iϝ��'�n%t��ڣs�"FD�
FY��|�@��B2�Zf��|�r���G�_:dZK��W����,��p��(��G��m��&9dv�+W��r��-�YT���@{�9�����,i��`
��RL��{<_%�z.��hQK�3r���$��Y��\�@6�u�ήf�����X�2039hh���6�� i��n֠ΛC�Rt�d.��L�}*,m����GzI��*+��Cwݢ(��%�fYA��{�����q����S���|O�����Dp�t
*�?�Tؙ���f�kC
zZ¡�%ʝI��MQ��"�"�	L
��*��i�D+~=��`TWNC�HC�9���R����N鵹�kf�dA*mD@S8�\��M���r�ǳ�b�����nӎ�]���u�=�<l�륜�0���G']��L��x+�вZba����V�R,��
���+m.]A/��K�"v�R.�R��OS�����3�=#Z��r�Z��o{CL[�αwP��b$���<qWVB�C��LW�Z?��W�W��;~+I��j�m'�j+�X �GGOd�_P�����?��?[
�����^ӽL�q7[��X ËlJ���RNȻ���8N6Y�o዁�4�c���ڊ�._p�5��iQ�n�w�ϴJ���>xJ�R��6 D�bp$M���,�qЇi��� ��$f1b��H��oGU�տ?�\HI�A� zc���\B��l�݃���v���[�e/!���]��7[MLZ&q7�[L�`�nH���i����:��P PA[O���&>ìp�­vu�NoQ����,[�����+�� 3�Y�Ȩ�~<��%�)�-5���jΩ.$7����l~b��ox)k��qI�#��@�m��9J����_U3>���x�Ƨ��;�ا	�3��,o�d@��� kl	]�����*�b�g��=�ʢ����Li��U�'�}��㉢�z��6���DF10���>h4<�$]B'Z�I95�n������Q7��֘�y甃� s����n2@�G+hS�W��X�n�W��r�3�:�������5�שׂw 6o�!�$�q1�����}F���3vw$:�����>lrB���^���[dU=����zS��;��:m���g됏�![�R�*�5̣�&��{uТ$w�Z1Q5˳�]  >�lC��CAb9� &�R��}�˹/�RҼuGY������ؘy=TA'\_������P	�$6u��{ ;��~��u�,��F�ƙ����.�E���������n�Vf#��70��g�d��%~���������Gq�]�� ��O'?7(��7�(��w���7�����Aq��rv��e���ʮ��� �ΐ�����/eDM4H����Gө�S�V�7,7ͭ����H��Qg�7���-��+A/���`TߪI~�]�	�bo�`�_�q�ݧ�	��k�V�۩����� yt{]�C�LW�&���K?�5	K�/�)���V�Gu�����j6���j���~�̵\\��:��ֵ�:'
(g,��e0���tLĹ�i����)��P�(�IPؤr�r�5�a��5����=�Vr�OK�4�ޥ
`}�&��BW��%9�$�HN	�ϢY�2�R:�fl�Bx*eSS�b���ʺ�aY��gU�Ƿ-U�R����VkY2�R�W2J+�N;&هa&2AL�͘��I��">�ܸ=����<vv�K#����-��O5׫�e��7f o��	P��n_�Y��L{�ȵ�)���J�縝(Ƿo,��%�.)P�V�qa�4������D*`d)��ړ�۾;z���~�h8�yk;�\ı�1�*2�yt[�;7����~��G �&�j��@6nQe��`/���9&)��{]1�r��j�>��3R)	P��BB`�a�d���B5��43��v�.h�F~�k��tA<�d14vxI�/�ju��G�����OJ�\{��j
��]Ob�_bjA)�pIos�5J�D�4.��ļ���'4m��ιBo�!�@�v��W048+�+�AO lR0����\z;�ˬ����ki�@ZJ��p�����K�Y�L�aw N[����_�hx�˹�t %eI���َ�mFg"��R�\/Ő���P�J�T��	��w�K��W&f��?��.��87{2[��ٺ�����>��e�J �]Lp7�6Yݓݟ1;D:��&'=�Á�/%4�M��2(WX�[խWȭ������mi���}�.����?����0���ھLtz�S�D��WEuG�\���sAN��"Z�:V���z"i:I�<@@D�|�M�X����̮V�/�dv������O��w��˲��pk��X��gX�:�?����H�{�^r����$�f�+�v0X���E��e����J	d�Z�IK�	�׼�S2�]�Y���o�I��I�Z���z�,`����䊳[�9!F�t�w���1U����K����1F�-a����4��JĻ(C3E��A[�gא_u8��2�
[�Yl��fϜ`����=ӂ�̕1�gZ��R�
�$(��9{izmR</�2������UZ�u�(��M ԃ��%O�Y��Y~���Hy��ի���6��N��Ά��]�ݭ�6��.요�
��(}y��|���U"%Qr?Z�H�	 |��?$��Rr��l%�9��^	�2�l���]M���@�`2�����ԡ|��Nyc���6
q�R*~�S7��؆^~�d�A��4�d�`Ew[ %N��j�7\�!W!fJaro�D9�����Rc��0f�PA��t��},����1!�^��񊟎P�.�A"�1�g��|r�cq����rհ�qw�훈�ӫ@d[����^��<J��}�X��Rk�g�P_��Ҽ
Uw@��v��8'���%�¬�3R/�����+%�o�t���A�]�m�y;��>��O�W�G h,R�!���v���-�t[�}B��z苊iR&�(��ךXT� ȢPA_}�c���b�V��,��y΍�a)Ht� �E䷲����+ڤѡ��i�1�h[RF���8nb6d�����09���{|@���E���0#�Nφ"%�*�{~�a|Ѐ5����=��9G)}r����ti�ϰb�w��Pb�،��{}�&��ߘEbqs��;�����1�i�Ed[���Y!\�qƾ=��'X��?�X����'����TV�W<`����&ME}ᄜG����r��?�(�vB���G��E��X ���^�c3Q\\��Y�y|2x�j�h�ʐ*�B��V��}5�4��.����+@����e *x-s�d%���E�K�W1����������g��)���~ޟΝ�%���'ǩx�A�X����yu��S���\�v^zs9�J{�Li�E�D1k�c�(C]��v'���;��h�,9�[~S|����3�弡�-��y"�s���/�oI+؆Te�C��>�ʞ���r���{yr�k�!�"�) ]�S:f�kd��-T��_�����"C"�t9�C����[�B���8#����2�fKJ�W�>qL���3�m
���\�%ueNӶ����a!d��~���8�a3aD;L�7�8y��~��(���C��zv�[������Q�Li�_��*3��G�2.`�GW	_� E�7���b+���ǥ��{�PXHB���j�߭V��/����S�����u)�J����D7�A��-�0�1GZYn��m�J~hoL\��[��6|���S��Ы"�zN[4e3=�����m=�e[=e(��!�X�}]h�3o9h�kX8���iPg@@�"��K��	�Q"P��G
� ��&��p�X�X�4�w��PD�y��,)&�OMh��U���%���i�)ծ����L��ME �S�7��[z�U�^W@S�#lGbu;K�l������w�𧻓u�#�q��:PP"t[O��R`�i~[Qї��þZu�"���\��=���p:����� �Yє<����7��0�by��p[yc%�-Ē<Z?���|����e�N20�|����!U0-s��'��0���ɇ�,}=M��tq�?�r}U����,p�6|�h�]�^�\cm{�ט؞D�UZ����K�fJ��}�Pi=P�z_�Z�
�
H ���fcxÀ�rG��&L�w�������%r�E�G��cUb�J��A���bz� ��<��I�6�F^���� TR-�7�61k@m��(Y�6���ک����Ih[��5�4A�B���ɜ�ӝ���`�Rq�趜���.�=���k��YQI�6`����G�g�`�_����_��3�>�\�,i_���^�T�=04��G��[x w�Q��le��"��u�M��Fr	2D�П`����z��{���[�dU.�^�W!_*��=�r9�>��ގ�]7��uH�ٶ�K,�h6{xl� ӵ� ���U	Ve }h�
J��rN`n��]$�
=mN�˔�
�]��$������z��"�x�L���Im��_���N��1�7�
���%>G�X��jU���I�_MJw�����0
����@�T���w��8��֗�����$40k�s����DU&��N���2��+�6)��5�f\/�-���r�V�8@��S�^,?���6����=s�$긱�_R��G����A]9]�.(&=#���8�j;��������_bkN���-M��8�R�T�a������o�N�iu�A�*a4���l�>XT�Z
�oK�OSF��\�ti�@�����kq4�M)��N~�|��e�H� �lXe��XW̲���@�r'��4��j/晟N���M�v2�SGA�񭺻<��F�B�����>�`j�%�7�x��	���dTX5��I$_O?��d���;�6�w(�b1+t�Z�	���W#"�����cEg7��*�,�������N��+Q�x�	��)��P���M�y�C��5�l�n�^M�6��;۩w�dJWmt���1��{���ќW�ro�~]I_~7I^,�Wp������,�{|c.� ���0κ��Q�#�=W�=)�G����A�C0��fLQ&�ET�XW�lc��s��A�����w)�r4���S+{���&�$�0�`��5�Ч.��NR�`bS�+O"�z�O�5��j���o���3GCp'p��ijS�r���EIǑo�ÒQ����!���H|e�t�B�5d���z ��,���i:�:�O�k]=��k�m��#Q���u	����Cw�{.�{����Fj�=�W�1�P�l���cg=6�0f2�A�=bJ]t9 B��k��@���<�j���5��
j6�1٠jL�W]N��'�?�&�%�����k/�h6C%�ڸ��o.$�g�����I�I�{�A��*1$ Ey���e���4of�k���@���h��K]mHJ�������aM8�5�}���b�� �F�"�#cd~����\���X&չw/s�K��d.��|�y�L��g���t*�C��6���N~��܉���r&���ܼ���^��"ܒ�E��3�Л��ܐU{�L�OHr�(���}��Q��d�g$����P�OfRd����R/o�$)��}%����ķ�����/�%�v_��K��d�ɝYa�s~����<�I�;c@�a�	���`q�#���Al[n��X����Z�0��M��Z.iB�o�O�� 4�)m�ƙ�*���MB.�O����	ʬ��e2�
�ME��J�j�'�����0�W�;�#����xn��AW�'#ڼ��w,&��Z��şߞ��H f�t���G_�(\]I������-w6`���I���k�t�����>�&M��2�k���B7_J��e�A������h{�L�;�3Ęз��/���ӭ����S��)���%�����*Y��xq'�={k��6ޢ����e�T�A���\�k���s���.�0Ǌ��D.�h�}F�����2&࢏(�mm�߃�l�|�".j0J����%��=w�k21�]kEwk @ �-�Ix�L�$ȬS8�n� ���0�H�>[�5gYKC��򵣦�r��b��tO!�Cp[��ld��'��/�j��J�x����̯(�?���Y��Ņ�����L �hAͅQ�D"�kEOS��Z��㍯�lOw��;�@�b��7�f(18(,jx_��R֚#ZoM>�s���0���)?ANJ ��P>�Z�@x�_�n��}Q[Ʈ���f��O�ɬ�06$<:K���kEO˵w�n䶗�]$�m�>ס�����n�Jw$\e���u
fIo�<�}�[�8�ښ�lN����CJL*��*í��D��6<�ѯ:� ������A����zRo�fa�	W��<�}Q.Zʙ��� S�`��ΈX�����s�-7J=΁\����V,%W!x�XDptȰ*z;�C��jB�{̮�݃�b��b�5��N��XlWT#���o��A;Y��^�c�����t�<�ˑ�O�g��a�(� �Y->TF�$���&)���Ӗ�E؜�s,tM���q��y@&�\�Ԍ���N  �W#NY�D?_�J�oϡsc�6�y}�N����g���T͏�>�4"�(z���a�֍\��$�kw��A΢ܦ�
Y�~�����k8�#p�ПP}��kD�U�S�UPFS�&!Z'��T�hC�`m>���!� ���'����𼂠��c`و�h*
��l�S^��mʀEa5>M�e��!�Ïi��?�L(���Q�>����IH�����{�a�tE��ON������<����8�>�ь@x�\2Y��1�&6j8)̦YpB$����U����՗���d�U�<'���P��������L��c�X^�b�B��E=!f�{r�+B�<�P���Zʍ��+8��a�Z>Ab��	�d{н]�bP�I%�����[N���>.�`�E�<���ja����,�۽�'h,���T��6�l�*��]��L�+B��p�D� ��).�3�5h%)Թ�.�B�w���L���C��rg�����%��^S�#���r�-U�S����m&6$:�)�������
6�<����SxG�3����q�F���b�⟜�
�y�$��؈B�@�����z��Ed���R���5���S}�s�6������]H�GE�Q��.O��S��2P��8cw�|���!�
�3��X�ǀr����� f���P�o:?{HCo�ӓ�1����;0�Ó�[m}�D"F�p��dR�Bz����G(�!(��=�W�9A�%Kf����1&'�K���P3Ci���D�/���Rd�L��j�{*��񞀿���^��^a��{@m�^��q�n���+�� � {����N�<p�ƺ�.-���q���KY��W��qtxOw$Y��
������g22Q��I*��v���[s p�(���� EI���yu){��j�=�a\�aN޸)��ٖ����7�f�GeiQ�j2Q�������2��,��Gk�z"�`�˒cp��86lkKs�� ����6�y�	T��2އX.`�k�ŧԟ��y�L�e�1�^����\Z{�F�r��Z�dO��.U/�Q9������"x��$�f�����m��$a�^C3�4wy�@[��{�v�;�◺g[p�p��Z��;������	�����N����{f�z��)��ϛmy/D%�C_�l��4�=ϦG.�5�7�5gѯm���R���@�e���-S��)G����ٜ�jӭ���`2��B�r�:Q�����0h�� ��W����/�����U���h�Wd9|�'�&Q���#t+�E���]n��I{�aڒ������0��4cm�O�LU6}�bQ�B'�(C+��BNէ��i����-�2ы��
�ؾ¤�Lc����Iyt�A��l��3��=�����=]����'�hea}�`�D�Ո���;�{f�O�n�E��w^jk���J���Ʌ7]�����H��͚P��Ţo��_)t����LUս($菱y��I��E7��!�F��7.��ɂ�K�/("6cΜ�-&�?ԍ��zg���ҹ�(l.�����9��""$@��>$!�QÌ��b��"	S���}��k"�1h��iC\1v��X; ,���`��%�8;!�5}�Șk*J\� �d:�y�������1�� ̷��)Y�}��xz�F�T�)��Ě�R>��`�=w�j�%�Bл+X!�xAl��J9����\4��7K���5Yټ�C�J�γsv6n;ܚ0oO���N=��. R��(+�gDt�#.9I�� )��nfy�m��8U�ש7�j���Pl�"�p��xe� n K❓CN��!���Y=z��n5o����]�֟�|���������p{�tV9n%a{5#��kP�oD�W��� )��]O��/SeX����0��5l���ˤ�]IDv��l>��r�`as$���j�E�����i�ʥ�9D<��f�������� ��a��MS�X���]��fq�_^(���"�yX����E ���j��(d|-�C�m��F؜�ʚ��\j��� ͳ�BK� �ƹ*��q�RJ��T�-�u�ݺ����4�|ǳq^�=����h�4�P�̔���O�/Ztx$��SܾUkG��(�}F�x7Ӻ#��n��R�=����C�y���9�h��+��@Qݙ'���֜�D2�n�ef^!�]/���&'�G��l���K��2#s_��8&lz2X�>�����|HX�i��I�Q9���FvԬaotM�C5�I��
�W`-ęO�O�B� cQ��.�$���f@����살U0=��W���}��T��a��Ow�ľ]��ؼB�鵀� ?m5]~�p�`�Jm��aC�])�9��(d�^�ݧh-��fh������Ǧ�S8Hu�Ewȇ��w��]��\o����B���}v_9�,O�/��mZP��L=\f�aW����r��%��sh4��ڝ�N�p�>N���fʀ��⺱�n��1��~ר6�l>�;eD�Vk���n9Qo����6�H&M]�Z��|�R�]K�`b�<7�L��&��~y�J/�����f���-au��p�w��b���������)Ɯ��P�#r���	�8�Qs��f�М�b�XB���}s��20�6Gh�9�<�d�bF�g.*��	��`/O�H0�&/J?����c�確����a���}��,Z��m϶ӷ��/b��j�K�݀�K^�uy�W�a@�b-��uk�L�{�u_���W��|te��P����-Y1S=P��Ti%�m��m\|�
��X��'�$f�?ظQ/���s��_"8ߔ���E��b���|��ޤ�Rku�̭����{�6DNzڭ'��Z�%�j4"�"�r�F{�����L�7��`���G0!VW5�L�g�Ӛ�ox�a��R��o��ls�٭w'���0�#��ղ3I�X�z+Ę�m�'RE�Չ�RY�6����39�[f/��(󜻣w��PA;'EP@l�����,�Pg3^�'��*B�V`�9�pb�u�\oXrh�D)J|�w� �:KϔK��!��8𹆲6�6�70l��R�%�������;�� 5y~�Ud DI�&�@AL�"��wZKu",�8�bR���Zz��Ǳ^^y܅��P99��ѹ׽nMY��ff̅D�%���?Iy;�����N��%�}�6�<�������`{� ���֚&u^�9���?����jp	�>�=� 	0��MA{�ɮ�H��\����� �2R�6�YD�v�����+�lM6|�x�p�bY��J�������7s�J7��Z��t���q\�gh�v��6R��às�x<D��3	M�6�����\�-\�(�F`NH:o��_��=W ��G~^�|��1���{�)hi���6u����y�w>������C'���:��e�X?��%�(��}�6y��>��jC7� �Y�.��s���5��d��W-���4z�dX��tB�j��?��F��(�L6V3����;���>H�o���h�pp'����EZ?��D�[i�T�.P��D�7l��cP���,�����m?�ƾB�	o�y����U�.�W9Q�(�W�DU=�z��/,ހ�RM$���khW�
i�������tk�s�(�)�B9]�1Hq��+�����9�x����4�u	c��6�_?�V��>�?E�5>Q.x̨�]6K�����{�~�h��V����t#r�[�껓ʙk�@[s���x�t��98��l�3`Mz�R�� �V��"<>/҃yb�-�V�^U墑�P�"�6�~^@(|�����}��s�me⛖�X���w�༔�k�ʟ��G`|��Y� Q�;�0���z?�$��g�<��n����K��T'���Y иJ�OɹZl���_�v<��T��yL��!~gH�7]b�g�)Z"�Ȱa;ʞ�W���[�?s�W�CֹT���"�i���C��$��;�-$�^��J�=|��v)���}Ӫz8IPv��h�^ΔU���t�Bw��� �\�j�����d��>q�A�lq�:��R�B]��������E��=��@�p�qf�����2%�3��@����'걐г�T�`
<������_s����[t����kԾ����Xl�I��iF�h�0V&HӤW���#�܍�YkW���ٟ�޳�InMq�618��m��(&{]�ތ�Mu+6���/>��?-Q��64 �~4>utE��P��N��Ww8��y��%�g&��M}�aUZ�9�"��-�י��1i����?C���_,�un��_����%���7�:۩�U�[E����l�0�n8U0�?�wT�Nl�&��.D��L������$K���!����9Hd��7a��C]�zru��1�$x6ṵ[��%��cR��2�#mE�s7�xT�)����ZP�t���f&dD:��T�����8#��Հ�&�x����6�k�亰ڭ�D�lZ�&^�L>��/�]4W�� �h|�ݸG
��ҤCV`����+��O�馔�s=8��#bMѿ���fUm�v��t����&�/<��*m���Y��1i��>I�֐�|��/�1#n�w�6>��ܳ��(��w�4y�k�G�-cN0r���$�P�_C�׳y�a��pЕԾ&�I�}GBb"�-R�_�
�B��t�W��*���BO�����q�:اFЏ��8w ']��ڹ�_Ӳ��Z��>�)�_;U�OίM��m��4Jˬ��z�5�|;*-��(�fe�U�}�!8k;��P�{�;����֨�&x9t�*�dқe������d�Q�m.��z���&��7ZL��T��""چc�0P�p;"u��r\�8���+�s��}Sv۟��8=�� 8K��l���Xf���] -����b�oB�j��D�U����:�U�b������SQM��]�ѱ Z`����ބ�oQ��VG��H,P��"mtG`6J�5��"\V�������$��;�N2}��b���K��z��=!�Kmtp�V1���p�a��-�:*y���ާ�s���͍��m뛣X~�I�k��i����iT�	jSvz���z�>Is}� �~,k�^�0��ߌ��r�9���+vw�0x��f���!�!�KE�enױ1�#�d�f`gT���ó>Z*��Qa�YcEH�����b�����h��K�X��	j�lI�WC�<3�=��h�S�_T6�E�UA`�8bz�����X`�x�{s���=�&�8�;��>`n�Q]�����r���)��Ǩ��s�� �Օ6���W�����Ս��	BQX�tL)[�d�%�O���!#���̑&��/��9C��ۮdy���Uz������q6McS�M��il�5�Z>/?�ꠒH;�J�3^Tc��o\Gw's�@��Qp��e�
����cC����Cp���N �+���m蠛?]	ķ^~lٍ��W�\l;`���3��d�Y_�œty���O���
�wX]�8P�XM5di� �i����*�fc�q>�	&�*8(gb��!�b>,�z�v��[&\|@T߹H�,�vGK
ߴ��f�#2g8�o�P_�\h8 p�R�q��{�Ė���l���Z��(��0R�1����5^:�պ����)�H��	��珙Ҩi�@��'r-?)�sB���w�.7\l�>/���:%'_I�$���؋��HJ�:� (l'�O�Q��Ov��!�������J?y �43V�h�F�O�2�8#�@��.bF�%�x���1��+��05}׹t�W@m�p�ʧBHr��y�*�x�Aβ-��6 '����Ւu�ՃOyT���αﰘ��^O S6_�3�8���E'�ݩ�:ь�	�o�o�Yӭ��X�LƸW����@�5���4}����hp-��EC�_>?솏�g
-��TE=(�&�Y���;u�>��ts��pvD L�i��ۥ���Z�
�dj�����&=+�j��(\p��
���c zVV`AP���p��1 R�m�#v�6�D�&7.Tt76]m�*1c�I'��2QnG�ú��p�}�MP� uWA�c\��֐+�eXE��PN1��"3�Ϻ���Ѫ`�5W�|�p2/�� �_r��m3>��k�u�x�P����G87Qz�0��Yl<\q�OWx�2��b���:��J֬���� ���uM��8�HU�\I��
�7Ț�TJ�%��YV`���|�7�к�5>�S�9ˊ����x�x���w?OW�
7���'�᪚3�!iK����n�'��vOst9�x�Y�(���%|��~)��(Ö[r���Z���[TR�F��*3��ܰ�\H�!���u�p8�R_�����L/�	��@/�����y�s�q��tO�tUQ.P�L����CSf��1�)n��-�zcG�#Z�}�n�u1A��I,�F��:���xѦ��{����ך��i�e�.�$b��Q��=�b��2�ˀ<U/v�M�t;<t��|��`,D��+ie�g�}��������	\��r��9�rF�(H�~U
�A�O}�ڂ��ֱ%x����ԛ.D��;1H��SXc����w7��l؅h'3뀤e8�4;v��܎��ȶyb�A k�(����\���<�Z��c�ǅT�ȌQ[V;���NT
У�"�coˢʫ���Y��*��.� ��$�2/'s���.nŹ���Tkn����ʖb,)r}�����b ��8G*�`�3�x��4��w&yk�XB@}�am�}���?Bw#��p'��!�S�3\�D�0�T�b�"A>�F�[g�P	�~ہ�V���N�m�7NV?|���F ���4n���qD �9�6�������4��y�^�l�qҮ���5#ΰՂv7GN� � �^ܶ#V�������=�����i�2ߕ@R�O�ؖ�諛g���Cv�� ��k�������,�c~�C�?p]*�gG �1Ȩ7R�y��":ш34�;z�0���답7fI�G�s��˧�	���)@�^���S��'��?��
h0�%���@?w��I�^�]�N�S�����\
p��-/*7���K$�[��kK.[��|��\�c2>�U���߭�@W�_��XrlF�#�r{=��?#&>;��K
!a��E��r�p~������|Q�Ll�[����WXj��		����2��90��:G�T檻�5�d�#�)�� $�*����B�D��c��	�A�A�����e�y�D�̨Q��X9f�G��m��3�������W�L[�!��4�b�m�����>�*ѫ�>\�@&x�܌$���NQy|�s?�� ,4V �^W�M1\`l�Դ�w/�m�+oT���3;���|L!�7���}�2{t��=,r�h��@��e�}�ްۃۘ%��K�j�,��pt���Q���[�:��`���>J�:�A�K�c	E�������[%�EM���xDW�h
�;�dV�tM/X��b&W�B��`]%����ѥ"-��y�=b��]��RNh7)݈���h��GgQb����� PbH�t�u�qf�M�{��E˶V۝�Q�*Q��	}���˼�t�sG��Λ_�doO�b2�Z�Kz	1l��i���J���7-�Ӷ�(:J9�S�b�Զ���G�؋Əp:LГ��B�X+,���l���9�^H#[�Q���0���p��owc��4]Ɏ0��X\�Rǎ�U�թ��ׅ6
�HGAU5�Ϩ�ϯ�J;7�4}?�WA{	�"{���c47	���A'o�y<݂������&=��bge)�|��S������(�@�~Z��)���1��
�a�w��x��e��^"��ϵ�qq.ܜ(��7�r<�����*z�G^�P��IM�nB��Ɇz�Ѵf3u�<������x!�#��,����
p��~��5�2���R���p��E�qӳJ\�Z��3>,g��`���L�l�Ġ}�5{у�$���|M�Qg������ƣ�DW���?�e��n3#?�Uo�~��ADE�fJ��OI���_�t���$ex�W]�
��ה	r~���rZ��������=-�5�v�!���`����n��|!�i}İ�7���:Wu�������U�������o����L���s��՘5Ձ��9�||o`��枍2��[ �1��p��k<�?I�z�lY��b3��5E�@�j)�����x@Bb����%���� 10?�}Mw��+%�}��kZ�*���5��~�R\u�~α ��($tZM����%�.�Y띨��J�(�-��Cû����^̳%[�o_��`�2����X�ޯI�&W�����Fm0e��[���F�U �WƧ+�e�h���~�z��cƲS��[�nJ���c�?pf�i���l�X����!T/1�`�j����~:����5#$���z��W���l����FYy֑� �;�v�L9�PEE�����j�@�ՄڢH��,�\޳��R/����A�����M��x~�O�!ގP3�As�,�G����Q�t���ό��%@��&�d���}_���ۣ��l�� ְ�(�sTo��Ɇ4� �]�}Ͷ*?���b��&e�c��5w�}�@w%7�4�����!7��^��ԅ�J��Q�������=!�7��A"�@�Jv�m���:p�v��� ����N���Zg��3nw����H����z9�b��O�)Q����A���r�q#��k�ќĳ�`�&�1����
2A���P^��8,���I3�vyȞ�N�����1k�'u�(`�D��ݼGB��Ч.����>�S�k�CB�/�I	S��z&���)�ii���d<$r��c�(����	ú�I�)�'k�5��2}"O���=HS�v�*�"'ו���~(~�p��J�x�+�wo�jLwE㟼8Q�|�Z���B�}�����TfU/qm5֥�r���b�C� �;�����î0�ӥ*��Xj��@h�p��{��ST�������ik�w��ϭ�wL�0���="�{M�y=����V�3��0N��!��7��������W8��!�z����
��o1ng�� ��h�	վ�	���q��38&��cuZ/�U�y��L<[YQ�Y��yì�9�ť#�u��M~��]ǳ��ق���S�-�sk����> ���:q�(��W�?"rjƸK�r����  w'+�6�A|}c��
޷���2�_�l<��[i��DV%��훋���Wd���*-DoH���hfAp6n�2�a	���ϗ��<m��_YT��&f��@o����ף�Nu��~��rF��cԑ���A"���+�[���'}�1��4����"���h�w�^�U���qN:a<�$�S��1J�DE���G�DIRJg#�"�"a���ڭ:;��]�.U��n��!��V��*yk��|����u�8X�=�	
E�����cT9[c��Z�����*��d� �3�N	h<7��L��վ�x���v�w��c��Ϳn,������b�}�j��qm�P�b�}�3�����<����B\�8��,�bk\�1k�u<[�4��,���� ?��0���\#GϫB0�7�V�z{|�r~��[�h�D �������JW%�)5X�f�)�h2�A�2Z����0�L�x� ��˥89�$�m�~��`y��d}�̑�qY�߳xu���8ۃ���ST�OHT�暸�2Y5��ʩ�+L���ůK\�,;��c
V �n���0�zo3���G��}v3KPbqԸg$� �3�>}ô!`dm�	��$vIW�`��s�sYh>|��d��}��t%/��ՂϘG*��	l�5#_�Dw;\�шt �>�ڠ?/ȫVg��Z��i��v�X�zj�����Z���y�g�S[�x��`�F��s�]XH��?���E�4���
E�*`.y���LD�������Ǎ����q鵔��\6�o�c��~0�7f�~9;��Hq��Z,����0�%}�?{vv8���BNyJ�v�h�ុU�$h���Gr�8��ʆ^���OSr����Z���ȇ�ry��`}�r����E�&a'������tLv��"-��>�D��r����S�	�s��IRe��#�B��i�e}���*?�ُ�ڊ���S3��Q�b��Rx�������E�#��Br�E�m��ڲ��[,x>��qe�a&�{��e��T�6k�Ѕ�^I9��pl𻅞�?�#��)�M_,3X��cX���~Y��},r���>�q�y�����4鶞ۨ���TN��y|*�� o������E�P�SRf�jb{!F����F���Z�S�N�4���p ٩��u^�<�w�*���[�ng�Q�{��I�<�ʘEG�cVR|bh��	�3>}-ڣ"����J�*�*�Jv>��=�k��e.�֐�#�pN�wٙ��8p��f.�i֕��A��B^�ݚx�����C)���B�������"���o&,�Jՙ�X�㊃J'G�no�Q�l���Q_�)|{���9�!�ϬmT���.�Y w5�I+f2�!�`�'�L@�w�ik�K�ܔ�	\k��tu�L
�w�Z%��s�u�N���_PC��y��9����I.(fi���-�Ĭ�4Z���?w�m������l�QI�ْ֬�*
y+l�X��WS���|h���n(��j�%L���L]��1����t��6	�e�w��(�Av�����f�}sa��[�;R?�R��T�e��]�4�)0,,Ci�8��c���FRBԽ�(v��
�{�=�-uu|���m7�N\�y��4��w�=���Z�E �7F�7���~5�͖!ḶKP�8?߲677�������}ŻRi����(@Ee��h8~�^�Ht�?�˞(!~+�
&�f? '������q�я�>�[lR��X$��,gt����� 0��Wt/�����ꯏ�;E:���i� ��\���+��K���#�oAfD5j",���*P����� c�C�4�,�{�%P�X���7�,�*+ce��ZW�o�4}�v��ㅨ�'�0�׾6]�m-n@�3��
�X*�ricJ�D���X+!+-蛥�q�l�q�� '�RT��n�tT�Gh$�՝��<�t��n%�I*�V�Y�X�����m�#`6e���{L���l�FBw�P-������W�C-�FԲS=�9̀�����[:��h�M4@��~���±�^y�ŜC��Q�"�?l�{�V�k��>�	'v�?���'��E�ߩJ�>�0?�*��sH��i��q��B�P�Q��o�Q>D�3mP䀙�"�zW?on�9gl��g���aa����.a����v�\��柑��o���^���I�:��-�
�J�F}��=(��H��b�#u?���*�&��5�o������BYl
rV��$�ne��i�r�d�����F�%5vL����!�<~Pt1ls����_.�ҟ�J�e�W��M)�F*�^3��F9�����Y� m}���~]9�}��)\]^�[�@,�g_�j�D�����K�n�ؿ,�lA��e�p��
J���L7��0J����f�7|���t�k����[5��Gb`��Zo��
 $4Y 6��#�d����#;p3}0!=�˳B/������,9�E�Z8� $1Ų�0�w�_��T��l�K^(����<�8��j(C���룍�n���0�i�sqN��>�l2^�a��^El> �.��|Z�#�_<�@~�.�nЫF�of�o-� 7e�q�|�k�s�ob*�䂍�4hF���܀�u>�]8�W����g�׺�F܉����U��]T�k���j�aM���f�Zb#h$<Qp����7
+Z�����WM!*84�(����
����`��]���տp�3s8��E��y���7��]H��)��1��}��*��G�~� �����~��r�U%Fu��)V��贞2�`���UV�@���a�y�X�}�	����^ag[˱p��ա���Ѱe/���F����_�<!�&�g&��pEG~������*�zM}I��\D�,㷔�%��+���VG"'&�S>�)+E�4��>��PP�W,�f� N�C�F����x7��#�f�rqx��A 'fp6�C|pN螀77D�T�ԣ��ܯ�hd��4-�B�٨Q�Ix�W���]�J���1:�e�X�U��}5`�h=���=J8�\-���9�,���Iģ�U�u���T4����ӟ��OZa�_g/��4!�#���A�iի4w�s٨��ڜ���f]v&�k2Q8�B�$G���+,#8�C,�Jr�㋠��>qfOR�f}�d��9$��v��H.?X��|O�J�y�=�o6K����������Y��h�ƽ���J!�2>=o�ɴT��<+�Ea�J���C%�mפ���AhB�F炅�l��XZ����wkuAi��P��W֓����F���{��Y�r#�tj|h�L�o��,�
tUAw��Q��mT��H6�)kb<�B��j]�����.�uyU*d��0��"��݈�
�yp�l�$|'G�٬I������@`��Hǈ���rSJK`���}E�߀-���D��V�$R�L�Cf�3�C����?�{B*��P/�N��EC�%E�U���i�W�p���<��H0q�3PP���>O�\w�#��/��Q7|;�u��������`��0 �vl�;\k��� ���1�Ro�����8�Q�8i/Q���G�(�;I�a�����
��@�+M�h�0 ���
K�T�czd�IDjO�X6T	���[%�xqk0��E�k�� �F��6�i��D^�/a8�C�f�l�e�t�#{��;���yF�F7�<�T�[y������~���Ph�S���3��T�hR�=Ѭ^��������r�D��� ��P���?*�z�=3��|}�g��HDT�<ʸZ��,����O�܄�Z�
��R�[���_�����ax='��:!
��݁��rkh�HHß���ڤU��z�`���H��|�('��jE
�aN|��@� W
��vM��V�`�0�7�-�l5�cܰ.��|�w`{Wa]�J����� z���xzP#eq���o��<�Z��sG��5�ѻ�1.x�hk�Ƣ���%�-#�B�T)�kE���D��k
�9W�.�<�ښ�������ujן��Ř��8P"�qZP�� z��s�������9�(�@�~�=�{��sV̝����n�SM�(��	��r�"A�,�e ���
kc��E ���&�D�N���;�OJ�ـ��|n����`�;n8`��/��T�@����i�.j:�j���ĭ���h��^�,Ts+�DRrlg��.i�u�Af'H����I	�����ʬ���K�/8�VF�l��Y,��f,9����*o�-Z��%����*;�P���
�`|�M}C=��f%�����td`3+z�9@�vQ�����,�0Bj]ŏ�_D�Gg�����������̋m�s�2�|��s��K9�@���saw�$����J4�>�m����Mp�ff���c|MG��3�GS[2$YR�^��̂{d��K���n�Jj���7I�-�zD��	E�F~z|�F��J�a/
���������qh1��ӄzN���;^�����F�.ލ8h�nu+�(U�	�Yj����F�5���?��(��a��vX�U��*3��	:��D5����ݐ�B<�`��:=�9k��Ȩf13�<�Me�J�lax�넨-�
A	����CD��0��ۘ���XI�&+�k��/9��MF�5x�3�0Կ���T���$�Ӵ��p|�����s��Q��ܶe�3��	�/}+��4����u(����!��]��n��� V�B)M��k�2����ْ?ǟ�������F��/���4��4T8�{��RuQ�0T�����x2�9| ��D?���V�c) s.��υ~�N�ٗ�f1.}���ɢ�"<��B�G[�1������ܰ�Mn�K�=�.IW���I�������h(�S�n%��ױ~�O7=c��`�ڋF
�ѷ��n��}���J�%� ��Fpy� ��wN�Ǆ��f`��"�E�9T1 \-�&'�G_o�x�g)btS��o8�as9"Dbl&�rߠ��7�� �8o�A�g�ϛ��y����,C���r�lW�M���sL:i�	���4Q����KX"G���T/}�"�0�ث(���ڎ�ڽXgDQ|�Z��N�s��xj�:uf����3w+��[�Z�g�����s0��7*Б���y L�s%)߀�`�>�)�,p�:t'��O3� ;��������&щԉ��F�]��1�K�����(��i����U*��+�����>g(u�rqq��;2��Tt_�%�hG�� ���=�`$���ׯ���ݔ������rZ̠~��j�vH�fЦ������{/�L�{��������4@��q��tF�xW������Dy�q�4��m��w����Y�^�@rd:�yT��j>���B��f��x5�>g�5e�g�>��***�Є��}�|�F����ۆ��^0��$h�FiG��À�z�A��� :,7�	N��=��BJ��"��.�!�����D��}�l�#���\3)��ٛ�꼅�I��s���0^����QP�#�$��S>�J��v?4��{���
��jO�;�i@o�����\��A�|뵻>
�@��dK
�p��b�§m�����A�c!�Yl{7����7*P ��W�:[/��g�5R�0A�8�j6�]㳒����H��g�sc�j�]3B����(�Lc^-=��� %#x�mȷ/��T������e��Y/{����u�*�\�Y����9]E��kBuw�6X�/��J6���l^} ���W�U���_'��[ש}��[Q2e*H��t\�0p�%f�w��F���fO�[��1�[������H��ڦ�e��2T<(�2wc����%�^x�D����cA���Uk�^
R���Dn�L��hp� h4,q���5���Մ6��:=�cm�/{��Y��룀�f�<I���6�AznH+�U�)�-M��5d��ju�B�Ɂ�mh(����'NͿ6����Эf�����._"�Ө�f�2pr�E�j�_9F�������ɀ*o����u����O�"C1�xq"ٶ���Ӆ������6���>�1�T�:!�_��KQ}�i.Y��L�2'`k%.�D���2������Q�Lsm�f��u�T�lYZwh��k�-E����:T�3krn�.�#ʺҗ����Y8{[.���L�\�Bߔx�s�5(�$���m���3�J�*�Ʊ7�1�[tk%��B;��l4"��Ս���"Ȏ�N����_$��ynH��0;pD�ëM��X;�4��C�^6���&��|%�dxӘ�F�\|�0�[nD_j�A�T�@��߫
$�Z�s[a>]B>���<҃b�>5���t��<)���@~�� IT����ZH����Ƽ�����$���n���)��p� =]>��T���@�^���GER�Ig�֧�7K:�,P�W����p�g$ult(�y �x'�J7�Y��L�R��Ds��Iw��L�����(a_�ą9�ː "�[Ӯ���%�elT02=����9q,m��+�5x�6?� ��]���Ċ�E�ڿ�s0c�+�Q+�3)aV�˖�A���f*��At.��~F�j'M���6�@cWڡ�h��f�8HG�n�d�u���J�y_���`��E��
t�������&ȩe"�	�޾�v�%�=U�A�}���_y���$�k�UX>'�������ճ|ܗx���F�=kWo�ӹTDU�<_ȼ�#�t>ԂU
����� ]yHnT�E,�@�5�4�35s�#W׵