��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���:����~׳�jB%�y���	��/o�5�n'э�5�a��U��<;�A���M�{ǾZ�Cy�f��ѩ�����@@�����2V�o�ڳɣ����@��? �bP�:d��6�t4�,j�1�^
�{-/ԷR�V;��X��Y4ׂ���.v�2:A��W��3�y ���'��hf���&U =6}�Ӽ��ԏ�xa��lɚU���[�H(�dܳ���R�~S�=�����N��w	Ș2��Ô4R��kі+E~�8Ƕ�R�W�h�4-M|��ʄ�4.�}��x�E>�ϫ�.�H�����Ȗz8���H��|ȏ���5�>קs
a����k������t��L�g9ɋ�X���kwc��/�6dI�5�D��(Yt�Y��?��={Y<M�v�4�`{1-�E�n�>�VfS�u-�(x���Z��O�\���{w/R��u�S��D^\�Z�6t�7�sWU�BO!��ݢ�WR{�uQ��y����p�=$+
T��r��Ne����϶GX����4�8X~��L�~$JsZ��,��˄#���s�	�#��$Ԗ}06@;���|g�c']���3��憭� ���ًrx���=���Q�3׃�$�+=�x�(]\��B��C��D��a��%�Œ��9~Ju�����;��a_P�*��*���	Z�r��|y�K%���8Լ�*�BvN����Z�4��=g\�T�+���<��paWa���nB��?<��=���tP�N�"�5 "���)-��*��XL�a�O]=�xw�R~��ҬB�{ܼS�)�F�~m�8�!\�/��pz4��(��˦�~�A+'F�p81����w�/Z1� GjrM^��/���#�P�2d�:�I0eٳQq���ə�ۗ���q��A��$��+�.�>@˔D��� �x�BE�0�ecV8��?�	��S[�Tk��E4���|-Y6��l���ż��̟�G�7�+�ep�C�_K���m0&�4�rHA ����� ���vQ�T�+�/��(Ґ��F\� }�у��>W}֭��3�:rL��g�-8�V����]U��T�9}~���a�;�/�C�ǗZ$�9�M���$[���p���%�s��ј�\j���78���mJ���� �K��vx��S�ڻfw]U�ڢwaI>9[��r6=K�&��Z}I҈��^�`�98>9�N'�B~�D�`5�B,�ψ@{%�u��j�TDUU=u}�5T�#���B����[m��yo��-g��r�#�ko��r�5~7�,bT赐˞�7gS��ܗ5˥�Nq����!��r��fb39�� �[?gQ��R�w��*�X'5�f�n\�� !����h���y�&�B#�_/T���+B��q�L��Q���X��"���y~�Jˇ��D#�Ӧ�#��Snݝ)T��i�u�|:����%�J�J�i{A0���h�1%�M�t���.���W�KW4R]�ɐvwv����Wɥ����{�����aR����M����H��u3P�*�3⥏
���:ݰ�f��[G�и�m��\y�!�u��F��[�g��'�R��Wnn����l��˾x��݀�r0u�]��X-p��n��U�?�?��j�*�`a����:��y��!o �ى���m/����3
g� �zPc}�l)�9�i�s�$=� ���#��9�g@�-k���i�6}���OvW[ƾ����G�w'��\��x��蔚a�6���	�F�#Gc�2t|o�)���m�E���l��<��)5��\���YLIz���{DЗ�B�1T0y�g��z@Ks}u>�na��Q�;��m�r�lKL���~���fTCz�a/Xm�^|�y�S��]ۭ�]�Ll�i_�����>>��:���#߉`��^�`m��ȨN�%�_~u�}z&��2-Cu2��5]wұxCE�U|���$�2&P;���
P��d�Uv��<e<�BHz��'4/m���ޚf�&ġ�ɽ����_�9��1���^u�;#���
�M*xi�J]�>�7�h`#	�\�ӨO_� �q|�����O�i�0m�q��᷁���)�DG�)!�x�a&�fPh�ӌLs��ҢҴ	�<:U��TnM�H%q�c
I�h3Y�( @�gg��h���<��uۏw�adI�ٌὢx(�'�H9�ʚK+��(
ä\OƝ�����y��T����bM�������u�J��M�fo��5����#��/"�-���$f���2�z�e.�(N��&����W{�\7�|5��&J[oW��Š�[���40j�ϖ�T6��%=9Y�2��x�W��S;o_q�[|�FΚ��`w���eJ9��?����35�h�?�r����E��%�u����I���H���5#ƈ����o����<� ��9��z� ���������,'j=L�4�����E��&�	�>�Ot��g��{UEl��^_M�G��9��۹-�Q!Inq�,=s��cE������47{�'7�t���p��2C�
��X����d��h
�/`|	��jJ9�6!u3���f����E�: t�,GR,�V��o�S��`k{
'�Ko�A/][4*Bp&�z{����a��K�;ѥ�L$�� �SjP�< ~�9cr{�$<Ⱦ�ӈ_�f�+5�q����5�� ��J5R�ZV�G�Eo��E�cgћ.�!F����F�6�G]R��~?iw$G�_�Ƭ��}r�͵�S����<ҙcZ_�1��c����LʃM�-tܶ��ڦ��f!=@"g�A`���{p)ԝ��M*���m�Q��ѥvŪ��4_kɴ!e��1Ȑ��*�B�	�]#�Z+��(�������=h�2���ǣ-E�oa(��/X�14�ʇ[�.�NC��`rL� `���KN��7ZCU��|�M�C	/���M�3@�9�Î�rA��q>�����Nʿ��;#/"�B �g�cy*���@t|�5��$n�5v�(Vd��ͯg�bEi���afG��M>�J�-�����x��p���_&�*�/c�?⤼pF+�s�쀺�p���E�}:�� ����<��>nϧ/X����b��y�d�HG^Q 1m'��娵�I�`�&���z�1�b�6*X{�5�[j�k'o��V.�L����;�-��[4�[H��r;�����Z��|Z�ߤ��\Ws�+@�@��H�S����Z�����!�'��M`�2Ƹ�q�2�G��D�m�v�]gZ�̣�:�
aa~�ȡ�F�`����6v���#�$+��!xȷ?��w%u%����P���T��B�}fe}vg�(��Я��j�Wh�3�J�=��G.e�Ɉ��y�x9uB�����Ѱ�B~1�����#�Ns� �s~�����Δt��ȿ����P�:rE02����$>b��$�,]�*d�/���/=�N��	�{�ŀ(��H����f����8)�����)���굵F��Y��ۘ���Pa��x�{s�d!�3_��@��� `��^���$��B�}���fwe�����z���^�������9�l~�=�)�|���4lÚ��D]�qT<~2�7U%S�Bq�m�M�{��Ϭ�����T��j��i#\�ݙq���A�l,r.�������6Y�C3��Ut"QNT��(�1x��3��2�O����¦a�ҾW$�y�͌�S��4��U�h
h�)����ZG���^��u�0���S����N�a�Gj|��'��%�ʀ�5�Aiq��ʠu�B��E��S$�E��P#���Eh�5�v��
�>�e���2�[�2bxp�o�6���Ԝ��c�P=�����q&��&�aW1Mk����;��~�o�*�z}��b�D6\�!'[@�{qCq��a!�^�7;�cZjf�O���mQ��@{R/�t��Y�a� ��v�SvQ�N��Q��
��&�.׭�n����Ӯ�C�܊�_���0)L���Vϑh��T��i��C3R�i��;;��t�f�A���_6��e#���J�~�dFK��"KHJѶ9�sǡ�$�^P��|u�`�u���w �f!���?�A��;�k[�)}2Q���d)K՚J�O�=�Z���y3�8W�<Z����}1Ke��X����k��R�B�FM�l_�.����>�$`H:v7��1l�h�b��"u�6�t��
��}IO���Q�+�T�(Y���.���a�V�}Q�Ί���$P��"�e[@_�<��㯹���Ѿ��f���NkՂAE'���"�_G,M(��Eq��Ot")>v���i�r�2��/nhí�����{$�&�vyP�lU�P�i��1<E�b*�+
R9�:`J���� ���m�����.7�
GGj�g8�C�C�d=y��e��2�,g(��V��
�M����
�3�OQ�A�����<9�=� �Ȧ��{���Oޕޗ;��k�+"����d��cHx	� �
y�>p�KAi���V�Aʐ!J
���|e�s�z]P&��s3ZA{�ߺ�ag��a{�
�x��1���R��$����[�<�Y?{���>.ŝ\n+{h���}�C�����|��g(n�f^� k_P5�����R+J�(���z�q\��q�W��G���!b�p�̬
�0U��Y0��Ql#Wn����r�ڸ
Ղt�L�ȉdgC6K� @�zVGS�h	��ӝ�|��K���%i:Wk]��Q>@y�,',����z�O4�Kې���.���_��-K�N����
TJ����>h?,�
��oJ��vey�J��8L鹒E���Vf������m[Q$6֏�0��ƏVz`fh�O%��[�)�7�vM�ըT��W�( �aJ�f���+nx������yV��}��"d�R!�݂�>�C����=	�;4{�ҕ���H\��)�C�᝝������<ú�^����{�R.�+�l��J�#"4Ҍ/��׀���v��cJ�͋����%�!�@^pïL:h���~��/TU!����@v�0�
O�_^Ζ�>��E�|�V���b5i�fy[��3�Ȯc��w+�����j�5�(�,�5�f9��.eE�h���}����g�l�����'o �h�Ō���x�(�m�SW��` /z�[Q7_��g�k�9��>�yiT����ʱ/C�
����D(�>%j�I�Jʸ2OQ���m���eo�u���73����y�Y����\�<BnL�R��P�;���ݕK+���\P[��W��dؙ�%�cwD��xO�܅��	�kv�A/��-j��<�L��7�����k�/��������{�AP��gS��X]%(�x�G]��ﳆ���^{wk2�8fcrV����!-'�0�X��*�]�y&(�H����#�_��f)^��᯽��ǝ�j�l���2����:�x��N��7X��Z���M�~�j�G�^"��ɷ�T3s��~K3�h~ƶ��7�6o]o����ę���ų���pkEYϷ�$ܐ�RI��n&���=JW>z�E�)J{\���a%���m��#�T|��)l��#
����-,��*Z2�;![��t��A��9����a��p7إ�ޒW�u;�-�0�o�NE��=�(�ʊ;5��� ��^7��au,k�~���?�����5k4�s�pܶ�J(�� �>���:�f�{��WIL�3ryYw��}�-��³�b�tyRD>,��M�I>��!I�t��RYQ*�␣Jo���a>�'�{��/5oT<�[�=r�}�q~�j��-�To�۠e-��ΗF,!���ܩ� �mp}���|#�^}�������!%�����zk}ه�@f�=ESI��N�������R?[�5P��ؕ �傔7��^��L��G�O�I�k�Éq(�G#o���o���V�"F{�3�/sb��څ���f0<������+���$0<��u�kpʎ�J�&�$ց�|ԸIe�c�ۥ�Ym�T	�!���I��C&�:�c1J��>�]��Cэ���I\�j�]��V�l
�s���a����N���2\��7㊪x	�x?c�����y8�uQ"�n�.}��)��m@e�{ ���e=���v.�;a	2�kK�	xӐ�-y��SI��Y'{�F�{�I���?�	���-�)(̱��}g��f��<�Q��V��#��'��D���~�]<-�L�2��hXΉV�@-��"v.@u���'�
�����T�p��"�'��!�i`�o��ݐ�D��G��j�d_Bf�Z\|������x���*��$,�zz��{n �x�7�K��Ӿht���T.+5�<X�� ��?����#��a-0��_�	�?�]�ٻ 溩��!dK���>��6QO�ZL��JH���T�M����c^m�Y:�x9�����L�A� z�V��i0�t���KN�?"WlS~?r�bƦ���m~|c�݁�5�!j��J�p�8h�U.�#��C�mb)M�������#��/ �T�����aK������4 ��J{/0pŔ?Wq.9Y��o6�;+H�>�1��;��}�9n?�f��\����{��]��rA��yV7Gב��:�7K?��4�a��B�2����pӕ�4�e޾�T��QsX E"s�`�b�:T�f����w,�.�g2����uL�F�'sY�����=���=��]��Z�8r��c�TY��{�q�V',Cf@ �d+���r)f�k��H�/�U�r���l*�ک��T��ڴ*�|��gc��$f�� ?_S2�'v�x��7F����0����yf+���_�Y�3���΀�'}�nWP!�.��-�_��QZ�8���kC��	 �����k�W�u���*�LP�"�'�m����A��*�&%�e^g®�D \>V�#[q�d����f��v�vĨ<3`eo�3�9�P,����I�_4_N\��5I��#2�f���p�Oeu��s۞���*Xc$2�w-SI�J�|���!N�!b��F�P�z�%�~$d��Rΐ�œ�?�@�_qe؋'�&��� �1[���z��j��v." �������˲h4��Yh7T�5+lQ�S���:�z��滆d�L���
�J&����zƃ*͡X�%O�ɡ���~������2w���e.��TЏ�+X[�g7���%ϲ��e����n.6�����3uDLc�_�M���.'��ڝ6�)]R��˼i�j�d;�ԯ�\�XO��r4��� �r�GA���WA����U�M�O@��ʦ�D�K��b���������h&�Niv5�Zy��(����9	�/�y|��oD��@��v��U���N��S�"�S���t�Kg�̸*Ii����5��Q�l������ͯ4�-�V�6���͚�K�Y���x���SP�]k���c������Ȗ��T"(� ���4g�^��U�~�_�+��] OJU�q�GQ�-1���gۺ$���׺|��
$ǁ]rvJ���*�֧�lKX����g�[W�T�ڲf>��i5������F�s���t��M�Ҿ�j��f�k����Բ ѿ=(D����[���Q��ַ=�d��祦��5�����l�����㳏��}a�~%DCN��D����{�=:�/���-N>���6���i�]AQ����x'�6��x������i͞EӉ��=�h��a�	���cˤ�?"���Gp,u�����Ԑ�� /K������TJdy~�;�!�N�\*Ǟ�\��f�|�.~�K8+] _<%�&�$߉%�o"&�O�UƎ�Ҩ��-�6̲_u�����o�!CJ	���n�HgC(%}|=9�fT�ꁯ�E�8ֲ���1�d!)?��HS�D`ۅ.���*�­ j�}��#hi��,�3U}�5@�#�<��p�h+�.{h�*#r�v1}� �ܶ���^'���H��豪,�~�xw����G~�R$q&����{×��F����w�x�U�O�f{LmȤJ����H����$�Z� �KaG��|*i�`dk��My��h9��4�6�p��'��,ii��w}�O�w��);;���F��el�[2fXP��0�ݧ<��)%ڄ$<��O2�ܵ��
�
��ՄX���.�@��_JwU�(�m$HG�au��&��n>
h��[���U�	�3ȷ=Wg���D.���+7�Doˋg$�Q������9�@6m��
����L{�ЪnY�o�j(Q���݋4�]oR%Z�֜Z��C|S�o��W"Hl1���~��@�LGiH=t��XY���IQ��kd=]WtX�H�����{ٛ��2A;Q.�3�e���Kz-��p�n�w%�$R��w3�ۉ�s��.������hۤ��H��ͥ���_����8%C4j��к�(+���tO�VmnEX�H7&��:]B>hX+p��b-�v_B�t��� #SGB�ֲ.���=��]p*�JfCͦӮ6�c)h_���t�l4�<9]*����SJo��-�A�� ��Q*�:mQ�w���BM�����m/xw��xQ���݄�:��T�j� 7�Ȉ%��BuE��V���ct��p0���7Q� ��]<��/�j� �TÔB����bn�AU5ڰ��a�w�xJ�:���-������&��G�/I�<���ȹSzA��r1?���`Q��0<���j4�W�\�BƻT�Oa�Y�b�껁Y�zOϬ��2۹�n�Ug�N���0 Io!�<�� �V�c���&�t)2�r����h}ɣ���?��+��=��w'�=.i�B$9�q&��c�糄��hKdb�Q���������-��6yX�	���>���~<d��94ǒzĤ�d�=�M�s�)��n�Z�� ԃ֬�$�4p�x ���B)9e��,z��`��I����W �*|=�x�IP�3ޫ�T8Z���j�Ì+��Ƿ��bN[E�c��w�@Q֛骣��'߽ʹq(���W3��}�GGAQ��ZX�� #"��_���٭ZM��(��m���`�96�+*�r�
�8X��a�*��gK��*���=Q����VY��*ӈ�i�MR����877��c��)*S/�]�-3�m Ϛ�x��^oy������NE��f^~�_ ݻ��4�2S"a�Ek5�@k�Q���V�ǦJ�G�����<��7߬]�=ᱧ���|b�A��:H�eaEi�x^.aġufq�Ԙ���V�j�c;������ �W�VGR8(�AH� 9���!����xF����:�����Y�:�	V$��K��٧�2����ĽQ��� Je�,�q���'�>?|n��y���6��	�r�?�/[�!�Z�s9R�c��m>i@�g\�Y��G,��'���ʎ'�3WC�(�^�cc�@���o�fkM��=�K�q��<)���~�B�ͮ�5���Ļ�Qx�,��GRZMq��ye�V胶�?�&n�q֙O�Z�)*���g�P�P�y�s�j�԰y/ߜF��$<K/1�E��e!8�ĉ?F4gA���r���.���5;􁣗����C6)Q�j�6� �{�a[΄�b��Y���qg�$s��fI��O�Z�~F���c�>
�m�FA+#�x'F��RP����.ʎ|]]MkP��2��� ���Hq��&�ZL�2'�$+G���/���\�	?sj	�9�l�����W�i�Ղ��dA���)K�nr���"��#`�`���N�H,5c��%���ElE�$�!�a�Ⅼ=`�%L.=UX��v��n#P�`��D*;�$�//�3Wo���;�ǏHEܯ�os�̨d�0�ъ�#Co��3��!Z1P�}FBN���G�Jr^S8��u��|�T�X8�R�}�x�U�QW눠�^vt�p�B����Y3��I$$��2�4T�Rb*B?��!�'���j�d#?�f�����|J�jWA�+����p��K�KFӽ񭕧�@;4/�q�a���s�J��z�ם��ܓ38m��i1�m�� D�4���P7�6�/���O�r!��JٗR4�Ҡ�;�v$�J�Z��=�Kٿ�[�8[���W�����xAykj�n���ew�ze�m����!��/�~�J�Jpl��F�YB��n�R����<�p�ǂ}�ƥ�}���S�j-ܿr}�x:�!u�r�[��փk��FL��ͥ�~��"45f>y���zl���h\f��n�=3a&�5p^Q�yRjKwZ����AT�c��!���;S~9'�#�i���~��c�(��@Q}&CA�R�RX��ħNoy�M��G�����u�``�tu�W��ܿTk6hx��#,C�5�f�P����X�ږ�Z��N���W��1�D����O&y�ɶ���km�I`�l^ Q�%|�6��
��C�q�;8�]8]��)il�ԭW)�O4��>�� �|��2��ck��?ME+ Y���e��cYǗ.��1C���3zr�VtGC�,<��0ͥ�G^Ul6���#�Rma֪g���*=�f��v�vAj������a�����ppM������xW}A������u��"P����: 7��zK����
1�H��N��~x C��}�Wg��7ɽ�"��<ؕ�ԸG�ws�ߠ�����{XT�Ȳ�i��??#o���UK�ܵ�� ��|(�6�Q����f�Q���)�������y��x�y�ש������["}�[�q�x(X��tBm�O�oD�Y#L�sLW��4׿��L>���e
d����`dޚ�7���;\[�4* �W�݁f$����䰲�̘��d3�{�؎����&�x��z�vQR6s>e!���l=�PC��?b���H�T�,]P�D��&v�)��*�U���%��R���ND��(���9��/;�I��)�/5`S��U��j�ɿ�o���?�E��5��	�Ǜ����4���1`�=�.���t�wsL�|��s��g4���%��=P���))~��۷����]"�
��(����� U�ry�'�H�� Ŏ(��[�6���w�M��mj�^B�|���G7�N&��K�H��D����EH[;��I�q^���˳��C���������ђə�umΔ�$�j�]�I��N:��^����ކ���
7�sM�	y�ۓ�N�ۿ�B��3��d?�{�ԑ���m�<�>�y�� +mg��HH},�0������i��z��GK0�[�������f3�\& =f<5���S��%D=�\-�j0�(�5I����<g#�5{"�j�/�S�X	Y��Pq"Ѿ^̴+�HTS��gw�d��h�^э������-��ݏH�`���%�UU��@�"��E�&�9K9�G�������8����:���@䬲���P��z%�q�R�R)�.z��)����!鏹o��_�O%7DZ%��~�JP�JW=c�ӑM�f ��)��iзN�=��E��	��}�~�u�����I&��<|�]:���|ˌ���@Os��}t�o�@�Ԟ:]r�q�٬hZP�PN� |�	�\�u=�w��#�(b�F'Gr@��a�E ��8�
g:�7	2r!g)r�����<�����p�2�{[��o��J%���w��VY���[������Mc��:\�2�~7| G�K�0�J��h��zo[e�{j�µ�Џy��BX�݈FX���2�~���ެ�CC��0����F7�wk��iq�J�$˞9Si���[��}�5ſ�gե	�#�%�
x���3I%J6��J9A�Cy�'nUމ�-���v��6��U#�=�޽7�2h���P�9��<��C��E��3���/��lA�N�|��/����n�P��a/�ݾ}�VTF��,�\/��_���ed���h�K�V�9���&���Uw��>��G�;�u���ZrdL����Ⱥ�#6u����Q)��#Ǿ`�{Y�8���-Kz
����'	�H�Â��Eu����郏�@�����i-��R�&�G�h$��<Q��h�g��1�8Fɟ�j*���(1�V�j�%=MA��o\�����Z��bfkOx�	���&�.��_]^B5������E<h��(tG s����`m~. 8{`lk^v����L���%��v�בH�E1���q��5���9���Q:�M/(B�l�NF[�k�'�����:Rٖ�z9쥖%}�cZu�kq�ǳ�w^΢��8�<!>$�J���gy�I��f�� �!�,�ǜP+�Uw�V1B�>֬-#��9@�v�s���'�'�(���XVw\��'H���'u��������Ҽ�UlO���{4�0����f�������ǁ�$V����4h��h��O�<?�9�쥭��U!�shB#��Jե�4J����/�`�&����HT��{�!���j ��w6��NX#� X�:�b (�Z�s�F��!�(z�?g�33V�&��˦'D������G�/+}.�
1d������/&?� �ߙx���:J�w�9٪�,	g��N����OEV#��!p@Q^���f�����J�3�0g�v΄m��rK��i�� ���k������y�����_�ʿ����hLwd%u�e��|��� �L&��Ɗ'mhI����{t'���|W ��3&��nnu� �"���e,ҳb�`�K�c�D�Bs���>�'ng�:����V�h<�Ϭ�Q�ĉ` ���^�fv�wJ)$+x�Eh�^5pX�9�bi����~�l�)�,��'zQL*T-'�Z���Q��u'?�j��(j��UԤ���9)���t�����}D�=I��3�`pj���EA=��q����ZT�$�_=
�P�H=&�҄Wp��z�4BO��L۔x8��[8B���B8!���Sk��}�(� �[��8ΥB{i��P2��:�l]�gxo�x�%bl'^K����\��N8�g��+f/�n�z��w<+�����:�FpN6{�%0�s�H��ܷ
�Ѻ����e3��x���yq�Q"v�dc�/�{���Ѡ�kw\�p�ֻ��l>�1�w�8}(�y%r}}J�O=���.�A?P:n-�I��v�7_zϵ�8*��w�B��7�X����w��{�X��G���o�V�-�\m�����#�iC���etb�L���	L�[A-ʟ���/H����zj��|�D~[�/�#:!�+�Gn�8��_'m;��-����e�����n�2��e"Dlg<k�a-'�-4�$]�寿�C�h2�)�X�Ke}��1[�Äj�	��ehs}n)��
M� CȽQ%�V�k�	�d�.oF��:MH�`�PS�iR ��h)���!!�u������ʻԨ,�-T�k�";wNos�ܞ���ћ��O�������iR+��k�����
�#�,.���jN����E��V�E�����!�:FoI�,!�J�Ĳ����U��*2�zZ%6@`������.����q��*Z����"�
��L|�	 �0�VQ>�)��;j�W��=]u��Ǎ�:7��y#7�u��l����t̔3!���u�3��oS�m��9�&�62=9{�U��l�DK�9 �NF�:�_��&b�m�7[ӂ��������+}��ˁ4 ��8�zm�6��Fψ����\Z�۰mT\��p,�_�U���F��]���x����F�����O��"<�m�{��Yz�/��wݟ����sǣi)ң�\�����hI��W�?�c�$ܹ���
c��i_���+,fb�SŨ���T�&}��Ї��1.h]pR��0o
�ja��~��92���wU��'�)�bP��F���-d{�h$/&�^��*o{g��R+
� \3�	9��~w�K@ ��E�b�~�.�5]�V��k�k)��g�[7�1ti�=R���Z9V�Xl�葎CY�ye� �k�<�c��u���	��8<�BK�z��*�.�	4;W���)�W��\�c� �6:�d�׊"�,�c6�~쇑>	Զ�?'�������(�3����"�/�-nȫ	�Iy_R��T�Hs����P��/s��\��%�~,�:m8v� ���TQ�����̻�ba�R���lr�|1��2N�X��<���Y/�)ހR��`��M#C�����~W7R	盽��d<�)�ς�$��>qPu �r[�μ��N�)Ź���ʭ S��[�[$|Mp���f��T�߅��hNhϯ�k�|�����=|�	��n�@�������;�����|7��E�˝TN�qjm��m�mC��֕��m����-�Z�;4$/Hh��h�w�w�`{�6ซ��i�;)�G����$��o�O!�Oz�e�#�/�  �6Б��(�׿K�L�|�é���Q;ʜ�y�����)ҋO��Q ����U&/�/[����`��s�´	����Ӈ��
Y�(�����e�M�)2X"M���@���%|�(��'��X��H��YJ����2�d0��m�98-���"��զ�9e f�C�<w���xO������3|��=�S�d���Q��:�rj�U.�|�\�)[���U�Au8p�8~З�g�%��f��DܠM �)ޫ*���m�Hx:�srو��k$�)�7�s��J'�&�b�.�Ab��Yp^���R(��U�(�@q�ߒ~���s����L�3��p�`�n8�W�K�z���/ǬlDVX����{��\�R1x�����G�	혅��g$0ҋ�ݖ�ǁ�s��x{�T3��-��g�=(�}��� + >�g>cnN��V�W��i��Ԡ��m�O[��y�2-t>ퟺ�f��NQC�境L��A�h����nW��F\ܳr��1�h�@4N�����]�\\h�v�![L�ͨ�sqNO<���	��n�|1��{��Mx�"G,Ϭy. ��Z�`ʺ��	.؃Fk�+��ˏ
�����;Y�Z��������
v�'��4��?�硫��L���{��u��y���:��Pr�[�ԯ��H����;�j���=Io:�{���:ֶ1./2*����2Í�܁��%��i"���=|ՋݠE�V70@߻L��Ti��*&���c�o
��2�{�^P0���Ԡ�����$�Q��+6B�VF�Ó&�N���F4K��u�1˸J�O�'$��4��"ξl	s�B�H��؈��=`u�E-0]`�ci"��`�������P�2,b�9RIf�䨱�&<�F2�3��3�4���ňŕu�D��0�G&)_�ñ�s=������
o\=��x-P���W}�2�҂|f�rY�yJ|`5dB��h<#�C�Q!���|{�|�/�-xS&Y��O����>1����6�
�R0\�a��r\c�eneљ� ������!EirH=A��@7.�x�g�/�r���� ��_�]�����9�uF��3�Kʱ"UOq����e|G��/'M+~�����3xy!�{����V��h\X��;�:���S��k7����gSLw�^��������]�`�.��+a呋�x������ƛu  q)S	r%��B(#w�GL�;��`���u�.6�f@�Z���)�?��.1i�$D6�ɬ<�;.��gZF�LXΚR��T�@����Wp�H<��?�1���5������	J͊ݟ��	��<�"�9���N	�;��g8�hysMA���f��X���O��%q�:��6��ͩ��O:���5Ĩ2N����!�k�` ��s�CG���8+�~�7S���J��^L 7��5&��x���=0�tz��-�L/:�=���"�����z����l`P�9�'5��?���:�xY�ʆ��w�g�N}ii��Ȏp㹰�.�D~�ݤ0��!��H+�h7w���]���Fq��;�,PX^"���#���C.xy$��hk� 3$�'����:�m�>�}C�︩H��C��8ˌ�p953:����D|���v2B$U�@��/�֖��r�M*��8
�T ��3��u8��b;X��*�a��j�]ihr�Ԕ�fH�Z�C�L��b}���:�ͭ���sF�;v0������ 6dh��ࠜ��c:;�^��#�k�������\�J��M釿���M] �����'(?-�K�H�U9�/���Zq�x��=Z؆馅�GwYK}��tƖˮ�T��7�/rr_.��q�zU�R9�����������,D�G����Wb	��!�G�6-�eRCN��}x y2�Z�P��c]`�ي�b�YCi�'4i8 ����/�և"��L�����i1Em�ȩhSݨ���T�-K)�$B��F��1tP���:Bh�J;a#�!�S�S�$ �l� �2�5O)oC����ݎ+�$�"�J�h|Ѹ�w���g���j�!���¥�F��X��ʾ�c�!p�]�^�n��Ph�HB���P����o�/��������v�gg�-��R�� �މ�&��{b�7���Ŕ��vO0=@SRV�R�+��W�V{�����>9����>����}�b�W;H7���A)������J��D`�\PG9	z����K"=Q7~f�A&@�WF���X����y#6�)���~�[��@��y�����u��j���Ee0E�+u���7��^�W��&c�G
%=QΝ\��r#Y���|�%.�VK���t��1"�3�[X��5圶�mu.K{<}p�8j�Fa���N��Tp�J��ce�<���i�Ɠ_@�}?��H���K��������ԓ������1������g9��{>f�x�F�թb��m��r����
��=�o41�n�: t� 5 �������x��Գ��L1��4���hW�$��ɵ�B�Ioί]���M]���� Sģ.��5l�L>3�c(���񹾎�;(@�̜�o>���>��&&� ~4l*C
Ȩ*Y���ғ�

v>+���Y�l�,֜%w]�G���൳�1��;~���/K{u\����F�pǂI�6�{<n7U�Q�j<Ę\�vXe���9��?B��r�[��,�`�	AL���1��owӱ�=�y���ȶǹ������$)Ҍ��#���K.B�B�w�#-���͙�G�t��H�(��1�~��
���}y1�^^����I��4_�s��j<v�5
�X>~M1�%x�\��l����q3$n
�{�K�ŷE9���誀F���w�hT�6R�$ş�������yS�X����C�,�Z/ ,����n���ÑD��K���þ�0�3�I�d��UN�����^S�iK0ѓ6P#�p�Z�^�&��3;z|ŏ�,��� >��hM2��IU��YF��})���3'�
&9�pY������n~�5�hD�"���h?���8n��x�q`��S۝d�Sw��t��U���R����@$1��b��\�?�5����k+��H��1�ZX0�:!kk�?̱��|�˷����9����A�p./��nv*F��*�ȕ�V��,��`8٤�1�]d-��@�̄�]ϱ�������f�f�v7�f)&�R��d<�56�#��
��\ώ�Ξ���e�Da�O����~��BKc�!�tT��a�)E���x:���	3�ǥf6���W��-�~�k�?^Z����� ;�E�i����O�Sv��9Q
��P�'��0��<�_�%��7�aw-����at�m�!�D�/ HI�01#�1\h�4]+�g��h�~�rt��Jd���o��vn��G��b�ߩ�E6�'���N(rH��3�o��}���)�_�UK`�3T�P&�0v:�I���iV�����u*,�i�D�'E"�]@)k��!&�c�Vz�u���WB9mZ?r5��׃ݼ߮�=}�?�֑߉��휗L�2�{���82p�K���Td9��qIQ<^�;�N�X)�_��AScę��ۡ��mӜ˩�Vq{�6��*�q����L�.J�W-k3#�fg$�U.絛��-
p:�C�Ь�����N@�Z(��j^s�'�A�	z���{�Mk��e�ۢӂ6�sW�/;��:�h�k���R7�2a��B��6��Rh����/��rx�޹nbo�1TŇ���{��lo�-=i���*�â(U���V�>A�ǁ����	����A��c�{�b� ��DXe�X�L��md�Ȍ\)_�i?١j)�����3���}�Z��hE�"��5��E)�^����t�*�<�DO/�Ъ���Gыf�9��S�f	R�#(M;���z�2*��O@|��S���K�o�����qAu�<�J��u���S	�t|�15e'1��ԕAJ�ʁ�@�:D8�{���rס��UYSX�����W��Ƿ@����}0U;�YO��6��,j�� %��ݗs`���,�Z�9�3���s���I@B�s������^�o��THk�<�I�q�,ۨ��̈́����A�j�6[�����"sٺ%�Dc�B�q�8S�g�%g��J�Dj�@ù�Q6t�|IX'OC�)�� �$r��U4�ެ�X�%'��
�kb�a_�Z�m��T:Ә��@���$�3=�5����˔�n���0��}xޘ��N� ��E5Ą��a�;�Y^2ʐ��,R
aאw�q��0H7�1
nK��%���	?�S\$�ÏKKF�O�#vM<#�`��};.>�s�-��{�7��9{�Ӊ��)���kD�'���=�Ў��b.#S��Į��|��`Ǡ�U������V�XqcO,$>^è��k�n'R� L����b���~�țd&���S��ؖ��op,ұ�Xs,I��$�ň7�qt�
�J�k7nh��<�f�Р4�Nv:�yI�$��[j7�X��7���q�˟�Y�����o�ϣ��$zG��anl�&1j��,ދ="����M%4��o�?�zyy�wɇ��c����J���Z�NtJ���,�8r�M���<�Xh��i,�292�;P�߰j@f+�}D�IR��G��i6u���˵|D������-.��!��L	���@7��F���Ǡ��N��$Q��P�\�� g�V��(���H4
��m=� y�gF��4q�1��>!�" U.E�\	��$B!æzA.�IO�A��+�C�f��,*�����܌���d(W��E��h]Ш�ja%�	r���S�M���M="L�����K%��%�0pP�����|P*��+o�0uZk�I�b��Qc��N|z�Omɟ����x��v:{��;G�j�$$��-��/�5�|�q$�l��}h�p�Y�}���g���$��@��Q�^��s��-���f�$ ��mk�:�S�3G�ӿ
�4�R{�Z�#�<�4p#�W	)����v�w�/n.�}oC�;.����AC깯n�(J����Jx'�A#�f������R
�.`�ٯ�%xY�	�7{�G(����ۢ^Eؾ�O��L�~|�q�ySa<�����a��r0[(��`*'�!�V�Pst ����ҚW�7ޝ@�����MY�??(��F5���0��)�z-,% �n�9��)`6O:�d9b���=�ֽ෼���!���zmgA^b��f�$E���u����K([�p��K�ĭO1�1P�. �F�_��@/��fb�� B�51,��Z	5���sg��H6��p�-b��E��n���A�%��t{�RB.�Ճ�d?��*' eJ�	�l{�d��걑s��.�O{h�yY�<���[D�t�0�7߂u�P�s��N�|��ߊ��V������$���������?��@GaQ�i�H���ˬ���ѻ�uƷ�p��6���KM+�!#x��N�E����r�+�M^.���bͪF:/���i��s�44�B!T3S`�L'���o2��PS�^�z���#p���#@o\h�8uw虥��<u޶��f��nk��Tj]T�z֫�l�t�.p����[�z��~,��g���fH���:�V����d��B�E <\|�->%ou�"�6��O��W^��v\s�4��%�¾������-{��^jA^��,�=z��Pg��t�m�E��:����f��:��ȭ;��)dL�/�<�2�L�)�+Z����G��ұة�W]�l>}�3ɱ�����C+���M�+��nXCJ5��_g�n�i�
�5n���M�C�~��K� 4M��K��(�5�O0��v�z^��q��<D��G�� �-m��$Wj��p�ot]�:��1��]0�U'A�*W��{~�8�m_��qq���
������9�^������˳��x� %.?�*��Fwy^�Hԕ��8A�y\p|m&�e7}�j��@&���K��7խ0���߫�T����7�<�`:�;�z�y����A:T����߿��p%n��˿�����wf?<�QO�5��T��K F�±�����j,�,���9z3���d�2TL�$������%��ܑ����GU9q�(~�>oC��?�饭���>w
@���jw�."@���K'=���/0�&n�1�o�,��6��9Yn�U�����/vm����^7䞘�zBMVꥍ�{#;S�tg��3 �&E��ظ��]\P�d}�ͩh��O�d�c�[�ܿ�F�C+
�����5\�;1"���!,U�Z���(+N&=�k��C�oN��JH�����AC8���P�Z��uz�-��wBug��R�t�����7DKV9 M��/�t�6x�hu��<
Y�}��Ѷ�u-ں�@�JW��ԩǏN��C��'8xZ����Tt��^��r|����_���,P��M�P�LX�ӝ�k����
��57(�i�ڄ !�B��3���ȫc����WjQ�bt��;�i�-�C�>����Kq;�|C����qʻH�<b"$&�ޙ[['<\AM��3��6�fi�I?�'���wR_�[D$���{7�i�>ZFȲwKW1n��L��;�+}+E������=�փ�Ƿ�����気r�h�����[��s�5�	�D�@$�:�0��m��0nSƾ	�Zv|����X�F�Au���.����K��~��*$&��w%���+ۼN�G��5��%a	R4|<�.��8 )M��&R�a�>�J6aFK��9��R��A��B��B'>����¸����w2`��u�^��]�O����
3�z�t��U�kM��z�I��h��CA����u���G�g[��A� ���B�v����ު>��w��������b׻l7 /1���0��&���3ݎ�y��`�O/6H%LN����ϊyB��ʋ�	�ֈ��C����z"�5�/��!��q��s���v����?�:�;w�=�d&�8�g���99c򲓗�h/��M�H�f`�ө)?Oz��+��~\�$��%� ���w�V{���e�S�K��l*��2� �Dd����L"������`:E�����x���a�U�WuL�LZ{�+1�Kf�T8�^g_�> ý��L��D�4����6t�Y+oC���z$�
��{mA���:_�9�)�C]��-n߄-#$=K�[��zU���a�AOz*.0� ��
�з�W�^��-a��_7�zo���x�9�?�*�ȮK�S�S0��F$Ug-��q�&0��g~^�O[�d�Eq��a&,�GCL5������Ael��c��n�5pFz,���0ȴQ�+ˎD�X5��A�i�%�P��m�{z(�|��x���,-��R�7�y���ѾR�s|
.=�y:
�T�1��ż�:�������u#U&s����V/�H��Z}z�:N8���UP�<�S�o��)F��p���G֐se���l=��R�6e��D��bE��fF4��J�EȎ>������g���0�\�*�&����=�e�B��q>�Q:�2ТtI�����q˻�*6]�pl\k'G�f·a�Ե��	