��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����ao�����/M�R-��TW*l��T�F]�{�UB�ͦ� O;�xB���0|C'i�Tc�w�����%����I����.��b鿼46���ZR�HH��5`��@�����b�E�����7�[3���oi����-ؽgO6c��J��{g���dвG?�^ʶq��-�>X�q��ǍBb�����¼-�����G���$��^IO��c��ƀ�74���$��}�N��d��B'�h����G�����4�2��覀��<���0��QpY�nm'釕k%��G"l�~����q� �M锂�VQ�����0����^�:�@Cۭ��։YY؈1����2=��o9E��ޅ$��Vg���<�w(�CR|��5�?����R���C��L�bt1�o�<�^g���%�hEe>��bid"ez�)�5c_���X{�CV��~�(��5[�ýդ(`�dR�a)T�@j7�%^�������>L��*��w�]K����W���Y�<�n��J@�G����3�@��АP-+�� V������m8_�Jo�ꭔ�"gH/K�jŞ��aRZD	m��ս��@1�]���!>�r{/kS.ja�2���@�N{9rc}�8��$S`��Hb{����{�w��p���f�AmQt�����~MT�E+�"2)�`�=z�EQ�F�u���[�;-�O3b���$� K ��h��Ngv[��9� �Y{.$�.�R�I�M�:伣V�`�	z<o�^Z��
�r�5���mx����iP�]+$I�2 o޶Y�?hP,d��IN��.���M;�?�E���C	�MVFJŢ����ط������퐶�Vm�j�\)>��T�������)�n�����q2�p�p�`�L�	��=�Z'�f�5֎��x��
����u(��3KW���y�X%"�UBz7o��\"�5��[�K)Ew%�I��"\1�v��v��R�wG�;�:;��@�i��hm�B�0�j砞���@?���:�Т{���1��(/׳����������<�]`!�.R�?ϱ����?�Ͻ��p*��)��958�C4P��tM(g�풉yZc���R�m�k�1<�����c�pu`�T�t�-��F/_�*CH�ZEMo��<"�iW�ۡ���<�Xru�Bnd�kgi]���������v֚ւ'��n�~aS�0
��F9����ˎ��g,�������_{�7�wn��և��@���%��j0��x�����sf;t=f������څO���LN(!�?;?p+�te�l�}˖�(G<�W�8b�=�?�¼
:۔�sYW{gzO��6�Q*i�R���6�ľrE�?�p͒��@���-\�8���5 �}\}=�X��~A
��@�b�%a�Ws���#��'=���v$,�l�Hg��t$&!,� ���>��U·}��j>��HRr�E�
fp��q�$P�c����8���U�p�o���:>�u"��_��*V$�eK�:��|U��\�8�y�Tr���]�f�o�V/���O����`�/EL-j,��7�@����%�~����kS[� Wo����k�'��)^]�����Qw� Q��A����<L�s�fW������ ��ƍ�_i�Vך*��e������rnGP�Λ��J��!��l ��:��yj��mVD�8�3-Z�d�g茿�f:�K�]+>4e���8���`�Y�����}���v���@�jZ ��E��!k5׶�k)=���QE
R߾��^;���(.��������A�T�VpD����L���+�������9.�m��>����#ν�D�U�\;D4}�ݳΓ$ �V���o�W���H �V!)�$�/]�/.�býJo~5Za<�І�Q�����翶�#d������i�N����Գ=�����L�X�N�/�~K�e�،L{69�@Saث�Cy���|�Į�	�/�V�5��!'�ݔ1H�+�j%-��Jڏ�O-jU:_��2[���4KMow��MI�$�^7�\����x�9��M���f�w�!^�)�M��
�5��
��W����XԊ���N�U���')lS�f��zq�Z&LϯQ����;w��g�6w�p���
?+K���=� h� _���ϡ�ވT�`'�Ҽ���N�޷�3��G
9��ت����ޯTs�����'SL��1�'��epI��|C*>S�&�c�����2ksԸ�\��A5���yF��5�d���,OO�e�2�M��W��o�b�rhB�oSہ�,�p�Ńfr߂������_�#�u��v[�w�Gv"��G����¹����z�s�~�1��&B�ӆ}�a����4�8Tê*0N0�i�;���x���^X$1q\D?�ÙrY��籛��l<��C_[�2��U����(5Yb����蝔�M[ R��	;�ZX��I��n�Z||���IN���
�7y���V+p��j��>0��?�b/�|5�����@s�|�G� @�\�*��,��_j�]��b��tNd��a!X�4�dds�S�싡��띌%*Ŋ� :��2I8%l
�;V�ީO���lǟ�Gt&^��-?W�:��uit (��DW�:�-yJ_b�o��٭Ó�4�|�:}�\oXo�������k�8�{��#��q�a^pJ�d��8�~����tc� "�@B�ֺ��*&�j�����W�a�G�X��Md;�e��{$��Ŕ�Su汇(�?lHeTw��ZMc�)\��`�D��!�J�>a�&����X�b!ig%͜�c/��-�Ƴ� ̩��Ţ�����<�-�]��j����z"���%;�H^V�ʣ�5I����|�y���nr��Xh�~�_%n.���]!h�"����P'8�pS����Z���A����«�7T?��}ggh��4���ͧ/���_|;�\�`1��{�[�G�  CG�%x4�m�	�X���ք�{��ic�q�T�SV��4)���,�a0?���.�޿$)�Se�yẩ���'h���"�F��%�h����7K���O�14����A-�;�N:�����a��(�ck>�juu��v���nl�ZdE����T"X-t��<ׂ=`�ΐ �v^�6h�W�5?ͽC�tLr���*�B��8�RY���K<����c%8˒oNz�����[@P}�!yw;����R�Jm�	=���d؀5�p�$�����uУ^{/��=�̥ot����j_Kd����>�g����'��73X�PQ�ov[$�Ɠ�'�L!��?h-�?�:9F<3��S�mR�|����>��������6Ņ8�W4k�1�kE����Q����j�vY���������gR��}�<E4�[hi�v9к# �s�S��7~��!�.��ە� z���"���yuX�q�	�7��YH@��gm�G/�� ��JbnxF���H�{M�m��wtj����ڕO��ɯU.���Sv�vV�+r�\NL�03]�������J�9�s��_�ab����|}�pϘ�_w
�'A�������#�^M%U�B�+�r(�fl��Vۏ�Mu6`��}�]c�7���x��+��*[O\��M�4oBA�M�Q��$��(�H:Xj�f�N�v��%���T���1�l���1�UÍ2}h8���� ��֏�|����p	�fl�Ȁs�aS9��}�E��2��U�!A���r�&s�l<_3��q�'�HX]�+����j^�W�_���a}����M�����ԅH}����k�m~�*���`y�U�`���_CakIf�ܝ��]��#]�����%�V߰��x��A������j���y�b��8/I���ƕv �gT�(
���
]�_
��Gd.���`��Qz@L����Ujk������ZO�d~'��v�u��3i���'�=à�.��
��.2�N�Cx=WʧFn���z��d����&�@P@=Bo��1�(��]��Z�ϸ�v���ڎ]^�w��h��|�?nks6	pC��I�T�*r�����8��Ob����u��$����%�H���6HA���A�`u|s�'�9y[�G�� �G�4P��B���[D��q���?�j��x�z�u?^���E �(����Z��)*�l�w���Z{�>����Do�&����n�����WsvF�o�f��DXZ���� �@���$5M�*+)'*���;u�ٓ�2�z�-�i�{�N�Zf�6�)"�]Ng�j�8�'c��67X�HG���'�����4���p��l'�	���Qaq�"-P�߱!bP��������z�8���ur�`gb��Kq��n������Y,{���nۋ�~.R�s�g�L�g��10ׁ�7���<�:U(��E�� Se�lf�Ժ>��C~��r���1Q��Bdx�Oƃ iޠط�i֦����A�/�f�Po��w��Z��6}���􄶽��PF��Y��u����ٯ�s	,V�/IV�-�X�!uȠ�vZp��*�:!����^�<K~�ۣ��Q(-���`��c�BV�	J�X�*$;���
�U�t\��B���+{z��XY��|ONc5n��?�~���B��={;�"������3��Ќ��۝�Q�x ��]Q
r�
޶%��;��:����w�E���87!U�w��h8��������f�!8�c�0��C"�?-�Y�q�1�2���ͪ�zd?��1&�d��}�g�mN�
@���g�����&��Oʈ��������(;p������v5Y��N����>p�eO3=z��4��\������5~�9b����T5D��'d�7ښ�/���*]���%? �=��*���n�G�u�8[���,���@Dد`�e��+ou�yG�⨜p�_Z��__w�#6���l0��=�HUĄ],��A�M��\^���a����7yqD��ļO�Q�F�+��c�R>%d��ͱ1�p�)�p�p�sȏ��3,~���Np|u$}���Wy-��r�S�}�=�a�o#�76����[\�c�ہiJ~h𜒷��=n�МI��.:*.�}oK�
�O� A�sN�W=}�3�s,��0�"�$�M��A�)�n8�����T{�"�F�����t�r�:���EjJ�� 3H�g�.�~�%�p�92�� �0m��I;����^|����t8xG����6Wl+;��E������A�2�v�\���
�P�%F��8�(�� �(�Hb]���e���J��bvލ``���pr�����t�$)of��PÙ���SonW�\��Fji�M`�.�|�qw��=	$����N&�`Γ�8�漢���w
��=��a����3Fj|�š���9��S��^����t�΄l�b�~=(�!h`I��9X���B䈯�R�6��n��+B$ ���͗�\�I�-ƨ*��*'�~Mb��Jv���)&*�=�#2ɘ��IG��v�H#��b]Jy%�3�Lw� "���)���/�Pv�hc�J�U���s/ɵ�)� ��'��蒏LYl��~#^5"�7�2��ă��N��
�p�:aHkV[�o���_��.khU*���B��s_�"�L����5�-���vo��K�,���oŅ�_8m�_Mu�k([���k5��W"�G-����:����`�h E��'�4w�B
�1Mz]p�%�3Ң9�r���2h�J��r5;��h:!�ި=�M��W�j@�h�I=���d'?Y(C��L�t��\@[)������M���pBC�ɕLCH�S��F�iIA�@gX��+��8��#'�״�kP60/]a��l4e��X��h�]�� ���g<��ܡ:�����ɜR�+��gV�R.�ʚ_�q��G����6=��T�|�.�ecy��uH�⹏�����;�e��pr�ڰ$U/4������=��Z�yU̠҆�M�:�C;\��硈K��^R +|��0�= �T6H�V&���IO�m�z,&�|e���У��8����A*���(�t�b`�@r)�FW�d�%T�c�oe�(�����Х(�kk��vW+�e�5�[��	3���ވ.>�Sb�������~��ζ#�mL�{܇��d�	�!	���ik�$��?d!И]�V5T[,��S6W\�g�<֤�,=qAn'a����o=M9���F�2����#|�Ο�?�����'� �;��J2\��X�=�����s����^v�����M�t���U��P�4q֜]�,Ӽ>��O��ޥ�N߷ͮʹ�RyJ�hȊ����-�MDjzp��x��;;��f��rLк�TF'|�Y�b�AC�q@��&F�~ej���VO��x$��c����y:�.h�/
p��;n�k�1���XF0\gQ���d��b	�+B�@��X��n�0�"�?�ɇF�y��ţ�Ch	�O?���|�k�Kx6�����SX7���P��s(ʵ�Y1_g��k(,`�iEx�W�z�J2��0��g��Q>L�����J�6���"<S�����*ޚ�K�C�{p4;�7�Yvq��#1sb{K	��c����;$�=.]5�HR,��4q�<�
�����,������Z-�С���t�4�Z,_w�ئ�t�F�"G��%9�3��殲|�V�llZ�O�jtU#P�`N�R#���"g��N�_����l*��&bisg���eaA��N�e��7��`M�]
A��tk��Qu@\8#�����۷�B��|S��S�$�������]�@��2U*t��鋻�ƽȁ7�����qNiR4��r1��vD��0~����$���ى�[R�{C��~>A̰U�T
r8B���`^��0�`g��Y�6��&����X_�B��"ll�?�\��a��*��d0RnC����_h��!�(�&Q���Hi�{��)JǶ�H �3��)C�jz����p�F� �3�cs{QА7�ґ��0u�� ۡ��/k���z�k�5��AR�E �`״9�t�x�n!�L<Ij�f��)!:�$�1�"2)N��}�	Q1�����R��X�Gw�.���B�&F���*�%�Vϟ4yD�Ć�iX�Q����N'5���RMy�'��b6I	�Qc��)Jnsg	o|���z��օ����
�Z�`T_l.v "���&�箉�ha�e���1����U�Wa]k��k��E�� ���b�n�cP�t�/��'W��׳�m"ƪ��ұ�iG��3TE�^x�sжՐPGJ�52��t7�5/�hd�@�q;d��!�0�Z������(�Q8�f�P���鞠!�*)�oل�7�%�$���Uv:��'h��	s�0Ta��է�cR V��� 7��,TF����y��\�IH���ވ�:-6\���8o�Sc/46�s[@Xܚ�i�@-�`(��y�͢WiG�w�H�y�諓5M�4~���{�����Ҏ���o�F�6!B	{��\.��%�C�v��%��	"(�"����S
�|?�g/�`U[C��*�G�E�<\}�2~bdIs������Ǘ�xa�Nia�Զ���HFjІ��'���B:pu���t2鿩|	�A>~(�N�L�Jb �lK��g���j+D�U��S�ܨ��aB���e:���?so�s�d����Й������_���6����z��5�A�^K��Β(��ٺl�F>���|p���^�(Z���0�X���]\�0�Q�-�	Y�d�<v�z�����N�Y�v<�I�pZSn�T�^H ���_�R;h������6U(%���y�K��F��
����7���,���^��ԋ���뗂��`�fj�7���C���I��F�x��z7��s2N��U(�j���xe�-L"������p��21v3@9�����w:���7Q.���ĵoK���U��w�.b�'�#ђ����g��"�,S^L���*U���M>�����Y�Z._�A�񞞰�@5ʂ�	���4���n���f�}SQ�+s�9��4m���cw�ul����t'Gs]	�@"���i'jR�EV1�M@��U�NJƕJ�������$�}]U "�|�%3U�"B�i�^*8��[�8%ke[Sݝ���=��t����Zx�~�����v���a��y5�(H�CfZ�WkbT$�Q1�p8
^=�љC�Z�IS��_�\�fj�$]�W���os.t���gn�g�l�?ʲ�vA~��@u����E�,�*�0$X�o��sF.4D�l8�T��G=��c�з®�g�8SWm�KTr�|rV-���Gg"����@��.k���$dF#8̵����i �Y�h�iP���0� #q���'�r��l����p7�©�� �Q�$%������}���ݷ��B[�d�"q��i '^�2�C%��6j3�-��~ �$,21�wU�03L��T"���n�/�%['��b���P��[qn�j�IT ��Ok��ݸ!������|�x1�="�+48*�J��X��p0�B
F����D���0Μ�T2�k��^�8����_�bmB9-��.�vd���a]�OБg [�`�斖�>����9�	�E�K���
��Ru����ۋP
x���9���US�/�O�W~	u|���	�;?|1t���՛`AN��`l��ā@y�R��xEJ�]���9���X�!�$�.�{0kwZY��zh+��nɮ\r�C��D����O,�� �����yk?ZY��#�PvBh�x9�]y�_)�����7��땫�&��"��E�����ݤY�~^~G.$��'�!pk{C�)\o|CxnpU,{�៮�VG�#R!�>,S��!H#�(�=��+A�#C��#c��#*.wtS \%�y����̒wAʋ�Y8��T�;�K�¥=�m&A_���_'�a�*O�W"_��U�����ټ��yC�N~�]�d�֣L�<��br�IV6�M�f�죸��eȁ!�����2�L��#�ݻ�Y�����C��U͏S�͢��u�n�aH�������+/�C��Cu��a*�wl��c8��D���Vڞ���x��SBe�V����E����>B�ǋ|��*�^�� ������-�p]-B�*�8w4Y��T���gH�Xz�fr�Ҕ�)��:���0꺢=v���WP��(o�G���G	/s}�	�r�%)��Y3^�ߢ�gD"��C��I�m6�N��#�%a�=���ư7�J2���\�lki��2�+Zf2��l+ǨU,H������;����")�+�Tg�(ŏY�n؁���8�~a�]�1#��g��U���T�2��꒚T
>�*�d�'Y��Q��80`�V�ٽR3�jSH�����~��jŰ�n�H��$���s���;�Z!��~;���L�Vc%��h�'T��K���iʰU�ƀ�KZ�U� ��Y1ӛ��[���5���R
�t��t�;&m�����--v�\ ��U_ЊN��*Ea��������y$�̏�]깔����
����Z�!['8C�?��ϟ�����R��h �!�L�7��C׋�y�rIS�h�/]W�%:�T-�UM��RA�7<t0���k'�G�£}X*��H�]ğ;Nފ��p