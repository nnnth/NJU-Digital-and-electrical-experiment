��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�_���v��	�������d��i��HO�4�H`���ul]����_/�ǣ�����J�g�����������Y��� ю훴�"��A�Fb,j��,�Qq���~G�4Nw���݂M;�g��X�}�}Y��PZ�?�������뇛��]b/��ad�b���Bpgp_;�Š�w%C�X����F����3�$��1��N�T������~|4^ǸE��7[�|�p���">���|n��Q���a�,���=�ٖct�&�` ��X�#`}�c7��G_�#� )!���P<0p� ��b0k�dϷ ���*�\gD<1~=U>l�f����q��V�_8��k�D�9M&b�e����A����7�6�H��C�WO�)���i��Sn6�<��0�Ӹ�B.)��"���R���� �e|G'��Ʈ��d�ʯgqPZ��c�m��*q��|hm��~&�د�&�6t-eO6
Ӷ����@�D���ch�'��n�V��bM�pS�p>��O���R6
j*\!�O��r���N�s���Mo%�#X������v�$Z����3��kY�"��(E,���t2x��, #��6�����%�}lS�/ ��{��Z�4��ʈ�|�l�V�8=U�*8+ˎ�2�c��;�
\Φ�:]�"Y�+��yqx."謧�(j̯�ԝ�k5�2����;h��9L��IC�OQ�j��L����b�^!�ըx}�<�f���ڦd|�ҋ$��z�@X�o�%��W�c}�΅�bCj\�s��Ł�T��/�E��yy6O.2��*�#���׷�h08h��P���t�sn��qQ9�Hι�`&K�\V~��k��$~���kmތ�w�͏ާoX8
N'��� 	��8{a���X�bҡ>���I;Mf�]X�uox���sv��i�ocH��I2q����O8<�P\�C��#j���e�װ"��IБ*���M��{U�jk|���W�?Z�C���EwUt�����
�ȗ��M��H����ΜT����#2�a`T��6�T��A�E%=@yDM�,�x�=��Fn�6sy�BC��`��vB�-�ǰ�R�MlJV_��d�a�����{�l����j/
��m����k�Y�7#z�B�̟���s,�|�v,��f�mu�"(Y%ݞ�uz�Q/8zd�O�7�U�4�^R��M���/g�&�lH����=�mo�+�`z_�)$�K;	�k����kuO:�6�,���&�;�
�{��~����l%عa����d��V��'����(���>�3M�Jj��r���T�g�F{M�ϝ�%��>;�'�+�b���o`��(�wJŎ�ּ�6^�����m����/Ԛd���4��v? ����΅�]��*P|1�C��̂ Yԇ�`��Zg�B{�e�ͱ��J<z~:��Svhx�,P��4�;��A\��|�`^%�/�o�3I���@ V�yU�mb(�f��))��dl#hFsk����j�	wj�8GXP��g���{779�����l���2�0a��i ��.�+Y
�kc
�eSL-����q��X�I�8�!�������|������T��)t���i�R��j�U��Lɇ������;��Z@G���j궶eX�s�S��Q* #miY[{�� #�|��Sì�B�E5���Ю�?�I��J�k�����3�����7E�4`,��H�����;(j+됑�Q���QO�#TjV�������G~4���^���WW���|"�#'�&94� �,2n��?�����Q���$���H��:s��.nUsN�$��(n"�ou����bEv�,�$^�e7���l�J�~-)�f.�e�mFZ�x�x�<��SñIFx���s��?�Us���F�^��>J:2���#+�o��x��X!�u���S��ϫpf�s�Dl��c��-��u�OɅG���o̊v]M�7���RP6/�^��Ǘ� �"P4x͜��G�zcS��>ԼoI����:5�k0m��3%S�uJ8)y/|��Y(H,�9��ة	���e�������T�8��#�Z��2���6l��4�/4z�F?�"�s�<�V@{�>�7*.��Ny�o�����]9���)�m������1 �ſ��-�&+�X@�|7<ہ"Il�Jvk�^�3Ҡ;J�OR�I�E��Y�.�ax�� ��i����c/:��}�p�r~p 2�wA׀b����a�~�A-�����Շ;u�����$�9��G����o_�:�G�
���q�of��ܰzu�`ְه�
ZE+��{�(���4b�\���'xOx&U���nv�O�Щ�\ #��o��~�4+KP�ƽʬ�P�@�vrT9�ј�ۼd�yU�Pt
�>>G�h�*���p����)��=�f?UѤ���'�U�iHBz?PV��Jj��oT2��)"6�G����X�^QB�6r���ʾ���N����w�q���ͲQ�6�e!���:k����2�-@�3K��X��t(f��{�� k0�p~�/�i���7�s����s����Y�a��/.Q���R�y�ۤ2�������&BIM"�Ɩ�e~"��[�s�����5�❵����5r*)UA(�����1��g���h;-���M㷼��Ó)e�h�>��/Ф���j���p���%o����Bʎ�;�8��304��%���r��ʳ���-@{��S��Hø�0O�����$�WH�����{[�/���_A���`�`�e쯔��f��v���!QW���+���ؾ��T�d?x���p�A$��zt�p5�[P��
q"d�ο/��-r|f`N�~�RMu0�Rt�@�߀�)`��r(��9�)K���)0�h,�Y*��,@����~�O�\�����43�۹�!����C��DUk�m��r���p�6��	@��WN�i��V�1:D%��q��B���TMK���5��$�ۉLc�f�*3���N��Q<D���m��^���g�@aꀳ1۶(���??IJ�Z�F쳐�}ӓ*��V@�L��n�hP�e�%02����t�6����Cڸ��/#h���h&�����'G�`:�@���k#�xQ�ebL�f�R
,z�zö�}m%R��K����a����V�fd}�C'��n�_��"#%�[8��]k�g��~�2u��7[?���L$�����ǔ[I�uU���I����v�s��М�]mʂ}
#E��\������[��� jD��Z�V;/n�G��1ۖ^� �B6V��"
���8e�~v��I��!	�(��{X���ܜ�=��M-˰bM�Ѣo���Y7ٌ�N�:��###�����s#��f�D�S��ejUa|������������2���+[���[��֕c^ C5L3������6ED��DY9rck03�æf��$�a�O�]��.K%�no� �j5�����lK6�NK���䗔�-y�D�(O�0��
|-5���V�p�a���$�����g;w��
�CV��R:��r�s0��ղ.�[,#
�
�/,3P�h֩�F��4{�L��F�؃_̺�K��a�ɸ���1�tlA�mJ���Ս�2������t�\RW�x�����3�G':W}�?ǈ?xE��܄i|8l��v�eĦ=�:��1�[;7mc3��[E����'�?3�o�R���w�� ��8#O��H4	T:�lಊ��m�Q�K���[y$��M�S�΃C�7ؓP����1�N�`���4����3�?�+�Ώ?�am���T�`p��g�5k1r�"�N:��C�V�}�&L���eW�4	X�ǟ0�m��h��W	O$�� ^�~��:.+�[Vka_���
Mz�)#>�V�߻}�L��Q�t�gGD��-'8X����@��L?�1���a�����Q	��<����mU���i�^���4�<��?�R��l�*�<�W�Z�dK�-ʰ�2A��c�:P��fB
�r�~�_J���ugBmH�������,q�T�Aԑ�?Xr��f��S��>��K`��r�%�/#��s�K�F ~�X�I	/Q�7��Ř$I���n0��� WN1l����ˬ�@���D�d¯�R(_�ҷ@��v�<ip��p����d�E��O"���3�$7>l����G��=�Z��ᇊ�L��L������|;�1���9Q������&��nW���Z���z��Ұg+��hJ���4�k~�]�*�W�pZބ���i��(��i- DH-�ӥ�/�A�Z=;
��qi8�
�l�ٹ�S���!s�2+�b#���,�=O�@��fDU2^0z#���ǫ�����z>��j5�ܵ�<��ꅌs��TnoM_Ҭ&3	�Rz#����Rލ�Ľ7
�R�9�B�vر����wb��<��(��6�T��v��0t�nW��/�C/�][�%� ���#'�(c~n:���;� �������]��})�K�k�G���� 1r�n�'4����@e�#@";d�:��>D��_�0�/ &����}O��=�䀳�@Ѫ����2%���V��g�
���o����b��6�m4E����wv�fVB&��^/�z�����l+�C4&����*X��&ڷ���Ɩ�6��{bO�!t'����B�L��6���5ۙk����{e����V�Ep��qw�f�f��1ޡ5�%���L��Tu�%_G}B-�D�qR�CF��?�H�f��>h�VR�B��A7��P��,-h��
H�/K�:x�P1t-�r�&g�=�4�eC�
�<g�þɆ�J�ͳ!׎�	tY�y�b�i��$�څ�l��Y;F��EȌqL���
Wzo�34z�
N�BFm�P�j�zC "������Ԣ6����Kj��z�Y�e�����q��pϊ�3��Lx��`�M�\�w�R����{lu��_�ro�v¥�n�DB�?���0a��6Ɏ�qq7��ʪ�9�C�Ͱ�{�J��Ӗ���F4;�Z��#nweې�����0)d����ӳ�ޙ��M�._³�}5���}����C�'�!��DVE�@z�ɳq��c��TmM�l'��+~Z���ydm��lKM�ɖc�"��9����sJ\v��O��_���P�{��w����EV �G�Z�����;:G���q�qn�G�`6�{Ԏ��m�;I�;^Z�y�%}�ԣ rω���͆�`�����D�Z��㐏9�X	��ҏ�Aɜv��$Z����}?Z�%����!!��s|��l9-vw28)�4w���a�AU��n��ryN��Ĺ*�?����!�ք���s���r�#�v:H�P��s_EB�?[־�'Z}��Ə���si�?U���1��}�_O�*hM�ł����̄M�;��W�l�s	����]{��@g�{�z"1a�/�ŧSE��g3,�4=��ò������	{&#?x(�e���_-Xţ��5��~|��zkI:�E]�0���6̀j9[D�jT�ס%H�ԉOG������)��	�q}'�R�e��ց���@���a쳾1�!OBZ�#6˧
��K0Y��qo�(���&���q�;�VR_~&z�/3�w�KF���}X^��㶒�\r�	�R�t<qKJ����lg�����xϡ��78f���3���.��F�`�9�PjNk���~��E�"���C�n���p�#�NhS��wP��H��+�늗>��p�MQ�H�2<��x�AіYu�J]#J7ӮȔ��09H^�)y�'���G�F����D���3�B7`D �e�H��Z�i_ܿ�cȑk�O�`7���5;3,!��)�7�U�Wq��ʿ��ٸ�6�yx
��p(4�ji��
xဓ�R��j�Df���Hh&9� ��؍�x�;�m�wK|kg��̸��ԫ})JȠ�ծƅ�C��ʋh� ��Wl��5�e�7Ą�.���Ĉ���}���<�X���c��
�t|�A�����B�o�����Z1�vT�Q>�-��O����z<6rW���e�9���p�\���4e��\{ �0��$���֊�ڔ=$�����E[�2�W���lo��y�	�j�߁.�]:y@���w�%��F��#�l��r-W5,�x���
��hK�4(e��[�^'�}��$��,�|s��K�.���]�yj U���a��abLbyF+��u���|��?��xH��]rS��m����5�6��]yd�;��)��S�0C��Q��6����e��`�P���c7�nW�!���73ֺL����?ٚcȶ�;��!$@�D���|Ya�`��uX�'?�6�m(��))jN�z�7��;��p<�~�P������� �+į��7�)�+�iو�4bZ��S�W폱�^���x�	��`����/��&�l��J��{���:���V1�K-N�)�
���s~��� �	�@��&|�[�ċi돮õ�RZ8�,�S�:�9K&��ǂ�5��@x�5�_矧���M������[��>5�J�F#����2*��6����=Z�ilI�ѻ�Es9ʽ��q��MK�-+�n������2';v0A3.ĴH[��������c����n��ߦ2�if��@ ���;������.�]eI)JoT9Y�%m�� ]MҷT%��'��=@\�M�=�y즔�vlK�<>��%�	�i�1���?B�@>^��#<�s��1�J�x2�=����XtP��W��'��/N��A�%��$^�&����\��ĮЦ�HqH�·���}tՕ�ʳ�S=jvɄ��s���ðq�T0��I�ӡ}>Щ��#C����|.��B�����D<_�\�>���b�:;w�'�"K	`��X]��`��ecsݦB7+!M���&��s���p݄�d�HI_�%3Kԫ����r�o�(��H��T�����u�<_7�P{фі�T7w���DY�� l�w)G�~9���f��,5!y���׃ ����>��{M��"܌g\�B�����t_��F�c(�s�S�y�逳k_o��#p��t
:J'��M��yr�u�wt�	.c��"{�F*i�z�L��+��H�%��d(�7 W��L��d�$B�w;�fҮX]�*�uaG��c�9���,~#�m�ŹY���.�N�L�6�-��'ml�B�(4	��웦]��>�"`,�ZP��w.��F�3���t*boo�tj	ݨ�Ώj�.��s�Y�?��{ת��+�ɤ�w��0\��߿��%c���YQ��BI��I$>D}𭪳,_c��io����󹥂@Y^�[�[�������V`苌!��ؙK	�Oyl�[��l@�ζ���V�,I�MY֡��Ջ����ر�'ͬ
�z�k��qbB����W�w]�|�.��ק�.����Χ2����Q��@�6�w\�(��P�hgi^e����@�x���ͅ���˃p�����{����4���= t �VBI.<�%|+A���_��z���M��Z�ًZ�u���r��x8��g��:*�.s�4��ٟ`�[�x�hS�|�a�MV�Y��B�jg.b۳*� wM�0��ߴڤ`�7�k%�u����k���R� ;~e����ۧEAv�-���H�f��D�oy^��G�j��w��ԛ9�}��b V[ z�~��:���Su�̯z�m���-��GB��Ę��>���Δ���<H襧ꈈέJ�*�j�ya�!��A:6\9�
�,��C��^�@�$�rr��v8<C��-�Nq><�����$	������	���@¥A#۾o=���\��O��9R��0�'ouہ�3��)��,�p���{~���N�]��P�<�3Ck�<�ư��^0L�89�*(�9^I{�-j���1C`ι2GL�:N3�����D^�\� ��pF�=.BRM�yw�;��Z�R�FM��z�Z�-R�B��$�ᮥ�[<��bfR#OŇ��}Y�u�(���������y�_d�%&Hފe�j\�\ũ:��e%W`�
��]o����qi����Í�\�T�+�Ԫb��d�Y������%�~a6��E�Pob�!#s��J?/{�0��%����ٰe�Y8�*sfwF�ӓv"Q�0���5~Ȕ������H��X�/�5�H4w�j.h�&p\'(G+�Al��E�[�c_��ٴG
^�ڱ���u���' "0���(���X�)a�x�d���c��!��	h᝕�k���qU%چYI��@�[�<X9�,ЁDv�jR�g~�[�8W_�J?|6ƽB��V,F�+�fc��/��T�zs���3�D�0%���ws�R7<$������j�zYc��hD�S����w|u���|�[���~:g!3W�OIܴƜ&�P~�G�5(`d'��/e7Eug��JȄ.�9�\-^��+�IN@^�d����m9\0k�|�x���_<{�ۏ�݇B�r�y]�-l	�m1=��Ul7�����~ӹ��p��k�*��λJ�+��?0���(�v�1v���@���ytwǎ*�3 \n�m;3#m�2#�}��`~pg�U�8s^�X�.�k�n@�
���ŵ���Y���34��~�'P|U�AtD�:"��=�bfo�N��?����6�	 �-������; �=b+B/��D�ZAyy���z�<i���*K�n/1(`����Y���V$��[҈���9XG�]J;c��EǞ��~��讓Ķ��� 
�0�B���$�K���M�
�Ié�V���Іu��܂��#^�_��G7���EN���	s���O!'C�A�hk\��Fۊ]�n#��#O���gi]#]�4GpJ�t�:��o�O�6�q@8��Bx%T*�nw���r�4���'K�My6��<����7Q�[�2A@��^ٜ��=���{JLr5�Ui2�
�*B�5F��j���C��3_��'�>�)��3��9ań1�s�`����E�*u��~s$�	�E������"�@]�G��i��Zᓺ����Q��A>����ֳ��WM��ŗT5=�gl�CW����N7�%�"����
�[-�#1N��4�,��x�%�kG�H�e}��̄�ՏST!-�)�h���E鑯EǷ��]���RX��]����T�fU�bw��!�ty��_��Ư@%��㍦�[�}cHYid#~�Ȥ��У.b���a(x�Et{��[�O��U�� F7�?��#G��;�֡)ٴ���5�!Mr"{��_���!��S����x�=`�r�:�ش�#F�v ��)ʼ�-����a-��*�CM�i�]X=���T)ol����C���n2ڮ���?��������(�=�g�'��k���U*v��!d>a��_�iFI��|9T6D-��-�%���� s����ʉ��T}�l��7�����N�����bc��!^*�oޭ������-���E��0��[���v���f�w����Eqb�./|�����U3d�����+ҙʘ�e���zO�c���Y�Y
M���/f�Cќ�G2�g;��oD�[�x0�}�uz�q�~Zh���2�-[��FG�B�N2g���V0Yq7k�xl�Ǳ�'��{
O_Se�[�����䥨��2m��u�(7�2�=�i�M��#C�ʣ�����$�"IW1�3F�
�*:��a���/Wi5��1�DS�	_�-�ɱ2�xc�!�ݮ�M�<:|��vFM�UAJ�Z�j��@���Qj���È����z. ���|�Hd�p�i��cC�W���* 'i�����2�(V <�p���?���� F����Y���r�Aܱ�rq�����~|��&�!q���:��NiR¡^逭ۀS�S���N����Х8�/��E<N[�d�mΪ�u�wM���X�b�8G'M�N�4�+�+$/.#������D���{G
�玝����@��:9����\����r�E��;y��Z��6q�Nr/#��n�,�^�C�S���D�cV��1��'��l�U'�O����<e$��>���� ԧa�/髪�w�85Ǐ�n�0������܎�Lnb�z�����$P�����W�~���q�N�C�&S��JIp�d�좩iT��V�)���{��I��+2�V%t,�����Ġ����>��>tp,?Ͽ��#ˊ�H~��(�#������ ��� ��V�Ubv7G�[EJL� ���%%�G�q���Ι��)���_��f���԰�9��o�(��uz�w����^�1d��ܺ��Z���Nԛ�\�bJ�I�i�R�v٤~)�}JZ�",T�h�{��,��7M����n�����������]�qè�!��ڈJ��s�S�Z!��u^���5F�H�F�$,�H�"�(Y�@�M�Y-��/΀1ǽ�ǈ�� �����s���ћ`�6
�h4�m!�s��r�M~��,������@+�\�� ��|���V��Qd��A�OJblFg~����ҸAV��̙Ͼ{�kRr4�T�2Xb���q��αg�2F��7�)Q0HΨ��2���6ң{�oe�k�.3��T@�0\Mj�$A�X���X���h�����g�;(_TVd�w��/P��|Vd���u�x;k�u$*O�@"�{�;������X�u�!`8"��fV�����Nm�.@7�/y��l��qN��u������m�v����i\��bp�F�G�Gc?0��aX����&��c�{�^��D���ñ(e�\b�f���xJ�6�F����7I�V{�*�)9h$����r���xiv~�D�#L~����e��LE����^���7r��0�ԋ�{p ��d�����<���Qq� P�D������$��iP��W�T�y�&V!�;�����|��P0��;����E�+v
*8v�d�r�� 冬�1v�-(�i�E��c���3�=���E%Z��ȉ�'�}�}ݵG�gDNf8�����=��|���>������הOdOP��� }��1ݽkh����)��->���%4�w�/Q�-w8W�&D�G��R�0�D��4:�_ĽBqIH�ɏ��,H��&?v����,9G��RG>L���\�s)���6�����v�.�������ɀ(��M�㔌��6T�F��g�%�ųF���ڂ��UN�F3&?��cL0e�%%S�P�5�m������w��������	�ˠ�X�M ���	�����L!����_\ZWT�7�}&�uK��v�bE��]�t�E" ���@$��*��h,���_exc0��L�%�8-���:��g5E@��@c�Ä&�~k	�ғ�LZ����c:+��(����\Z�*��Y��8iԜ>��l�v��&P��/��Mg�et6�r���\z?��QR�����J�]E�����/��n^xI���y�[e8d�#��J�0�'@��j�hJ��$�KJt �$���m�e���36��Ѹ
2N�-��߉��?�?�V��c���?�fŠBH�����"F2>��~�4��W9�J��}-�N5���4�u��ܛ�78Y�!��M;��L`|`��Ya����\�2�Ȕv�t?�	�
��r7�(�l��~����1N�����h��W�)�u��`R~SRƓ�:u�}���k��`]�B���j���E�4Q�ቛ�N�!r�P&���D���A9��:�5�;�DX�W
����LqmU��P]/�$,(0�ԵK�2��TUr��-�;Ө����ߟ����d�JY���8���7ߗ��]���6��8J,�y�z��ǥ
���c-;n��F�Yk�!׀�s�u|Y8I����z�L�d��z�<��0�����'�[��T,���%?���t�\�I�"o��47�fP��2U�te�>l�a~o=%�1Ng�/�E�>��z8g�C~���y�=i��M�E��C��J��qA���Sg$hB�g�c�F����`��R�1r|�~���I���S��'��R�t$3ZO��d�b孌^v����"m�#�(����:e��	!�n�9��9r�����p�?k��O�����gx�4��*l�U�;�r����&u���S�1�o�7�ں��6sH��P�f4�w��F�,�$k�eT�O���X�ʉ���y&D�6���¯tsy��w_֫��X�0��O��L�1����w���C/o|���5'_�<܁���؏�L�W�ނ����j�<?�}9SB��S��7͂&-҂���_�ʪ!� @�"��k��]�i����M��^�^�G�
q��I�J�%�TS׊l�G�pq�Ȇ���zF��"AH�B�l��&��ɑ��c�0|���jfRlI�N����N�&P�5�U�P�M���6�V�=83mn�L�ebr�Zub4�
U�O����]̔�ܡD��&��~�h06����5����%��`�Iq��Huf���kk����oĀ�T�\�d�$��=�iE�961B�t-(/��I܋Z���ā���@D����u�KqL�����&Jf�����9Xpq����Oix��S��E���
M4�D��a
g�U��q"g6�"x����&S5��FNS����u�<t�t����J����5q`X��^��3���81`_ Wo�L.mV��XN�.�j��]�T�� (����P����mr���w>5��I�]쫐�:��I(��V����ۿ��^��G;x
:3��LE�����aI�Ϳ`ތ�LyHHS/�y��8�&E��g�R}*���e�"���s}�n�Y�����zT�e}����$~Ϥ�Q��C����P>�����`�eY�S�`���x��T
*п��nIR"־q�3SY ����
=V&j{���$�"N��|�����過�L_+5K,��ǌ�m��.��L@��Uه�rj@͇�H�o�u�a�ۜ�6�d��x�|ٯ=�8C�f�s�x�m��g�i(�m^R ��ذ	M_�Y��d��	��4�n?^c�t�*mYG�*s/9B���)w�u����=0��6MR����)H<L5U�;#�ȤZ��%c23K�ZN�h-�D�1��Ls�W��5�j�Sa�C�Zč�`	�y��W����.�6!�{����0ḑ}H�E�#D&,�Q�����RtS�%�����I��f�����.��P.ϩ�_%6vs��\<pR>08�G�o�^�{���Y�D�
��]+۩�w��|��<�$~������8]�s3-�9���������b�>�e4!0����G<�ë��RI�Nhp���'/5����;֣�G��zJ��x�겇Qc�yA��Ī�8S�]���ip2�t�[���/ X]�w�FC�s۰��S��H�/��l��~�L��U(�Y�d���cc81���n�i,PMP?\:&�ף&C��3<�=�n��������}���G�˸[!|��"��ޝ>)�Pu���2�/e��I}���"�pk��,;�tr���)@�D٧J��t~Yj����r���M�575OK,�~v���E��qa݈2k��.�(���^��u�S���I����N�����p�Ĳ{ԴX�r������W��Ly���{�I���+:ʏd�*TZ�nl�c���	}yE8�<	4`��Q#9��@���:����V�$XI����[��}*��1�d�o��PDr�V�Z�SD����_�k��ЈO}�LE�ܙy��B�v4{K P*
��}��FN?�t�.eo����Q�l6ЇUjjq3���1�{�Н��s��q(d���i���ˤ�⿄Ьy�v|Os��/u�Z��G�^��G� �
i�B�Rz�9�2�]l�v�r�"6�ٴ-�w3�E� �޼U	��[^�o���!�j�Q���ar�m���Kka� %𴷢^b�FZrK�i3�?�G�����T5�$�}��k�!s���Z�e%�K2'$�;q4