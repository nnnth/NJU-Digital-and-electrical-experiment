��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�����U�|4�}��3w���n��B�2�Y��Bر�An;|ܿM�MT�[�=��Kv^��L�`.���kS� z@����$7�.�'@y�>Cf�(t�-��D]��m��f�b"��G���t�:���bf�3�%��?�lG��nXI@@�6�~����2��Bt�ϱ�qgc|D�k!�a�����#%�h�z�eNd[_�S����(���o�B-���
��T�!�zvn4��3I�c� vl�<i�Јs�o��Um�M	�{��"0H�=p�0�˼�Yi�}��佖]a�Ǘ��҉�Zz-���&*݈͵�'��\,����u<뮁�ӿze3&"H9��X��|܄1��_�`D���?)�֟iӺ�cA���W+�)�}�11.�1��j��jꈮ�o֩��@8F�V
?�?��5*��k����)i���	�.��2���/69uMd�O����s�>,\�~�,�|�k�P'��a#L��m�;�Jq��$rE��yX��T\��p�'ȉ\��~������PK�S�z��Uu��!�� ����B������&�H��)��z�ӵ����s���5�F�z�
oQ�Z>��Z&%��LV�y��+��3(�����j����/(�F�l�=����E
��K��	Q#��cKaP7�)��T�Ji?������;N���#���	����+C���5��g����@����F!oŲ�|�+_?� (�e�ֶ��N�I{��		��)��68���SH��?ȒZn�f�=��+d}�G�ձ��n�*�tF�qX���P��7��
��#\��s��}�=��V9I�#[���(���R5�;d�Hgs����0�"
��2Gq~���Lf��,�v�i�.v9n<� ��B�STҟ�p�B.�r
�w���N�i��mY�]�֗�Y\=ȋ�Q' ̚F�oz J�TP��?Uhi ���~O��W�:�`�6I�R���α5��Or<�qP�N���:M���*�s�et��<B�����;���ro���#d���\X�T�~x04�}B:Nm3iu��ܽcL�y��v��;��`�ͅ!�=�&��'�J�Qz�n��?��e. ��k^�wb����`�tb� �[������ـ��i�8!���Z�P�7�TӪ-s` }~���9 ���{$1�)�D�2�loDǷ�;25pڼ&��b��YL��dF&�Ĕg�N�S\�Ǟ:t��r@2#'��d�Qޥ��aq�:_�QNP^I=Ӂ3E���di{��4O?K ������C�����'w`�&$��Έ��~��u�g�����r�J@�E��R���9*��d,T�y(�c+�l��0�Bg>?Ȧ�^8�����]S:�A���\}@� d(^'
3��*����`���́!D�V�#��S��@MOt��N��EH�}�W�=<
����
�Y4�-RT��-��BD�s�]�7<.7\O�@n���"�
�>�J�ˏ���Wے?/'5����(�/���Sa���9>�� .
_~�Ɨf󾋪ͷa�VPu�f�ip�Y,8��|�M:��w�k�1�_�P�l��!�4��ͯ�.�#MPLU��$�G�B��P��^
AR ����EBH�D¸�C�ؗ9윬�t����
������������!�b���\?�6�h$VxH��hQ̥��de�`*�F��#1�zo��Z���Af���1��a
zE�I��55�QE�O�4��bA\ve\����}��Z3(�|�;坚a���E~�r����G�d�AL�.���� ����9�6���NB�d�W�o��� m�!Xv�tՌ���3���ZyX�Q���rz�ѽf?��Üi���(d6�2�n�>tpǪ�?.I��J�1V��<�����jh���0�	��H�t���֟1�c�:������̓;G�@|����p�_/��c���F|��iuaHqrѶ �C����S���t�7�T�H/I�U�х��v�ύ-��w��7��1Frӂ���E��#Id#���M:E/�}:~�;K(�-3ޔ���{�[Z��v`++��o��+x� �a�f�;lu/�����u��G�
��0Y$��ѭ�cԸ�;Ͱ�^���a�6���E5L�醵�GD�3q3�#�H�p�
1��py�GLg4�M7�ݍ������=:5�΋���w�����f�sL� Gz�sW|9��	��&����������x�^�
�ⴉ���a ��&�#$V1?�IF��Gy�@�++��Tr�uY��E!��Nǐ�9��{4Zi0;�ŝ��0��&��+,��w�-F#���c�����B�J�D9�@NQ�f��-�0�'f^�΃F�o-d��@Z�
�嚡�R�ǔ�;w�[�����J)�T�g�[]���|1<���;�����Q�T�  �ݫ[�į��풥�/5`5N�g�.�l�w4^\��`��k��j\fU��R�v饶G/8)% o��(I4х�ٚ��x���Ӈ�Bo�|$Yn_T�]g�_�W�u��6=�H�cl�(	��{���ߎ�3OY
�)�Z�+ͤ����u?A�m;�-)��	��S�[T3$��J�V���\[�Ff��X���K���t���6��.�o4(;)�")#�o�U�1�1=.�X��	*�iŹ�h�⹗�Z㷡�6�fZ�f��1�9n�L�s�3*S��h���`�1�kx?��P�]G��GdZ��擪�d��N�m�:���y������J�����tuS���¬��'�_�ux�f�C����yfjL!ο���%�*'I�"�ӎe3�dH�z��c��o��Z�B{��Z9q�T=y��.
B,�Y�5׃�6���(�u-�X?mg�D�ǀ��[���dD��|�'������*���7� �%Li5��x�#�to��@�K�kF�υq�ؾ}�������(V����Zs�lDX�P�d{v�B}��;�ld]&u>�Y`Z�K#����>�:s�q=�"��W��dS�Pٗ:�������w���������a�e�/�q�s�/�C��9���v��cv~�P�p%d^D7Z��|h�|ϛ�y	��R�ZU^�4<���'�l�AJE���ã�	�v3�1N6)��t�ڎRr��n֖���$Ͳ�7��MB��"b�]49�����|���X���Z��-�&?��[!��ńC����O;u}��;-��\��pڴ�K���}.�#�S��tv{���`���
�R��_�,��iM�d�X7�nGk��N� ��BA*c��+��7'������1w{r-�E�x��7v�]�Y�O�1���^A��ϗڧj2���@T��M�w�]�h�1�����|��D`ϡ���TFj��Cm53������SC��[:��v�p�L��)w�i�'$������ŉ�Q��t��ɱ����@5�UFϯ6��l�����J�|�}U#{�P*��^��{v��*Z�QZ�hk<�p�ۨ�����<Ui���~�;�v>�J� ���a�,W�ı�OiZ&��E�I�$�]I��qK��J>�?R���VY{���,���.ω���W��D�ܨ��Aa��vJ��Ex�2�����D��Tv�,�]8��u����+��33��.&��B��Ҙ.>���h�������ڒn��J����Ʒ�t�'���T���%����R7��u�h���6��y��L�&�G$c��P��kG�B�����������S���]��ᇘ�P]��vܯ:gy�fB��[t�ѧ�w�M56�E�S`�43I�`�P��g�9%�o�:A�-��:ZiL+�Lp����������]�"y���#�o'B<'6'H���<�(�`;6(aΊr��r)n�x��>��"�4��<��?��״��Y�7�t~CCuc�� J,{����]�����X�~�!/H*3���J <v��Zޅ�&�҃���Z��K�_�[V�fn�<c;���dn��Կ̋���L�a>BHz��Sao\G$P��|/�����O���[i[@�Ŗt ���Z|�9�7�8Wj���	����E��^��}�A��4�����T��������5T��һQ6L����|�����d��d�"�w#����V�o�E�n�아�B�Cv�~���G�r��#GV}&iS������J��UFܫ뵸l7��J�Q�k0W�/e��7�]���ϖ�����i����~M�_�4����@���WYm.��1�zô'S_U�a8v�p'~@�=���j}A��k8�@`ŭp@��{ ���s�r�,b�&y>]iDi���.3�!�A�����m�b8߻:����ia�>,$V�[||{v�i�@%��'��١nK�:}�p^&��?s�*Wb�R(��\jc���Kb ��i|y�x��=�9��t(��j��������uA�+&��)�wʩ�D�x/���R�A�Ć�0!0��qB*���kac���
���q��q����4�"����ng�0�ɇ���V"�-!:�Z�#��Z��,�M��B�:�������!O.P' �"��Gx)������&^�1����ŏ(rd�e5*-� n�ދ�4WBT�3n�v��~���w���B�!'�%�/p]_���m�,|����@&��}x���ܓ��_�2��gBN��E"a�v7+/�͉+y��n��!ιfa�d�M!�-�JwrN�2��ʵ�Jˌn����_�B�ͧ?�Y� �^u�8d1m3ÿ�����C��:����&S눡�]�|��~�TB�~���ώj�ܧ$�1߮�\�ko�S��!��W�X��Pvvm��0aD��+gE��,ˌ�*�(ӵS\��v��bD��7{>��k�6���^K�oΌx�<�V�^�V�<u
y�P�_��R��K4����b��=ëdU��h�>��S��l:��̶������_�b���*?�{U|#��B���%e,�\f~	s�k��5�ߴ�� J��)���S"�j̊\h�fyw�-q�k]<�Nn��xz�q�[�&.������SN>�\傋�?,�T�M�,i���x�����+F�*�_�2�mƭA�N������d��\������{�5�ԗBB�34Z�V�)���"����'�8\�{w7��e�H��|A(	E��d�*d��b �J��i��e��6WU�2�i?�������)�u���#3�&Pv���s�A;x(�Ug��_xߝ����={<�����Pr��X*��#PNى����RZT��>��B��JFBJ��KB�%�h6��x
�,
��lJ�޵�R%�d�}��o��@��|[}d����j^�����e��%�����v'��	��a4�e�3�HO�U�GZ?�	�
�ۦ�G��'K$o5��o��fo�s���+�G��z��'U���|�V�Ԗ�8<c$�_z�]��-�} �vs�����Y�iZ��lg�����o�ϗ��������z|6���/9��{��h��b��,�C�<ņ��=W��,y�I<ȉq�x��Ղ��X��E0[}�L�G+�j�0z�y�sj�FQb��j do���z�к���|Z��#�W���Vs@�UTyq�g��.��j5�qyq*�"��0� ��_��>��a.���k�5ེur{ȓN˕R.I��bh��#������,D�R�9���W�����s}�K `{/�׎Y�yDq�s8۽��Om��Rki_�9%-@�X��ar�l~��%�H�X�Γazw'�*tt.�����@ I�D;%Ƿ���i��J׋q�7�H�]S���H�E�r�&j����b�g:��f8���x���K���_Cc	�P���6��}�d�0�1EC��p���?ͦ�d�D�2+�O�f�	�-�".Oh�x��������ke��HVm-���%�N��%�s��0�g�il����E�@�;��˳fwgC����G�\�[C'lD�$���ߜ��͍-Lm�!�],��덟�����O6-�SX ��N�e��]�{�����gj֔�J�tm��aI��Uj���[,���9���Ej~��/��KIau�C7qg��P��u�n6���*��9Qm�B��QK��:�vypg�W<�_�t�Q���A����E0���7fO�tV�q1 ��J�V��$�_�T�ԟC?Tr��2��\��P��55�e
���Bw�jG9l����4L��m,v�?~�g[:f��HV��Lju�l>���Q|�����l]��ƈu�
^��u��x����q��_JWx8@��#��a��<SV�ĴW�Y.^[[w�2[#Ŧ$z,�|�I�;+�:;B?cK����o�t��&�yEo�?��*ց��� ��6��_���Z�^�e�`�(���lD���Q�2�(�feN\��W���鮴�7��-�w�Z���t�=�C�__�.��h �m(>����k�s� w�'�!m���Zp�Jp�XOfR*��"#8�=������"�/e ,�M1�k��Ъ `\�O��|�[≸`��������L�Z+��ҳ�aN�Z�)�/����ZF�~f����i;�!O�⌇�4'�z���~-ބ�4�a��J&��+�J;[WCL���Ugf+��ɽ�]�:<XO�����������6��/r�Yt�����g[�'7�3f�_��[��c����T >�"N��U�}v��5J�Eh�����;n� �X(��E̩||i"]�c��!�azK�{�{�M<�����>��-H�#�W����P�XK���e�7$�~�N��� �i��&a��*!"=�S8 Ncar6��:|�b)�yV�A5�B���:�u��7%�ܱkq������.�T7҇���O��T�
��=~�V(�V��
	^���ظ]���L�!�/@�q��L1dv�>W��u��o`j�r�f|Cjc�M�3�]�i9�3���D��D�Q��?�v��Jc����P�Dfe���7���[����B�pc%w9�I�z��`�lH7�LzJ�Xz�/��ĸ�U�I�,�z����u&cē����릲��i=�8�+�W��^.��� L�W�V���1�Z�h�M�A3~��ذ�?ˣ���s"�c�j=��D��n�#?�M�šl�N����w�m ����ﴇ�<�L2�Hkh�8&+�4�a������ �ŀ�փ��px�_#���0E�$s^��|��k�Q����X��\+�x8�������rBJ��������3;�$ם��w�gvX�*�ܞU���J9̍��"]d!=�;� uJ���K}S�c�f���86 6�Cb����� z�1�H/�1���L�:�	~ ���@�0���	F�/��n����ry4�e�kN�Y��g��D0�΄s�{G����������������Z)�&���v9}"B��p`��g�bz���m-:`R�p#i(mE� �>>��:}x�Rj��vd!��}� R`͏9�>����ϖ" ���>cBF�
9S~k���hPl/�UsB����5jW��|ѥ|P�b�S�S=3�1%����ZM=�9\>3�*v��P�}��4h@�h�\�8N�=)��\��l�e�F0�k���[3�b��k�ǆG�_I��C��gp:#��ͩV7���O��P2�AUR9:�[���w�v䵪"�W��	������Tk?�t�h�xO�3�X�3�������e� ����潮�ύ�3�ּ��8@ �|;��W0�.�t�ò���bju2���2�6ٽ��:ޏ[^3�4Cd�UI;�T�P2	���9U�tKCG�Q���7��p��ډDٿ/�XG� i|4���_ ��-�UK�O@DΪ�a"����kj}�+�B��.#�ﴒ���kԲs�t]�\�
p�ک�^3~&V�z��VA�X1O蜼q�w�0)k��^�؝`J!��qQ���i�Y)�t�B��Ր'�5�^-�0��e����m�E"\����t�RUOf�iM60؉�/Nǔ�,P�E�9Gh˫�ۂb�a��������õ�2Q��&�w3>c�����TƷ����4���v+d�B#��z��aXi��$T��'����7��W^JQ��i]�(�")����{�Zr�M!�F�z�0֊��ٻ[9[����N�*i��iV^��׌#C ��w�}`%TF+\�(9�vJ�F�)"}�RX�9�y.�^��N̤��Cf�U�KÙ+�b�`���k~i	�%6�����{UNI��1 �����6V.(ag}@r��Vj���+Þw��������[�F#���(���(�=���&� .�|H1�Қ�:W�bs����|�]|ki�6 M�yN3ۢ���_-�%���k��X�f�+@aZU����Ç�:7�j,d�x���m���ݿ�/��h�@ꅛ��*��F�^ҕHr�u�<Nԓ��-[Fm�
˦B>���Ma�"4)�J������}�_n��)�MUA�ۮ)R��x{U�k�f)B�f�Yߊ���� g�G�.���ke�I�D�a�)n(�r/b�֊�����ы��U̽'`��꼺<x�n�B�Ֆ�#�J��'� hS�JEv]b��_��i֫mh�#�D�t�<�f$�S&� h?�(�[ӣ]|n6"���m�#0[�מ���CĤvu������s�eS�.m
�ޔ�Bx�S�دV*�kT��J�|e�J@�a�Le&sРibE��CƧ�Qa�V����u&Q�Â���m%j?<�O̎7׻򈢒�ȩeC;C��h��ts�M�P�>��?h��QLĹ��6��$[�6��#)�W����lF�,ͪ<KIM�2l����[�qani{�
�E��2ѤP d� ;>¾�����4�C�T�-뙱oS]��τl�w!��c�G*�d�9F�u��.]�&هs�i�៫�An���6+���=�;�h?�I� j��:��ؗ���|�r��i�ne)�	A�7I��7>���8��tD�NS�z���;��={zC��A/�q�Z?B����Ш�P$����@|�a�Q"���s�Y�/���OQ�W��t՚j��tO<�އP1YqPnz�[���h�?�L[�'���y"�`�����
Ǿi��AA��ny_�:4[e�X��=�$�J������R�W$�
`fu��9���&���e���L#��6-!�X-��Ǩi��8�!�ᦉ�Ucֻ��Yi�s82�u���BM�hwih)ۄ���Si�Tk`L�5>f����=�BP�e;N�	��~gY�Ca���<�ˀ���;���a������ �|n�tr3d@uR�(ŗ���H�:�]ůE�B�ǚX/����U�Y���H�(���!��M�<TN�&����+�O�I�˽�\$�< ��p���e�|4��ϝ���������#+��t�]R�Z��荲�����D�� ��k����{S�4�����}L��M����YD�G��D�/�c����������Ӛ�����Y��m�`a�1l�4FH'6�
�"��@��B�bBޥPV_��Tr�Αy8x?Ydj�|)��>'�1�����+�W_r�fK���>�j=�A`�I搙fV=	綳-�Ҟ=��X?��p#�{,#��K��gK!��!�3�7i��\~��]� �P�C��$���Jn�)$3���jy>���a��,2Tʴ�,h&�}��ϱl�q$��uq��ws7��y(��?`yܷ5!W>&� �@%�(�eRXQ{��Ζ�V��d`�=��I�B��Aߖ�S�]�������@c�?�3"nc�R�eܱ���P�{ז`RKbW��k�!�ӛ#��5Ҧ�h�y2��ڑ�#LU@��.ɲTH64���b����H�� ��Ù��49��:z��biVD���X�{+|dV�BNJ�k|r
��l��r�@g�����)BЙ�D~�Hd3�E1�.H 1u+�k�3k���;O8���������ݫCY���L�RO.���B*Y��e�<����N�U�
Q.�)�7��Ŝ�2|��ȬĞx^���l�5�#]2��5���>�@p��J��n.�
�2CWF�����
�zJ�ktT����9����S�̅��Ơ�7�����`��$���m2����TLW݆�Hbu	 DԷ�@п���Hm��)��X��I�3�W���v�V������~ 5m��~хa��s�˓7:�Q'��i��0T[�<��EP�L��?A�2f�?G���Q��>�b��RK{�.(��Ͳ58�7Zk	��|�Urd=D���~\�D����AR�q:�\��S�o+�����Z�.�&�@9�K�[�B�#f�C�O�%l3��FN�w(��Lo��ڕwBeo%@B�<VQm}�}������rO�l��^.b�D��Н1�8��{��gK@�O�׫�{k��jY�8u�^�S�5��Qhz	|����%O��N���emDr���|_�f_,�10"F��F�يB��Tb�m� 2�ተ�u3��t��|��p�
7���S(^sB�h1�3��B�G�{{��r�'�T\�B) ͚k�U21��WM�d��s�ѿAQ9?Y�ɜ�^ީI�S�,5�j�`��m��-�L�H�e�O���Fl*��î�;��G���F����_�b@i�%=���(���Ӫ�`I���ri"�jc��Y���.y/D�:�ɭ���R;�e�θ���g�o���ntMF�C���l��	�N��c@OA��3Qe�5���sv~}��nz�<mv]��u�-J�	?�0,��?u���d�al���ܛ�(��A�V*�����x��z��mjH���T۝�}�����I?	F>�Ϩ��#@��)#~��"��L:C�~wm����P��:�M��1��A p"'�op�(�O�y����Jr�u��B�x�*�E�(�NJ�A`gr���k�JcI�1��� ��VLP����^f �.����G��tl���xZ��b/�}��t[�kU��_3�t��n%��Ϊ:o��]�Z���L��R��j53e��gw�7 �ǃb���M�L�1�`��n�Dp݇vѾ�&G|�&w�7�b���'�
����.���s�����r���OQ�7�<��y��1��ڶ�����,� �-+�+cV{z:%̲Yxح�h��Y�f��j������j�Ǘ�}�~-6��~� ���Г"���d�<{,ȝ�cmc�;@)q�}v&��H4�>��M\"Æ:�Uz`z02�^yu�k��b����-�#A���Q��qGX�f=#o'�E,���!l.$��\��~fV�ػ�c�Ny]�o=�׾���v��s�&�a�T���H=I�|D;`7�H�h�0��FX�k]�{O�O2sP�[=��λ��Z3t����a�20f�f_-7C�q�K�% !�֗l��h�9>�Dns�v����z��`u�Hp�nX��%~���[Z�y�X�%(�^�=�uC��c�^���h>c$>%Y�?L��KW"zV�~c@Q�ԡ?��z��ur������� G!��U�Ʒ�G���%F�7�xN�1w����X1�כ8&�R�/������J! ��,�R�`�8�},&�8HXU��b5d��SSo���^�XNmM����	:ъ)��b���������O��
H�����'�%Й��'1� q=���2��L����Aҝ��촀������n����� ���:�D㣮EF֠�C��
�x�B�D�_�\Q�og7|R��q�"��#?��0�A [��j���eՔ;2��<g�z%�;�C2�'wТ�O�L�zZ�F\�B���l}��oXnz�T�趻�1!��g���&7�8&+�@.8���WA�� ��6O�Ԣ㰌��L�H'Y;H�aO7�LK'l=j'�ē��Q' n����(bf�;Aƃ{	�`H�b	�2+7-�.�K{c<ۆ�Qq��ư��Q��P�����c��wh�'����pڥj��!�2�n!�i.�r���xѲX�f�8 s�6_O��E��|����ΈQڴ�xA`bB1���������3�Xy�n�@���us�wo��t)�!xC�l��M,�ܞ
#ըV��@4E-#�>*�� �Ƅ9s�q�[� ��^�|�Ҋ*�e�SAn�6����2�P�m�)x���!M#�n������@�&�*:����7?π��z�.�R�%3��ne�?Ol�u�1���	��� ݤV"�i�{�&jcEʻ���ȿ�w�E��S��Y֤нQ=��If^�AH�&DG ���4ҼX��-ic%тqx^ū� �'L#}���ȅ��ڧ���#d�k�S&!�yZ��[�
�����6O��I��5��S��1e���\�[�Al}A)_r�L竑%n���~0!��W����0pI���(�pe�Mޣ��"ib;�xCG�ൖ� ��X�aA���ۼ��o��lT$,w?Qh�	�TJ�:�7�]�� $��G��L�}VĘ�/[��&�4���*(�цd1g	�tr�,�v�C�l���MK���y+90��8�8jax���!���r�+�o�	��x~�����E/��U�Jn�˝ҹ>��h�*w�A�e4����]Ľ�h��['3i��k4�q!�����%耨e�\*x/VO��R�Ԭm�S�m��3��༗��f4ɢ���=���ϩ�P�4o6�t$K�-5?���O�~�E<!c��dP�B��Z�B=ܬ]�H��%���X+L>C+l2��`�2HO<��'0;{�2�D�NW�G����~R���TA��I;S��}v�?�)��=�'_�i�2^�yhå.1]㡴��j1���*�3T����������qܑMt�qj�0���y�}���(e�M�s�y`9�n8V�@}�w�7f�ś.1�L	�������`�e�yg�ݢe�o+��0��t��&f��/-3��ӿT��K�N�|�R�����|�7-��ɂ�}j��/���b��%P�?r*>5���3�i
���܁��^�"���d �H�:+�����T�}�����*���]}�v	�y��W6J�$�-�G$h�kDv��u`��1��ے���fJ�1��Vi���C��������q�H�elq?��t7��3h�Pa���Y#c7�=p����+�5�k)�{�%�I��.xo�R��n+����]��{��Y?�+�w�- �U��tk��Ǟżb����`h�-�&^��Չ�e�I^>CƯ;��yS�5{��OR�rŉb/
S�柳��V�����h��e\[�����X!��I_v��ҹZԩ�T��G��g�?���4x�_~hO�v��}j�����;�:�ze���2�~!o+%\-�b7�����|��H�<�N�y�k
YK�kpHn~�]��a���q�U�r���^�z�:0R#9����z6�5/��7"w�-Ȉ]���C��T�>�+.��r$��H��g�5�~�.�֬#*��e�%�󫳣��n��@:Fr�K�@�d�6\Oq�i���8���:��L����Ў��yV�p'��wST�����+Dam�:���sjg/3��Q�X`��+����5#1{$�"���#皧JՆ�Dnh��@ˏ�̯�JOÞ��=���Ok&�+�G휋�`i�
�IE��A�(���ѫ�2�=	��t��̚4��d.qն$[P���Q����$Y}�yQP�n�z�ew��$i��a�~W�Ö�<��/Q����&qg����Y�
}Y��r��A��X��괗�L5��g=�-Z���?R����ǅmw��Ĥ��8�j��� �.FɈ��i��W���J�Q�Y#y4�M~�_z�w��SA��=�����8,�E^�Q��麥��Xa�3�͗�4N�� ��b���7�ڝ�%��Ǜ��p�޾�����&\lo`Ss5����O�F7��a9/�J�S�0e��*-�oحF��7�~%�������C�� �p��l;��b2�@��;�X��K����A	����;�FU��ֿ��*%�eZq*�pUF�!��]�i�[y����Gva��.�&?�d3�A^��kU��(��ͩ(�a�7JU�J�FI�&*�t;Z��0=4�x��<��f#آl��kR���
�#˞�;����,6��i������b�-,��1��i�����+��|J�,{��R��Q;�O��lC�#{�C����u9��)T0<��U4�wV����w�m�a�vIF�m;H���d2u팶�`7}R��D��z/h�%쇬�23LO!
=":��{YP�1>5c�Ի�5A.Eê3gY���8�ҡ��a��J���!\��Ж-:�2�4|�(�7C�c�v�+fQ�O�mZ��y*Y��T��t�=���a��Q�^�Fq,�=i�Ғ�I�O߈���[��n�{��,lr�wC�������@0\_A܄�E6U����m�9��)9~Ʉ�	�Qy���yz�.���>�;�m(���XV�-�C��UI�1&�;��j2U�4힑G'1�D�`,��a�/>I��VSQ�lk-s)�#��.�΄�p��)�-�kya"�g��!U^j�}��ן,�F1�]8��)��䀫=���۬ �6Zv�*E����Xj#���Z��tZ*I{#�htAlZ�Rڐ�)�����7ZZN���$�ɰ�V˼r��Kk���Q���,�mc�����^ns��D]�dU#x	�{n�t����	�g3Q=�O���7[O�l�,�~J8�Z��>Ḯ0(Ԋ�hxC���U(�tp���Jy�-�E�3R���F�Q�ǶL�V��Ԅ�y��:6��Ζ��5C&PU�-l!�����d�?��aj��Y��j�(¶8����@���U�� ����H�dhk)$A&����n�0bd�!�����������{�%3@���B��B�>��7M����ę&P5��J҈&��H�����TN|�X���t$~R�H ��EY3��L�[D�=\&�8���5-�P���NEe$>[g�^9{ڮ�ػ��c0gb�c��%`h/?��,�V<��9�ҁ���j�a�7?�y� PM�Uu�0����f$)x�	t�4'��C�i`^���aՉx�|G=���8��MQ�U��	�,�֐�$�[5�bqnw�j)D9�*��Qa�l�`X�?Pn�[�de�Ua9YGt���uHE��4qMґ�l�Gr1��.��=*���q�����o!��x:����_�f�#F<���wSBS�?۫�����d�`@:��p��q5��Q�K�CW6�G/(���;���D��5U��8����_TC!>�B���詟̺Ǟ�S���U�C��#-�`%e;Q����H�b����z`u4y�y���cU&�Awēr�&ݍCK�ۣ�K����2D�%2�\�<W���JH�|v5j��3Ѽ��?6̈����L&|��IS�x��d%!ޫH�W�3��z3�R�Xԕ,�d��{��8�]kJn~\.6#�q߬���c�b����u�~� �T(>��Ю� �|�^)��~O`5��t
$��n���{��GR�bК�%]ն���%���Ht���DaO����%�	�*AA%ob��)2O����[q��k(:Tm���_�}Eg�-�[�|�� ��`�����S��)�U��,�ۿL <Z���j��n��c���J�k�ZI*�(���9`'��g��4�C�ހ�����2y'��.�So'�B"���ο�{G��fQ�^ێ,�X��N��sQ�Uud'�;ty�d)|/�j��k�!3眪n)���C��1 r�srX+�E4���k�MqŨ\+��L�|��=P}[)�����dSZ���Ǖ�҄�;���œ�?2f�n]�e��~���~�Ôj�7���%�M�P[��GLXc�;R��fH8BuLRF��M�S�\�$�δ��t��VDC�$�k^�;6(֯�D)4�L��5��*�	��Ͳ��L'p�q�y}y\r��<&��(S5�jƇ��.H�E��%� S�u��6~('񋠞F�=����Zң��JF���ّ��ȂL�l�;{
�&�^�n��'=��qx�%���Y�$0�ڷ�[~�ł�<p+}Җ;�pv�>
F��1����'*Sz��jl�KW��)F%�{��� �{��9=<ώw�O�Ԝ517�B�,���A=ȗ@%�P�@[;�y)t��fZ�u���Ļs�=+Zp`{ f�`�;�©�v,���	���t��@�^���������Y���G����D�i~R��i��@�j��E8��)WaNs��`�"����22��Sn�����Y�R�9QӬ,�?��2��{��!a�����cA.8���$n!(��-7�Nސ�7P?%YQ}��4���ʂ�OJѯ��d�.�������h���F�i�\�Xa	#��=b�JЖ~���g�J�����<u�	-P�Ri��x���ӒM�(?�ϣm0�rpq6(�oO��Z��*���� ���{�(���0�"�����t;H�l5ΏNGY9����Z��v��@�1g*E4�h�$_���
�ܻ������MV��0i+�x�f	-<w��|�RǄ�~z.
-d"�U�A�[�����G����ŷ�##�Ӫ��Mv����r���8�4��3��Ҩ�d�'�
ﳦ�W��(RD�qc$��$��� ���� �"!�(ߦf�蟵���A�P{�2�DS1z�e���D�S��\ g{�jZ��l��k>��n��+����#:��/C;��|����qQ�r������Ov���vxm�D5]��t��(��񺵂���5�_���u�����g$�G~�oפ�_�������w��'C�$���h��Xy�5�%� aa���:���0A�k)��;��QY�����T�/�W��7����G����G������:�>L�]�9���m�ʫ�T#|�q��ػ�5����L��5��ՈlL}�4�M䟑wZI��i��Q¿�":#Rϱ�7l�2�}��El�áдr�$��x.��D�Q�	���S���lejD�A5C���&�/Y�Fx�S�JH/�X�.�av-�P�ַ����b	[�C�o��pJ���}�٢�s]#3Aڋ�1.��	��\n,�Q���]���g)J0X��A��P��wJ:�e$u��a�n|�=I��p�6��B;1�#o8���UALud)���#m�SQ;0�?
M��)�� �d���-^��s�e�E@M �_�H7^�����	p�ϑ��2�
#j?}`���5:� ������;7p����I�^i(U2�:EJH��b©n�6���|��ӵ��`:g~:hf�]�Yo7��2�s4����4L�N�e% Ӏ]z�D��T�{;8ݝ��|'%*�^i����ne}h��۹��-u����r��JO�|����2X�����DVK����
�v��(l^�=���Tz���?�?Z�./7���wq����H���Ь�@����$�p�%�Cf_��S��&�F���۶��=��@鑟�%�t
���s�Sea_/T?ޚ�-$�[��1\-Q�#��T��<��GQZ��V�o�r���z�3��wb��A�ri���K�W�
�~�8��$hw}���r]�L�O���7�|���1Q@ű�|\?#��Sn4��fs�T$�ջ��q���Xg�>��122����}�����WE����Gks�v�wS�'V�:�ݑ�� :���l8=V��Df���=��؊i,4�ē-	lX�=���m��§����|�[�r|��]/1:u�F��U��O�c�.nn�8��e���i����
a���B�l�E����QQ���m��w����=�-�����/�hK��L��U�}�Ҩp��fb��48E߱�^���Րf���^�����~��, �Өc o�	�mB���Sѕa7k������U�G��]�r-p��|q#���6�0����Ċ��/�C�@k�ħ|-�ײ����d?0w�Z��+��jU�4ԍ��'}��i_�+��M�ڮ�J���ڌe�K\^0��z�eP���@�n�:�=/ut�(�]�H{�>�Y���w������/1��-_��� �f�+�P]��rasHф�E8��#v�w9�~מh���<�2������+"����Kh1nc.�3��i��;��aq�67�|�8� q�qQ��79}�ِF*����%�'�U|���1�E�0��i�|b &�3uA��e��_��#9�n����홢 ��3L����5j�����	�g+L�F ��`^z�+���<�}T��pt=�`�m[�ťI�^%��Xa��W�����c��ӳ� Y�/��I��E�(|�k�Jt���0�>)�.���O��ei�$r�A�+�+9ۉr_�_uU������J��^((IT���W�S6ݙV� �j�=�0��W���R7�� �8q�?�5��e/��k��/^�pHu5m�?s��$M�g�<p�|�/$���w^������C,Q4�-�r�d���������>���ԙ��aa̶|��qifBҸ���������A�B��g�w%��9����� AFB�r_�ߺ�X5I9+�WM�_����4�wsA�81������T�˚�c��Ƒa�L�	����8
�|�6�%:��S��U\`	����z�1���h�|O������3�2#��,}W/�C��_b��$f�7�(�	g�������y�u�`���M�e|<_��5��Kj���=��f����ɬ|q�5zV��N��V�����z\���6n ԁ������%�d�Ь��<֡K��i%�%�*�#��9��8��x�u�n��5�EU�֨(�S�'f�E��D�U��U��TK:)���B�|sx6�y�>�7�2k�F-��[`����+���*:(���,�.f0^���N����77UR4����N@Y�ꥣ���nJ�C\�!�7c+x9�o�  ��)n�`�,�kW0e8�h��؄�y!�G�p1���I�Xm��Ů݆��<C�oy��$�^j,h0�tC���M5v˫�~�2��9��l��E�[K������(�=뻺�q�/�D��S�$��üm�o�jЌ-o:y�	1G:��L�X���&��rk�PI���8ր)�h��9ch;�{����9�>�t��CQr���_;��<+Y��W�	����uf�5r}��Tu�E��� �˜&D.3O��vr�k��<X+g�UzNU�І��`�cQ�fy]*��xͷ;;Y�e��(����$��2L����nlH��5���)ۥ񥎖�\T�<cG�������M܏e��"/?s�pJ49C��o� W.�����}m���FĞB��0��<�^�]��l%x��	�H�Ky.s��Q���~;ظ�ʍ&�u�y���\�Ȼ�D\p��ݧ��:#8�u����(t���u�3��ʤ̂އ!
V;��m���Ռ���!�7��(?�*��:V�ɯ��깏:]��LG���u���ɼ����x��J��!��$O�=�43��S.����D�Ff�L@
��.��M��O5y�^~?�>G��A���¿���؋�c��Rdva�vL���^���G=&30���[�VYd
�PO�~
H0sk��w�)ِ�g>P�;�mIBX[�Z�g���e�Z��s�2�b��}�5��hG"1r`�Sx�oi:�lp̜##���0T�{��N$V���Ѝ��|zp����8�
H��HPY�ל ���ܫj]�l~g>��~5�Y�=d�{0�3�<F���n|e�~l�& �a��a�tw���|�����uJ$�J*��ZCg��9G�����h�i;fv�<��/�ц���#^��П�A���Z��6����F�E��Q�zH֠���07���U�|��d�^�ƆJ`]���NG����1?�-63�H���	R���f��
>8�$Gȥt�/���궿;�w�r�{��1O�UjKv<5�q��وz��m`�4YS��1��S��qv�^�V�?P�.]֙���gcʚ�\b���t�ڊ���H�1Ȳ��=0u�6A�̌%�{]O����\����GQ�ٺO�;���$x�̐f��yk���s8;S%��Pi��#xҵp���7	����:LB&	���]��A39�U�@���eّ���"��nD�f��c��3��_Ew�-��f�Q��nra4;��b<�DO��EB��T,ӏ�B�����f�`�Z*����{㴮�!e��xgB}�b�f) I�ݧ�)[��hI����>줭�* /�EQ�Qm`���Q����Q=� A�o���.�G���
�UM�+�w�-n߹Վ�]���=�D�҇2L�:���w)eT�ڐ����U��U[�'\�Y7���18I)�����Emj��ZR��9	��
�B��o�'j�&1�� Ӌ�,0q�!�v��*���qE����U[K�᾿7�k����\�׮�J����<�9`M����BL�)��ԝ��YYJ��kJ���,��*F1�$�5��͕)N���=U�3P{E``��H�X�9r�N��~oُ���߷�8�A�܁"2q�{��A�ݳ�/�SF��k� �Q�w�"In(ދ�*C�6�n�DA��N��d����=�2�M}��u\��׽g��+�~SE0k�5�ò�p�ѤJsi iB�e	r���r�&Ĳ��1�j��R�M~��Xִ�ݟ�ri�yȭG�Q~��}!	�'�ι��y�H���X8i~��&L�T�n;��f�&�Hп�Q���r�+r�"n;�4ߚ�����o�׬�8;�WI�t���؄|ol(c�Λ�:A��䯹���y_x��{���?	"ҡ��x3J&�-��ЪB��ಗ��l��;Y�n�tӪ�s��Eڠq��	����h�B�Y�2�ܤ��#yy��PX��ܞ)���,C�FPY�mA4�[1���ˣ���s&Ks�Z�o�1�e�:־q�Fŧ�48l���j^�F��ő];d?)�H�2��1���j�J������U� �I��sS�˚�M�j�S\c��
x���o	\�n\���/a��Gj�3��P����8����(gƖҼ��X%ŕ7�D�S!��2�U���ܥlS��D����H[����`
���oB�$�y�C��*���_Tе�Hj`�.�_0kF�#B)+ʹMVv� 3ZjyC�������?�4���{�q�@)��\�E�C���A3%4��3|`"� t=43W���u!6F�vv�S	�_�;�b`�8������[����5`����d��_�p,�N��;���N�l��"���0�x�F����\��/���F� {��k�ʵj���a�)���'f�Z�Yc�w�Mq@�]F�>��@�ץ���=��v?�;F�e|�z��KpfY~��f�xN�o4� �������9v�.L�@����TR��:�.U��� �����=U�u�)�)	8��&f�?��P�<��ʾlR�H��g|��QY'�Șb�7��d���-9��7% �+]��@���^�&��B/Йs`{�V�-+�c���?LWV��ȻY�b�*3E�r6ٵZ��;
VՀ��_2��= @tQl�@9�'2J;����G�<�a�@1�̵=�Y�]^FL.Q�b�:#R����2��B�{5q�^�E4@i��2�\��/}'}<��^�6�R,���E�紦�a_e���p)��3Ю�I珽��R:P����b�·�u�:q��X�>d�bU�5`H���;���khSb��E{:l��1�B�^oY9oB�rr�,�j��l����F�Z3K"�z�ߢkq��
'~˭��y����/��9(���d�}Gn����L�C4�7V\r^j��"ʠ��vh�	'�/�"IP%�%��Q���d^��l��㙹a�l0�Y9�,�ģ�$��MP�e���8ImcM��C��| 4L?Lw��Z�Y�+p��]��}�;$*�Dl|�z��������?�5n�0)L2r�b�f3�o g�%	�I��N�h��B#)Z��H�v��HI	:E��i�lȲ��3�Q-pȃA��](�-��|D}3���!�P楁�"}�dx�k)%u��|���9�SǤ�v����s�;?VB+��ʥ��YC���݃X&����F��qypͶ�+*��R�����:-rB�-P��kw�tk&�B���G��u5�lH�X50���<��cط)5v2����c�O��f�Yw������B�2�EQԌwR�Z�\��S�Hh��S�΍B�!;�ּx��S�4�̰����@(����:��H�3��o8�ž��:XJ^>�yk����(�d9�,�KU�s ��$z,�:NƝQZ�3��d���{��Qe�|�Q���x�M�
!��`;���>��?7TÀ�6��D�@>x� }��{��h��Zơ}gC�t��z�f4� ��w�)xhRc~-LWى*v�����^7Y��u��U&����JP�I'u�g����suȷ�,tɢ���Pc�a9�N�Z)�R$�Q7����.�E���&�ԗW�B ��'�?F���;:��K/~��3���!�&�?�S}s����$�+�-c`��FV�)<��zF�i<+7�<�A��3Ή��p�H��ܚ�v���d��ƊC���k	�|�fScڞ�
�~v}���9�Y�q�+X(@RP����p�(+.�F���!���lE��Os�_�?�7A��z>̲5�l�v��8�?滅]�Y�;O#7��J��?#>��8+"���,�*h�?dejt(9m����7,{��ιs��me��/���U����� cO�d++�XP�b������9�k Ѝ'�&J�{=g�ecT�/��t$1��:��7��s	ݹ66���k��j�+� �ё���`G�"Z��/�8FU4S�F�Z.+��װ�������h�_㨿�˽��ᢥ�y���MJ\�2┕�$옃���Ҳ��]���s&c��JI����5����5@8)���N�Hw��~Cx�ͮ�� �F{uj?�	�|������Fr㇮�q��xr�}������I��<`߅�B$	���ط�U!�A�u%X���6��R�"t����������5b(y+�����q�-L��/S9th�vW���1���mPC��,f���|��@�<����x�, ��ɓ�#����'�5-�]����g(�c���׎-D�E���O�^:+'x����Eeq���}`D6W/�(�x��z����<XP�҆�W`�:�;-a���G�� K�G��چ���R�������<��B󹠉��66:��������9P�ݶp�Q��>Œ+�����n�y���s	|Ƹ�*�M<��	�xeo�y�"#f�A���=%�w���'**Β��A�Q%�e�$�-�o����߈:��gTrv@jz�*�y�w"ډ�%4��"bKU&��	����WU��J.�牒j��}(F��<4�1��U�A�E��x���_�>[����Z��
�|\.߭��t��o��Nx+�~�Po?�aM��y�t��ɯ
���{lY�]��+-���9���Ǎf��B#H�4 K�M�aE��k(�,w"��n���~Ǣ, �UH�-�8+I%$;���_���(�Z�׎���oSӹ�#�:-�h������R�b�g#�:�L�@DH������Y�8��i�Ci��C���Xرy����j0����Fnk��0Jw.����椦��`_k��Hr᪀�{�V�k�<y�;�}��)'�>��M���~����Σ������D0Z,A�E{�����k�\m1�����m<��Zx�_�v^�=�=ҳ��s���Z}��D�=@D���6�y���YXF�+b_;[�e���bI�|宿�m�@xgdv����Ĥ�̞����5�Z�G���L�M1+~w��Q�Ӹ)�dw�z�}���ӂ/�]��N(�=��m`���@m�2D�)xG�̅�C�/��5z�u�B�/�Q���n��@ ^�q���_�o�@���Ț��L����!Փ��r��mA�K��%�"�Θ �X����a?��V#�:�|a��㽈j��},��*��:$��0�Eo�ʩ���̇�c�	�?a-��2gf=�:�c$��[�f�D/#��ۆ�r�8�{z�,��ޫ��������*�k�N7�ꥋj��
#����!��+�ģ�	;���b�y�r$�D_��{Q��1O�i��+�iy$;5a�tY(�����ו��_i���<���8:��Qd���+�?�m3�^���5���6�t?�$�X�l��)]"�`�!�R�#���Crn�-�0qhcr`K�R	��7�y����N^��i(�f@"�#��{�(�5ڇ�������w �xG�F1ʠ8V�.�Am� Qf��/��	�f{��$�<�[�����QI�b�i7��1S�a��~�����;�g�w�.�q���H��;���J�V�H�)^h�%�߫=�⻥��g�9x�e|E��;���d�ZU�I�y��[�	q+�B"�0���
��o���W���G�s�H���G/�g�y��x<=-	�1���~d���ƨ�q*�xMeg���*wd�x=Rm�3w�Ӛ ʻ��U�JTvh�B���5�3��:�g_|B��<Ide����a����06�bX�Y�	L�.9��DciMs�v~%������pq�ziK(��V�ߘ9��v�V*�v����+,vAD� �!�pף��e0o������1�N����-K<w��j��ĈbN\ʕ���Ѽ@��o`�%��֞�oc�2n�9��r����<W�sW1��)y�ơ�P��)�+�q��}��K�7�)��6s����t�����nfț�u˄ ��Vv^j�]J�:n7짂��qR��H+�)p�yu�Q�[�Y�1���*�[�}Tun�EFc�	"���_b���	�}���0Rh����)�ՄD�i=Յ|]�����<�X�y9�#����޲�S'�x��a��cm��Z���T�	�X,�z�r��jx� �v�t=��t6�	"۵�X�+������zyO�2j��m��I]�=pt\%�6�'qA�NƄw9�A�3��^s|�����"!϶;$�F�Q�����qU� ���z^����G��U���@�7bA.r� �JOЉp����i��f��ִ0+R�������&/0����N�L1M�ث4�,�X$!�/d�	2�GXôD7<hn�?	�U��F�#2N�7��L��k̀Z���iO��ۨ�W=m1�@�Pq�$�M���d�ܔG��U���
4���O[4�U�6f'����kgVT���n)e4\߿�X�V����&@�P oŦ�NUv:i)"�C0���Ah�4\�K��'�*@�� �}�|��s�g,J�S������i��0�g  �$�$/� �Q.]��?�,R/Q���wε1:�Y�^�o���x<Z�Ř�ȃ��02�_�WK��۱�ֺ�@�F�^t].�6B�KW!�'��Wo��rlB��W��|v
�I��Җh��Aj�̓�=8BъMƍ �`q��!>:�0/�&"�/��*���u"�S'��^12:�F��QE���D[��_(�����_�foU��%�f�����p<+ea'eن���e��	�1�	c�!�0Z#!@������ׯ􀋀���Ӌ�g��U�mi�^C�1��=�seK蒸1��%2�w�̗����̂#���p<�,=��V3�"�-&GX��\J�k}�����۴≇OpiNhê̛졂oxq����B�|�o��S�4
������ւ<j�3���iv��;�{ן��^*�%�9�>����S�����]]Ե�p�c@e�ʚ�Սٻ�_�䤊ں��"��M�<5����k6�4�����䛞�Ƙ6E���5�-T�����L��$�P�oqzg�Dy���x.�,\��;f':�H�X~�>�|�ƈe(�*wa<�`8��e����;]L	���C���Ͼ/��c�_x)���p�>iy������w!��{�`L�2�{�q׃urB��u�",����V}��?� ��u2<��3���� �/P��g/d~Oj��0h�
�_�䶵V5R~���Đ4�8p8*�	e�Y�4�ʆ�Lb��w�x� B�w��&��C���c�`<(������ҿ�,$�Q}��s͸�$��1��<Ni�`��p���qw9��ÿ����ߗ�`��EJ17� ut�����j�̎+�`���������_l�`&w���i$�����	�)��f%��"�g�32"%���n��d����y�-�
x����֑�qh��~��#̧���Q�!rD*��=Y� �\e��R	�v�h�;��Ef�<�Iv��&�jp�����hz��>C��f�L�¶�	�֐�A�)e���#�a;Q�C߶���`&쬠"=�d�,u�G;
��^G���p{Ȍ!�P���4y^<������1�x@��/o�;���ȁ`���A�n����m�-�\mv��B�2\ �s	�6g���g�Z���QB�ܰ�Yh�=����0 �oNZ�=_�\ �:�$��������u�W���ķ�3oܾM�o���_%-�(��(mq���u��㨡�0��R
��a���:�	�Dwx����N�c=h&�V) wӍvCm/Tp1.��v�pR���9%�:r��b�.^sL����%��ul&��n��s��!��� ꧹��z��Dy.�j)1]����P;m�Q��������^�l�R���"35��	�*9A�`o��ޢ���|}��5��R��SI��L[�Ҵ@���w6( g-&95u���מr� c����.c}���E���W�{+�IP�F��'@�f����64�eO��I�fɬ>�	 "���˪6�OL�}�i���p���<�������h�2��5ҧ<s�e����RAg�4�2K���"à�q�И1�����O`]���R���v�¥��a��`S����(��m�E4b,�&���re���T3��_7�تB�'���9�Q&���L��nf؀��jI,]�#�Io�O6�K����03���$t_OZ�k��NT�@��AO�����FӮ��V?eT 1���&ɟhUe�{�#���W�2wxfQ�l�\	�
gG�V��^���C��bm�}U��6�&��<h�K��(%�Jt�zl+u���0~R6���Z��ҷ0z�'����
��;!��´��`� g0�g�"s>����T@�����],7؁&��FPTIueN(P��	'�p!��cS]!%nrtʀԛ�1�7�̖�J	 ��/aJ��*��9���,a���(rP�B���J�⮩U� ��W&��5�]e�Ot�=�[��^�@7��JB�D��6�e+z۵ʠϚ���8���*�&o1Y��"XЙ���)C��
�g|(��2U���7�($�r���7ݰE���1�d�ђE$��)�P�Z�Ά~���ǝ�V�mfA�懰���S��_�oJ~��#���S����4��8���}��H��Bt�}]��zN	�:�d`n�^%'�I�Ңr���S3x���O/��b
��D���B6:[�5I*����U~Hb�oM9n��b�Z��:� ��V���*���JBf�//C&E���♺�w�|���#0���I�5}?�8% `�)�즵��� R�9<]�<�ς�E\غk_�M}<������k��@B��G!r�����eԵd+:{�u�x�7�Ʃ�����B����Z3fA���Ւ{�k�)!v߉�z������y�ԩ<s�!r?S?0X�ӣ*���$/�q�+�R�o�׶0�	
Ό�a�+�G���`D>v�X�Q��d�V9��������E�w�]ix���
+D�\�q5��H&��N��؛jaQ�˚
̺����ӜŖ�����G��ҥR�=���F�;<%L�~,ʭ�~��VG�?�m��Hʔ|�	k�3M�hh�������&�>��x��4��k�{]mq��;+�Tj�Y"�����ߚ���}�ݷ�9аkc��8�H��b�w�� 1Z�܍�YH�	-�C�-�g�-.KA,g&�7׹�Bk[v�B�w�3`k��nK��ǒdBbb�����Xroɼ�HG'�?���iI2T��Ÿ_Z��ܮ�u��V"���rP�&b��\m)2�Ղ�م���.����=�A�L�AV���M�:]������,
5���)��Mp*=�d?(
�8��ְ��
�Cd�]b���S7W}�mO��u�	t�K���㛳�8�q�K f���@��n��Fǖ��p���L:U���d�io)O~�/>ꃿr0[��G3�owL8�b���}��أ�c�j\����`�H9��+�S��MYe�^u�^A��Ӈ�a����x��u[�)��FR��ލh�V�:����H�d,�b���|d������!����޴�t�l�hq22��ONEiե�&�E�ǓY����\l��(��iJW�ʰ��h��G��/�������6:��w���%�oH���k{����ɶ ��,�4YaŸ}Ϣ����.��L�xI�͵�0Dc������`p;�!���P�6��C�U�5��)q� C�D,ǖw.�	#=�nzԑ���'0�0&�R���;���P4|:��Cg��n6}̆4��_9`��|��p4RE�o�!��9x���+ �dtcw�}8d3�?�(�,[;�c�_o�M/�H��E?�4�����t.�bhiQ�eJ�+�S�F��l ���*��,��|�1�I��v�w2����sW�S��!�;��?�*�aU<�v�6�h6��.5tݯ&�����7�f��4K����	��yBYn�-�]��ݮ�;�.�}�L�?$'�o�h����. %ƹ�����W{!V
����vN [���j�E�GY���-����k�"f�(!<���{cA�?Ku�Z�0����h$�����?�Uã �� �H��}��p��H��#�P���A���Ms�����7�����
X����pS�x��L�En�.�!���v=��'�q��]�
'K˛*Z�	��[�M�������0d�]�$O�]�Y�b�UK]x�>ʀ���B޽q{y�򫪍�!G��-�JVi��IID��3%�L�f������f:'�G8[��^���}��5#�a���	�Т��a��	�*́�U�7fv��L�d����޲�n�i[�S�p�����?�ù��×Vn}����I��{�aL��x�K	�vp���y�m  ����.G5q��AY��84zRHF��遷��YcIa�>�L���[�bw���^�Z����YM	�#~5�����#�� �7,'��qI:��
*����d��R���p;򛐦Kȗ��Q�R"��g$�r��ڻL�^�{��:���O��)J�:|�9�{UM�=�C9~�H瑃�-ۺO���ә��������e:��VKN,E�`Y�|n�I]���{�ݗ�J��v��
�<�(�`:nbn��X���u����[���8:O��Bv.O ���ҁ:�?�[�B� f3���k��`U�<�Q=����ެ_
�R��S�a�]�c���DBY��,>Ǆ�k�֍�{��Do&�E�FB�x��$f}7��^>��Pq�k�9���?�䍷 �8i��@�%�,
��u�07�H�6�1��Hꯋ	@-H�]Gf�\�CpǞq�^��ל2���k)`�ً_���h� A�0�A�R蟮0%��(�颓ߐ�x��#�S84\�JI��'��B�|�%�d]��+ȵʽ�
)֡����
���C�])j)�;HlL���TA�3���$=cA��Fi/4H��:�mgm!�s$Ϊ)�UT���'E�4�K��&�Q��IL��`���<����AWl�Ȱ+�����=�:s�h�3�b���W{�ٶ �p����w�NsȦ?�dE�,�=
.�LO5�$� q Ĳo���ȹi4�n^�Ig6R���w��l@�R�K���K3����S�G�ᳪ ��.�&E�NZ��o>;�8�~��	�8<�<����jz5�����?��UfL�.��F���s}��]o�wC��ҏ�7�h�l2kpM--�F�����\�/�2�3A��$_���6��n�cj�;1e`�!v���q���������f�+��gB��<�c�}�?͇`�P��9VG�����N����e��E댐z��Rӻ��A~7K��{NlE�t��5���&��o %����n�<�_��"
��@�//�آ�|���OrS���\�Rي���P�Y15�H���Vl-��7Y�/5Px���M���tI�h�c.����� P�%?�w�@o�2�I�S�kj�h,�I�N���Eb���_��C뻁�ڭ@8����16���M�RS��F��n���:�;�d�wP ���4}��P��|75�[��V���Q�Oūd�@~u��������`�,��"��Z������C�� �C?%�R���T��z����K�� ����� D!JG�7���&	�.]�����A�>&}�C|7�(�V� �q�ƿA����m4o���H�z�oC�NK�0hX�|w��0R�/�ԼK���ɩQ��Osxi��N���]��5��%
� 
��������Ã�I(��l�I�_=[��&���jrj��f��HW:�|Оx��2{�͞�A��}Z��k����%2�qw�5F�s�L���=	�1��8e�=\�: U����{�j�kȵ�p��R�]���ۭ����!�x��)_0T��O.9�v�t �f}��%@�x��N��w��)4n���(A g5�ʴR��*��֭J�U��S@7��j���/g+~����w^�����:3��v�1�U�Z_�u����w�������|FV?9x�;Rw_��>X%��k�H�j����}0�����}��l6�,_?���+t��������խ@
����y�RqB��E1�*���d�˼`8�9��
0K����x�N�ƅh��W����ǈ�ƓA���҆e,߼l�������Ku��� IG�X���ߋ?����a���m@��M)P�L��W���;8���Hi�<6��=�9R�e[� �A�Cn�#GX�Oc�Yl�K��3�1�6_G��[��ؾ(�+E�↵楼���Q�m�{G�CH��w�&�:�,k�½�������<�x�ZEIc/��T�$�������C���z\5ߦnW�Ol@r�f�׻{K��l'�*{�:���������L_O��k�熬�&��p�I�����Pe�F�49۔Sƫ2���	���^��Gm$��F������}�Ȅ������+t�.��i�U�}�Λ���aM����7X#x���ѣSB�rq�X�&6����]�Jm����4&P�� /E�4��^ctN �����2����Q��#�����*ÈBp�����L�w.��h���N��q�Ν�$܁�6���W�A��Cݰ\d��y���z>�᮴�;��Y����k�b����'Jv3�&��cߦ��p�dV��\���H+C1,���� �v�D�:2���T��ӇK#O}��]�/�z����$5�c��]�O'�~jAJǹ�6�;���.,D�]��r�M@��r�����%��xə1nwh䢱�w���O���e��w	�8>L��O$YKָXn����y:��I�g�|դ@V�~^��j�ݮ�r�79�b5	��������?�!���I��2�N��M���/���P�ZGl������Y,��
��k9�!8�-ZI��@ c���p;YU��V�E�چ"GO:�����&�*�j���o
X�8�.�\9�JMl����d�%*U4U����Z�&��ɪ;���w��&�����gq�FQ݃U �;�Ӓu Ժ��&�@JHqRJ2�6���k&�Ӿ�NIm�hb3-�JM�1�����9�3.��'�W�B�v�"����ݝ��wJ�j�М���磥a��|❒�-=���%�ҧ��i˕�b����x��E��Np�F����?����'����Zk����	N��."�sЂV`5ڂP\�9S<dpl����LE�b�l�6<�,t2�?�]�\m�7�����FKX�f�\�{I ,�TK��8��O����t.�n@DK|�\�8?i�E��\����lf �ϛN\jө)�����F��xR��{�E�U�����c��!��Q�H�r��>���˲Rd'0���t?��u��v6퇫";���3���=��"�+#f����O�,#��(h�ƟX�Qpf��PV}�W�ƍ��9��Z�d�X�ݐ7s<n&ۅIv��_`#�^v�V!û�������,J��G��eX�Gɖ�l��f�=
h�����mݍ���S���e�xN,�1$�t��a%:\%�aG�,�n��FP���+��Y,8|�mZ\�4E>>f�iyV��AG7f��jə��&���3? vB.r��Eo�_�uֈ�4OJ��"�K}Xl����/���A��ܛ�l��Ă�()�̕t�x�,x�Tʴ����>�hD\f�ᦫxU�,yZ����R+A㺞X^�Ģ�5됙�MEs��?1�8m�L8���U�S�1ddč¾��M�p�3�^ŗiT�?ߕ��8�  �>^E�|q������6*n��_��d�Ecg�b����%h�v�P�Ios��g�͹+6��;�w{-���1�炘� �	��u&�(d!D���.�)\H��#��$���#�j�'�Z_x�=�k���ƃ^�8D��&u��\J�ZVY-\��A��
~C�g�߼1Gb[�<�3\4b-t��#EGI�YbuUKY���p;�v��-Z2��u��8&���m}��C6��M3R ��s� �H�����l	��
���G����'�]/Nr���F.ů��E&p�2�����a!�	���l�u�����Xj��	ZJ�~�F׵F�<t�����V����c�\ݖ��* �L ����M$�1�>LN֤3�`v00�	�ӥW%�*�T�a��� '�zl(�A��.v?^����=������P�\n.1b��?�SO0FT�Pn`�v#~��mHĝe��\��xܧ���ّnU5���>^Q�P�Pc�(j�3y�4��T�[3c^�[�������7��\iP�P����\5�Å��5�/�bӉբ��d[b��g{ĝw6W?H5��>�KufY�К��ׅ��3�Yn�ut����"�Dʹ���J-���O�խYZ��4��Ls^DR�&�Δe�B���M�>/`B�̆얣Y(�Bs��A��u���>���@����zGy�`�9�MjDhcǄ���BZ�	�̴>�2v�6��@��s�F)#!��{C.uF�u4킺V�S}lL��	�^$`�u�/�2�F�)ھ���ݸ)87Kbi�4��'K#J� H�� ��WW'�p^C�\o2����!an�������J`!8���X��<�7�����`�/3�:��>@�p8�-S�L� nC-~%/[�vh���<��r�t1��=�f�&�U�OG|�]6�zZ��n�.����bw�2'�����%���BNJ�Ԣ����/66g��g{k��*�NW'��������G��#$���z� c8:��n�(�
CȔ��&N��%���=/��5��<h&�O�m*�Hv���]+��`v7H2�{Ӹ��zr������e�j=O��Y|����Z>� 23�;�\���Ev�c%i��,o
:<|�om��}D9/��,x���r�vЛ}�\l�o0��`�v��~G��
A���wpO����o��؊ ���k���ʿ���ƀ����(v,��U�m�
]W�N�إ��^pm������R{��R��������&��Z��`L=��	��x�LY9B2|1�r�	]�Z��hao-p\���c�'X��O�h��A�Ș#B�Z��U\a��(�2�)�O;��^F��&�J��v�+�z�#d�!�x�gN�u8�ϛ�~���|�셎�Oj���X���e�L��e�dod���'�ƨR�?|�a�~������䤬>��qM<��I��H�/j,Y���Ǐ�:�p'%�:�I� ��0���-&w���#_��"p�9��,�
[AE�
��/�ӂ���'P1٩n��Ni�"3�Z�B<H��e��q�:
�ģ��U�o��P�j���ԣ~�&
A���th������ځ������Ͼ�O��
������+�!��`����l�.�M�3%,�tc/-A���}$Bfw��Qw��Ǩ=�3F#�{G z��pE��1��%`���$KQl�YZ�m�ړU_�z �>��$��/�͘�Cwn8װ��ҁ�ڑ�R� j7|f�+�B�.���n|Ò�-�V��*�.Grn�)>fb�z0�u)ɶQ�`�jXd���>v:no��eiO+��s eN{�V�m��Gd�&@�B�4é٣�k��_ҫ|9����Wz<�-ؒ�
�����'���f{����� ���֌6 讀��0��H���^b��I�Y�����ޠ���J�|���+�I
�%��Y����cp8I|r��>�n���^��6`a͒/�&j��o����߯��N�l[�D��h��
:Ű�?��v=NI�  0�S�w-��,�[Ӵ(B���݃|��[�[q��A*4�)2(z$����G?���fi4�� i~�u4�`/8���I����t!�S��vWx�����sʨ�I��Y��p�~��5p�^7>����P�C�I��wj��T�i{���u��9!3]	�f`�`P|�iv/�������H��8u��zH��=����"w�]�xV������:�}F�-���ё
�}��d��IlK�E��^�n�	ti2�Sߢ@/�H�Q�X�����-� o�%���mr�=J���+���$qN��8�Z-(�K{���2��C.f�>$��XH/*N�ld-t�d&HI���#!����o���{�(�t�z�|����+67�g�{f�,��D��D5R����)-Rp���{�B�c.1��5	�3^���T�b�C��G�T���#�=t �0�k>��q��Qȣ2ɸ�5���2���Gk\���Jm<��b
π�'�^�A���}0H+��I@N<��_���k�@�/�����{cX�Q&`,#_',�c��.�Y�$��08�/8����3��~SK�$𒷳��A�/KR��[�w�qȴ 3���b<�x�sEH0e�(�i���(�v�Y�܎ڟ��s+�w_�k�D�v=2}���'��1w^ww��R����B��8��nLBBW�Ӡ�XB����<!�TE��.
���5t!�*^���߇<���.:�!3cSdTN�~�$���e�}��T�/i��IU�!}Uw�):��y��?������+�P����(G��AgE�{��iY4��C܍��8f��r�c'M� "����N��f~�� I�����E�FL̶:�  �@/+��y�pc�����c�>i
����Uv�Y�cL��ƪ)��3���H *[\8Ơ����Ic�������؎Y-p���
���r7��͈�� ��R?v�RP7���i�c-g��UK5#���u�^B폖��~�!���f-9%FzL�0II���[�k���|�gsx{� R�N�Ƃ��_��sa��Q^�˴'&����YK�����*2IgH�Ḡ���?�G�X��
1� ��e��9��u3��"����8I���8^N{�=����TF.x$�D��U�� 	�sH������v�1�l��bOL���19�s��N�\�m���E6�����!�Il={fdih���L$؄�$L	oش ��C)����x�b$�qy��1�ۈO�?	6�<ʄ��Isީpȓ�>[ m����������T9� �m��7'm¬�ק&�Vh���*��J��mv6��\�s[�!H����u"Gn���{�u�"��c�a�^m[QD4��S�R3
��h�����t_ok'�y�A=	 ������L��cx	���H�����P1p��9k�q.�i\^ /���p���xN]���JT�U�{�;�rE�X^������r9���fa�βGvc���j�ӻl�w�¿SO%/�A~��]o��a�p���".��\g�c�g��*������ڕ	}����K"1�'�d���[C�畡!���^���f�=��f��:�%���m#9�E��
O]��w�rp���a����E6���lBj+���]A[�����*/<qN����&9�<���hlU-�a��l�F��j<���P��)�:>�֤Ǫ-��Ծ�SC�|L����/#VFh��z"%t��,^�A�����?h��' j�<^`�7����ǆЉ�� ���0toD{���=�㴦�Y�I�����iW\k_��T�T�$����N.�$�H``�@Tҝֶ��uzU^4T�;�W%Z�5}y/�Pݘ
ܒ �o�>�P4+S�?0�9�e؜��3�OPz٬4V�cTyf�Y�p}G�җE�Mn:���뗥"�./��Rp��D3���bλ����� ���UdN`���!om_)��h�)��*��
U�v��Vǲ��C���j�-މtɮ�jAqJgq��&4���/��D�Da��h��dh�͛�:�~����g:�e��v�2=��� ���3���������̿4'!�{0�;`��8���En.52� Y��%i�Z)��
!��^>\��Z����fw�U�H��#%��]Y.V�%r��|��~)��	�#S�z�9j��O�� (z��z��/$n�A��{����6't˨^�lTXA�������������UEU���Pc�z�e��Kl�$f{�%{1��%~��h�O ��`E����Z�C���9����׽��Kp�]R��nB�kpw7�~]鞁��ÿ�0��IV�}�&����C�_[��猚a�6��>�,����M٤L{Կ�sD�$�TPĚ^+�#�c�ym��̆t��rږ�<˾�3�>���W�D���fZ�9'<wD3��)R���b�fh �''�n�c�z�O {bq3�BFb4�2䡼�N����=KZ4����Ur�����tp�8+�.�R;B"/��na�沎�&��8��-7�-4�T5�U��/� }+�eZ5�o��ݗ����_f]}��Eқ���)���*��L�\���x?�3��G���8hqhe'����W��X�k���K��EɠLq�!���ꥐY�������h�:�r!r��9G�o����V�]���16�ߎ�fZtm|m�&�{ ��OW�)V�p�a>��*�^��k�U�[lR�0�AEr�,,������\����%��4ml�s�� �2?R�/���-��~!1rӋ�ׂ�@��2VU� _�{R5W�Fv&�|�m�{N B�&D�?�õ�L�����/���mnk����"��j)C�an��K��<D%T�� ���[jE����������� a�"xN�"0{�X�A��j�0�Z�+co��E�N���5:�f�N�ʅʪ?��G�|�Z 85^A˄�a���/���1�'Z�t�H�h`�����T��&{���XO�k�v�# R��2��Q�P���Ȩg�
%vECݲ����M�Vͩ�����-2V�N뭸�L$�� !U9B�F^������UF�%�k���!4A�l �Ƙ���j�'R~�O�GmL�:��󈞢�FQo�H�͙�{����R�ͬXI��82�4���Df=a�'�3�#&��~��ᩉ��S�,�\�Vd&7��=.�M�ibϥ�Ү@`yk� ���UR(lMm��A~��-�<� '�@�,�~�����0�`Rs�8, ?�C����_'��lp�ЈI��X�2,�6�Bm�ꂙ�?k�����xǴ�	 ���s�!u�%���@9w'ED����'4«pO�Ļ-6�� ։6�Ƕ]7��К�V ?w���Z>d1J����4�#��)�c��w�%w�=�u�v��p�̥(
��zl��!�[(����A���$�s4�Yf�f��w�"�C��%�_�cB�R9�>���=\]8��:�Z:<�u��:6B��V�\��g�V`9��˖��]1ڠ��_����u�Ӏ�>,�E-���m
��fU@}�#��<�T���!�_�޶%����a�S�	�룪�x>O��,
y0�dS���n`��=;*B�f�'���EtO��fu[�]�2�h���^$���@���^��Q6�i���c����W�p�8����UK֗�m�/�e�����W4�o���5  �G+Nk��xT�T6l;a�����:q#;����X�_,.�/�՞q]�9��+���=��	�GaAJJ��dM�;:�f%��>�opEEO`:Ӭ�bfM�����M;�����L�m�R/\Χ6	���ر��Kd��>�-_�H^�*5F}J���MI�
���E�?�Y�*��۪0o�!�(\ ����S�\���e�V$k��nnN���Aï�ad	67|���8���aT��zLq��� ؃��H�H�=4�%�0���&��ZX�z,9ׯD%�Xw�:�y�:�tR���C?��%��貺���w�G�B,i�qU�x�}:�שS�vr��Q������'Z&�E���~*	!�4��ʵk1�XZ�rSR�X%ݹ�AԞ�lKKC!"��Gxܳ��'5���S�ԛp����T�V�f�6�U �Mٴ��D��$1�H��8Ps;+�Y��P�2p����ʽ��:ro�P@}^�\r?��ᑇQ@)F~&�vы�� Z�.n�!�����	*6F*��7ʹ��pc�T{��Z�@gg�U]T��젦ӛ� �14.���)�:
!/}�~/���&g���O	���J��̸̚�� ����ݔ �j.��ty�b/NC�.�k%��s�3d���!B��Wy���j�y���T�R��B?Gg�U��8�G�3����*R���z(2��nE��ئ�4�Y�� "�� ����h�=O)�t�6��,�Sa��@��G���!�U8�B�	_wJ�T=����h�Aw��桧�율�t�����7�s��K�vQ#J�| ��^��-��l6l_+Lj3+
��;0������~��U�3%��G��3�ģ�E��A
qy+&@����� &e֝�EVE��0c���P��@��bUL��qQ�ܽ=}�BAs�O�6�h��0�v���2��!�`��GH�����5>V{'��0�1� ��F& �
�f^�s�2�a��Vڬ�tБ/�5����HX�����s��Q�f���`� qldk)� s>�۽	�Q)a!�A4���s�Hrd�-k(��4�=��6p}a�Gے�uz@N���@v�cI���B4��YHȓ�-}���75�)1%��XT�S�z»����� �R���=\r���ƖMs�VH��R�����ÍNj� na�e��H&!��+`��q��}��� ���9����4m���R��XCE�i4%N.PF�!���?2w*��M�-Da��� �=q�����gZ����茅7n���6�NC1�G��o`��#��!a6��y?,���~��1�8 [�2M�X�m�M�ͭ���>!C�3D�Vg��t���wR�P�&�09D���8�G����o���0wI�M���v:5礘�$߂/�H��l�I��A��$؅p)�=4�a����$�I��*5$�HU$U�ۥ����h��k��>_�l�$��X�.�b������X�]�!�c/�'[�D�pP���7���Ĵh�Z?�}��k��\B���2�ԍXpdN^���0X|��x�qn�����B�x�o=���|UJ�Wy.kI�_A�6��I+PO��oǶ���M=���D�8�Y`���:��YM�	)Í��}�@`b�i4��;�%�"E������������'����Ȃ܅6�4t:>����MK�	�'{嵣�Nz�y�WI>"Q�Ϸy�sˀH����Fy���gIl�0�A:�`����噣x����bpT�,I�����#�V\�5t�q����q��Zݏ0�Ӈ �F?��T�	�ڍw�a��'�QC}.�/�B�䄡^���I<�$���T�F�F�Y�9:-�>��3�Us�|D�f��c�-�w���б����Gz�o%���_��Ȟ
�vva�\�,�6����d�@�Z��D�}.T���F�0MCF_��R�����m� ��/�3ũ2� �"��#CC����N�rVW��Z"���*M��(-a= l�r�"a��5�� �H���O>�M ���-���X��t��^D8���VD��`���)�GG޾�T��q���ks��|�v
�Ʒ4h��+"�q9^V�m��o�g���֫h`�f��?�ܚ�CU��"���ۏ����g\O�"��P=+��o<;�$H�3R��=��$�ne�
H��a�F��%�Eaf�Im1�f9GCď�o^����Ȥ�Sw�����"�]DB��F�����_>�����F�$W��V^��(�/՜��I��K�v����
����LQ�^[h)d��ﳿo��Gf�'�)F��}��}/�Bh��O�Ӗ��눚�2�C� )�9��?qţ�]m���y���=w%��s�����4_7u�N������	�2
j�5�;�&ۡ'�}7	����7�,M��x,�u�++ދ$n�f��0������}-[��ns�ᶸ؉�	邟��5M��6��Gz����O��a
�"
���V��/:���ܪ�!`ZL[yʃk�11K#ﳗ�[9����� X2ibr��xWM��L����S�$]�1tVlfN����gm�OF�h#� ���%�44kj�l,:��z�#7ୄ`O-�df���s����"w�mͳ��bJz���1>�MGq�D�����3֔!����Ȫ��s��7�1��V��(��d� ~�z���4�+=J�|<�݂�}�~ءl��F_[>g�F���"�,#�V��+�3wc	K���K�X�[W	�!�է苪�£Y)�=�4�Ģ{0ҿ��h�w'5B˟��g#.0U,g�W�fZ6`h����^��(Sޗ~<Z��W0!2����i�/�V��Y"Q����/c5���������VĻ[�_s���L0+���*~�U���݌g̨º�,'�\_�H9H�F���o.�\eK�e÷�`H��ۺ�(uT���LݛC��5㩊J�����(��6�~�`��U��o���2�dF�t{!����%��Z�==�\����#V�^̮�МzH���ڍZ:_:(\h������(7:����lN��F�@l���\�N�T��؆Wٵne��ڞ��$Tj?��6_���{v�VҷU�h�@�eh[�I����`oh���������5���}�mt� &�5P^D��R���=�Z2M�(P�Ӎ��TPbWN$^Hݼ�<��+�ړ��R*6��/�)��Y����*y@/7m�(u^�#*��Zw�W4�E�b���Y�N�t9M/G2�̒�0����Ơ{�A4Ui�.�Q�ګ�&|�����d�a���9N�[��c2�s�&�;�겋����a~9Y[L�P�*���J0�w��N�>#ڏi�3z{�=l�t�64O\�L}JvZ}L|��ggf�97��;�ӡ�4)yHP�����i���D�"�k�u��o��|��B�p���B����b:jf���>f`aM�ԟ��)���ђ�̈:<
���Ic7P��vq���R״ʨ9�U��d��tڐ|��I���~�	3��t֙{��m�L�TQ���L� �3��h<�1r�4W�>��6�/5� �+�@p1�U˽D�[ �u���6��8<�#l=;_8���JڲR�d�������6�m���?���q�bj��Hm܇��/��Y