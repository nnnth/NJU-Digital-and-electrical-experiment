��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��ϱE�e��;jމO7������@hF��g�qd�8b�-�wV�q�V�mhd(��`S��`�o���(@�]º,i�S����@��P��o�3���o��yOL�����g���j���l>p�N%�'ʆ4/M�D�z1x="F�V�)BG�,-�*��G��Ʊc���i���hT��� �x)�s��	*Z
��i&W��7R������������E��t�+R��]��rB��,�L����Wa�m5jn����C�������m|�0�\>�u9�I�*��A��.E{� �q�$bB݄T�8a��p����h��j*Ht�d�D=�6�쮶T�A&���JGѩ�b~�?�����DB��=�B�L���!�n��`�v��`�lg�e��>��'����C�?��3.<Jvy�Av%(�W(�0d=�V�J�N���%�ڽ�����l� �Z��h��z��RQ��B Xe� �]��H��%�!�5)����z��9p>���+q�EԟY%���+{WHʵ�Q0���z���em����.���E;t�[ ԇE���h��ǳ'^�@����kՐ�X ��g@�;�[k�o� ��Ⱥ�iE����R]c�6�l�Qar/O��譢y��V�+�̄�|�zl`�8���� 0\�:'��vQ}PwG4b��t'�`*c$����5`��9��G�w}-��X����+:�A1'�ͺ{�^�A�sFD��7ǅU�t�Ώ)\�<ۚ��
�m�+Ю���Z�X���0�o�Q�h��:kc=����8N����� �WD5A��zf��I�a�)�g�"��8�7p�E��:���v&��$.�aK|kJs��l|%�@�=�bE�+&�����a$�-��%��-���HQq�H(��*|#Y��G�B!ebY�@.��g���[|�-i~�-��xDj8�eMb�u�f�ݭ�^��osnM�t��*nm��K�c@S����n�""��v|Lr�<Et\Qy�I��W�	�a`RߋX�P6.�����gGY�O�
V)%Ѹ/�s>��I���ڨ�5
�r��"$1'��X��pF,�T��4�2´��rTX�����+�5�y�RGĐʄr"X*ؿ�(^�⬫$Ϗ3J�GT_����ʼ�����g�� �'�I������6{x&��kG��y���eN�D�aо*�Q��7�5Ps���a��������@�9�WQu�0C���̍����#^�;���Y�߻x��b��3�ݹ���2�t�S��b���3>�8���2)���.i$f�4�z�?h|s� �VW&���1e�̽r�Nm�ˠ��ŵ���tVD/�k��A˖~zO�R�*��vԁL�A~OY���ƪ��fF�����x���W<�����ܰ6�e�"0em�'#j?w�.��A��Q����*��7խ2ö��%��01�R��^����JA䶤�JY�,
���S�����1�ru�;���qBi
�nWVQ�4���W��9Z�0�d��׎y?fo_��,�w��u������c��p�>��<L�lV*[#���$3n 1�}�^jA�c�f�h-Y(��F�ARsRs��N����h��e���(%$�ta�&��<�����U����+�n�THC�T鏅���7뼖1KxN[�PG,|�i���e�⫿Ps�ɶƊ���7>�ѩ��,r��t/ҫ �I�����؁;�U�	��-�w���Z��؄=qn�L��><N;^E�a�4#+T~Mn�@���>���F��D7�R*�UZI|���͈3~�>��'1���gg��1[<֮���9M!���U!.C�!O@�&�6h�h���;�:���o�AǴO?�XJ��%���b�]��;*OF�ԢQ)�Ű�;#�+E����O*��A'��0�n�},=����(��A���]&��� (\=�0����z���)j����Q�.@��"��;٥�n2�9���8`�3��p�E��a�Lܳ`�����Y�3��i�ߖn����\!�_�'ul�`/�:��w�~�yK�ٱ�_���($$<캍5���]�!J�ED��vɧ'��T�_���0fF�qPr}����/�P�'̰�|�B�nDMl�j����&��m���c�n�S��{�}��$7�3}MгZ�����f�M�o/�e�7I���p(+�t4�Af0�������LS���_�5��;��[D`���a�D��FQFI*v�!>�n��p�D�bZӄՄ�B��-_�$A��1w�:��9�F�T�P0C���������N�1���:���_�8GXr#T�[�ڎ׮�5�^�����o�z�[�����i�3�OW�1,<6��)��ȑ��R�����O����oݲ�8Tn�{���OPU9�]�T�`���d���}�͝�U����\��aҤ���Ha{\��|���_<B�.�n��w���&:$�%�u���ك@��?�s%�n�Ǫ	47K0it���	<�a�Z�;Q����H��+�#�����"��m;�E���X��m�x�/2P)0���&�\�����O�`���CB�5F��piF�
O�f�T�^��N�3"Hd���,��f�@�1p<�8Na䐣UhD���RG�G:��<���?��<7�{B`���bk���eEqՎ�a���!\I� ��ަ7���*�ڂ�J���]_���ܖv�3���6X�J����#�5�f6F��?��ߢX��BE�}�� 2���-4��ǲOӧ+`g��_�ӡ�)��P�h��e7�����-������.V�	�$Z��e�	aV<N�>��~8�QM�Y�F��92��2D�(�*�V���Yd�Y�t�Py���r ��eQj���j�yߦ��9r���}$�Ɵh_vA�Y4�T�_O�^R�|�Y(!g +��EE�&8;���WI�x�P���VکA�g��	^���f�l�w��oHҔ__-9�1B)/�� *U�\+�%?�f�:QTZ�4�~�6��t�,z?\�,��'�U+�szP�TI���r�
��s ��S��xE҉K�ї������T�:�K������I-���٪��香���3;�>�O/��d�~��(4���	����,���].E;/;��1��1�`ZE���`�c�wq�w ��LV�z�ҿ�d&����[�~�{NT��dt�A�>� Q���D�K�$�� ���ğ�dlq*�.��-��?@�S�芠��0�(�(���X�v�����G_4�r���J6s�*��YR��]c�9�z�])��J�PQC�w��u	P�f�l:��dݘN�p������Ey�]"`J@c9鵘G� @2������f����u��T�Rx�|6/�t�_0D=;8�R�ը_���~��<��E�2�9r�יD�y�K��%�	�iJ;��p��f�لέnC�~;��Mop�i�8����M�}f��W��+�f�y��뭃�Qn����E����6�����M�	��X	c6<���_"㻹� ��,��jzY�	���R5Ԫ�W�<��[�!���bY&?l|N~o*�'�Q��܎�������J������QnZ7b����Q\2��iY�XO��t�z�)X�ɉ��=���_6��P:+��14�	{��-���bJ���VGI�j���ȷ
��y)����j���:�)�kz��T���!�ETHv r�r���q�#:��UH���u�z��g,�0����:��Z�4M��O����c�R},�e*]�I|� ��k7#l�q��W}K�����ZÅ�U�5NgA�V�]R��.��Z��[�R�{��7�ų���G�����д+N�q�s2����6"� 1[qc�DN�Jv��q�O�MY;�k�%G����j. �Rd�J�(<i&l�@�]w@���s��ʬb��b��+&���͚~���&�:*�����	J��q�*�1�	~����u�C��n�q�"�>���*���h���en���u�>b�f���)' ١�≻�$N�?_��Ҕ���̭�K(KG)u���d;'�k��d�s�~��a�ef�z��Wݩ�.�x�w��4���q:x�#uT#��u���Rd6ٿp/�ՙ�y[ցr�3�VaT����fR(``U�@��$�.�B���G��y"W���7���ѷ8��g�p��x3�&�	�b��_m�R3_������E#�L��+�zwD�K,��x/�,X�$b�p�&�-�����{�!pL��w�k3'�fr��2�f^��`ކ�D 仁	���M4F��a���!n��A���N%��r��1��g�Ra
��JG&������ ������j
f [�$Qq�
1��;���.ϲ��eH���Q�hD�EȰ&{]ٳ��uHfF#3���c�#��=�Uf��͹O�?�%��|Djݮ[���>w��"���s�F	��P]a����}�5X�<6�ǘ7d��z@���ȵP?7��X�Ĉqcl��7�=Q�9Ȅ�2��o�+=��� J�L�`#G�Z��֌�s-��[���љ��kiB���0��Qr���>��9A��.W��U��:��B$	���ks��ad���@Ǐn���nLB�
���!�0.�����ĩK�S���L�ςb<Q)3��rf���H���
��m4���8��Nf��q�Jƴ� ^Hݓ��s$��!1�j�(4�z�~�P��d*x���)�)�{`/Kόo5$.M�Nѕ  ����d��n�#�ùi���W��YA;ѥ�ћO���:�%b�㲪�p[B�ھ�37-�A��F-Y�$<Ǡ�63u@u��/X���!݅��%�'��rj$�����ʂK�j_�MM��q�&A_ ��łn��,؜��+�7�%���L��as�I&�2�{�?ČgXtn?oӟ�ƣ��T\�1V��Xay_�+e}�]@ͥk����+@#�N���ԷC5k� 5��g꒞f�1�,��{ֽ7>�vFa���F%W��1G!�'�Ƙ�N����bJl����H˺���c��c��������᮰����*@�9����G~����>	j�w{�Zg�O�S%Vv*� ;��E��r �#KK����O׸܃n���,tv�BW����h�A~ ^�!L��02�F%�M�5|wܮ
�yN�o&�B�f �2�А�=?)�$���l8f�V�wy4L
�Ñ��'N����"��?2Ca��N�IT ��f*�\����~�B��
(����7��5��͢y��gO�����4N�M[��$�-Bj�����O=&�sxpU��ÒM_Am����<�T��-Ã�_b���[���i $�9b��W�K�,�ݤU�xm!\օ�J%"!=�a��E�+F���Dk�I_g���E�"�o�����ë9QJN�����H$�~H����,듷���D\\T�:�hZ��G�7�Ew�>��ޛ���2��sK��+�t"#�p#�YSh=�l>J07��I\���l���9Fu�����T��lo�;k^Pi����ǈ�����Y�m�\PȀ\�m
YԴIa<y����� ���1���K'��No����.�����;����7�dͣ�ɻ�1�{J�^�h�^ix�t��y$�!�?�k����#�#��eu��4>�?��Ȝ,a΍�P�KI��C�4��aZ�2��������
C�'c�0QŎʹ�떤�w��'���s��o_5u�=yy�z�d�D8�Eꝓ$BfC��>��+h5�X��n�L_��h2Ȕ�m���i��?I@跃�q����~��E�d��'e�q���K�&�ZiF�n�sb��Fl�:�	>�=���C�겟ߵ�\�ɬ��*}�hT�V�o�����`�}���+�5�:sX(]��:+���-��������U����1�9駈h�� �*>z�F�z�v��(��æ�Oz:k�R`.�zL�X{w��51ܫ?҅�vE'�}Mz�q6� 5ϔ��;��B&%4,�� �;�R��rP���Ɋٖ���4%�~E�i�D��`���y/�ꭝ٥�=�r��?����1/P���:�w������"����5
\(�_x]t�s��L��A��M���Y%S�2͆�1��m6����#���Z��E�LĐ�N��ɛ�9�[���H8Ȩ��˜�N��Z���Q�x��U�6�=�|���Z|�R������j)���3�o��6�'4H����&����+�O��8�~�L�n���]W��i�f�M�?�	O�j�a�LF�G_���sxK8�Dڀ{��d~>���Y�m�߈��t�R'��*�Tk������d�E��e�
v��Ӻᕨ�"������2N�BVj�6��޽�.�|jYҺ�o����n)<"J<�(���B|��2 �.%�=�c�Կ,뜌����AF&�j�M�m=Zw�N�,���p�\�"㈪������	�^h�%����"ZR� �@	�9=��	���1�G�W���*�W�'��t<;`���Ó58��A�>�/�N�jw�	VΫ�S���� \S�Ƚ9�������{�	߃Ȍ,\�u��'6
]f[6�)����*��"t����s�|�'bK�*��Ivx��3���ֲ����}h
��Kب g���g�po��VD��Q��8���aI	���^J��`A��,�9:_�/p�L�(����HG�F�.�[EN���ďx]&&~�����]|C����`$�h����K��Y���j����C�WDɹ���ƌ2�L E��c�$],�,�W�p��]K��0������� 4T�K���,����>�ʴ>��eH��˺��b�Ɉ��_O��<}��"�hfs8�,z �$@ع(���S@_K	��qn?r�:J����@W�~�<�C�&ßфQ�Q!C�������.�j�]�1U;+B���ҫ;���*�$��$��%JQ>z���hʵ�RP��!�6=�$�2�\�d�'�!�#���ɮ�J7�����w�_�>�,-��ѿ��!�X?�.ϱ�/�og8'���%K�Q���֯�����"�k�p�7a�8G2}�$��f���T}L ��� ĵ��9�^�6��!�/rӁ��|X��k��L��R鵁���78�чg��.ooQ���ᰁ��~A�F
ѢK`��U�|D5�e�
���U� �I%-���aF���kA!���o��4�7:��H_�օk}�)���q˰�u>/�~�f���f9&����(����B�c�϶Ey������<H �%3:$�����8&c*q,K�О�ɝ#�a���fˤ
�_Y�9{hE\H��?(:|a�wq=�y��<�h��^۾!�o�Yh%�2:N�+�w�$A63�Uܭ��HC��on��%�8�\��N�B�qN_�� ��5�Q�Y����[h�G����?X./���gMp:�.����l��N1%�>�RB�M�"c'�ᢙ���!���eچ��q�U�zQ^�!���/�*oYl+�d��6S�و��.֘U�i�3�%9��{�����+MI�����(�L2]^K����4�"�����g�/o��8�V\�_#�,xڿچf�%@�xPg��,�n�	�~�
�u���>ھ�R�k/��u�q�/^67/?A�7er�\�#7���k�]�8��[��+�)�V��Va��(.�T8
S��Y���� o^��v
I8��"����m9�:�D��L�����:��-�s3�GhΤ�&M����'�M����|�)��P�
r�������b�G�Ö��~�����s�	c��"Me�[�M��s�ϭ|Y�����[*����G U��N�<5�E1�H%��N6����1�¶2�M	~�_�3���7��?k]�S���5q�s ^�V�߲.t�i��S�KLeN�	j'�$��Ci�Au0�円'jׇ�y�k�70�-)\���i�>i�Q�Xt6q��,����[��F=���t�m� �=�GU�i-m �:��vD�7�Q��'��wz9�@�p{Ah�ȡ�iIp�qk63u�������7*��N
�B����`nu��M/����Z�x�N��lH�'����=wp-����J�2���
��1=Jd�-i���=j�3u�!��&(�8�6���4�Iڀ>���Q.xȩ�fʛ��b�����4����yTi�<���0!jztY�'Nj>����P���{��&���Qhk$d��\1��E�G�$�:z��r�����ld,��_m�&0E@�!�p��93�-%t�=7z
��W�erwa�v��d�=���1�8U3�k��s8����Á#F��K�������!b�@�l3��O�.���{��Ӷ�0$���uhG����%14����8ŀ��2iw���%�Wϛ�wL�Уj��"����uJ�D�$��g��F50 xϟ��j5���H���z!�ɿ��I��Z����k6�I�ԭ�����s2IgRl^]���Ɂ��ں��H�� ��x}�us2�����$���H8�ַ���7P�B��6��1����z�nOo�8P@���7�_ݙ�b��o+��u�h�ĿɁ`�kW?��8��Q�Rd��?����X
����#̄�=�q��N���3LJ���c�J�P�$@y��)�b�{4��U�N#Us�����dJ�%���p/���z�L��q�t���l�]��H�FA�G�xZ� Yi��<U�+�AH�q�dl=#6|�L�{L�g�A"F���D��Ts��)�vb��D^�\�W���F~�=�_Ϫ��=o����ܥY�a�R�"���i�-࿡�tz�����s��^箊g����KPW�a:�f��/��O�]� xl������I�v�)�~���ɷ �|�yxF�[N�э*��7����_u���6����������J_Ty�i< j���lg$�
:/��~����ڿ�t��%�*w��!Ɍ{T��w�U$��lr�C� �F�ˢ�1�2�]Z�޶lYℳ�Y�Q�aV/4K�Fs�[[8T�����JZ�~t���_P<���
*X���S�V�,m\%�|��,̜��ri�83	��7^���6��P�W"�:�q��X�3C
�#KQ�|�<�i�����K�>,��;����=mK����6�b>
�UM�A�oh�P�{5��Xf�~���[5!��n�԰Io�>)(rq^���=�X��iT	�T�o���{\���Β��U}��/���q7����ag/�)MJG6�����v890HRj�>B^m�ss�q�	�k��5
i�k������[���g ����#���2������w�b�F��f��<�(�O=L?Qz���̎�Y�2"E�q�Ư|S��J҄J�<ݢE�y8i�2�Ù�R�+B��*�%^��Ԩ0�/�mv曆�a�:~,�I���@�)��k�N$���\�#p� �(7_6�������lC���d���=0*�C<"����A���&�+���Z����%4�\�L��Yږ!Zy�A)��]s��t�<����'�}w������v�I�j���O!;n�5�d'JEܗ�Va�J�(�>�ؙ�v��-�җM����zb0w��Y;�c%b�����B�`��:�*��x(�)k��8�N%�O�r���^��&t��yeTt���y����T��m&� &��q�Y0-6�(�r%i��Gjp�R�1���=t"='��]-�����e3B^���&vjΊ�^��G� �Eg �#�@-��l�X�m��a ��L���B�?l��z82��&9tD�$k�LCC�0�5���2�_ ��3��uF�ϲ:tͫ�㨹vp�#k�ה���Y~C��x��v?7
d_����Ò��C��+��F�D�=�8��?�ț�{Z&9^'o��¬���W�o�W���Asp/��=�>?��F�s
|l# ��s	�A��	����$�bK��~=x����1�
8���* �{U��m;t�����д��td�s�]+��R�D8��eH���Afi\#��=��P��m�l��e�G2�G΋�*���O�_IG��Y`��&^xB�̷�\*�|S��wD����XB��`$+z���'�
���������N����id��-o�:$Ȃɝ�Y���҅B��1��!��Iǐ��J���?,��p<�pߡ:�^8x�6�l���{�Q��O���hh���)u�ßd�P����G��BA�I����y��7g�]�����ܩ2��>��֐�m�&CWVI Z!6������~B(���4oF4@����~�N�?�A<Je���AB�����P��yu�W���d�-Ӑ M
�f��n����m�cf�:�B=�p<�P�꿷��s��_	-��<_�M )hdi�R�P#��^<I�UHX���Z��B�����\���^Es��0^<�����c�)��#̵9��6m���ީ�2J���9�xA�vq��-��t�6z^%@QH����U����Wd�����l�7A4�����5��z��;��S5�lV�3��-��t�����W��s�G�2�m�r:���?�"!���ҩD�!�=�R`���e2�P�q�Fv<qf�R���ֱ�1�o���6��:���Y ��&r34Yʳ��� ��AC<m���ޣ�8,���\{�31b�_~!峴�iTr������+�aJ1�Z���z-%���Q��c/��.Z�t��y����1�t10F�m�S	��2�-�Tb6ӇES�闃�F��#�Ս��4k�`K�@�:DT����3)1t�����X���y�I����p�7O;>ݟ^�$11N�<��u_XWAa *=z/�s�-=�r�Bj\S�fw�?�p�哊{D�Iw_XP��>,JO(� m������'�]�$��@Lj�nhF��*%�C����$ơ�Mp���7������}|��&n�Ɵ�t&:�~Fm�W'Ut̉�Gyk�M�L��EÌ�ˁ��,:6�b���*	����G��]���[��;7N��J�ۋ1��"�OsrR�	���B� �63�zhTE��jeZ���P�!F��Ƴ�.u �`|&�#Q��΂cm!+z��s3+�Z���JU����aWׄ`���1�䯭��8�.a:aՁB܀����� �R���QT
3ҹVڙ�皠:<C�}m�Ώ�9��w��� ��S��k)	YMS�9��n�[xm�"JZ�>������e�o�(�)V-`���B��{OQC4^�ի��� ǂ;��W�;�Hw�'�;��&��5�`-�c닝�����n�{3��meD��dP�&Uv���"<���4ofC�A|k��K�ɭ[�ҽyO�XU�W�>=�nIB�U��`$����OK�7�=�Z$�ɤ��L:L�Y	�n;c`��LS�G�'���i��סeP�0�pL�?����T��ae�F�,�v�s�H��$�yYV����qmY*zD`挳/����/�u�#o�\��X��$X6T#�5i�3��]��xSY��Q��V�x{�M>�Of-�R ���J�4b&o��7�F�*�7f��*f��R��*�g�I���=��ޣ��>�n>s>��ʐ��}�dC����-�y��jF9�p�	��Bg����)A��,��}��RH��r~ h��H�+\n[`�v���|�W
�v��(7�<���:�C��|ƍ�e�c|A���ly���t���ąm��� 6)�:����*<�G��i4-��8mZفV�d���O?�k���(6>�n*�#]�>3�hG���"M�B�"p�>xָT:P���ثjE�����n�o<϶ٲ$VE���X�*_��8ε�4
�'mr�%��� �~^�IGv2��
f���ꢈ���DPDas��;ۨR~��d�f\��+ ŉ����L�![�~���UQƑ��ϑ���=E���;�<
{�e�B�<��m]���M����U����\�@vV�eh�Y�VQN,i���ܪ�Mz1�e���X]��xV�%���/���|�{���kz��m+��_�K��[WS�uf���ER-�@�|R��$�e6ł��oMS��E���6*zݑ��|i�:�*|��u�"�'�Q2� �H������UL,>o�����̎<���S��\u�w���� ���ϽL��kF���`��ٹ`�{�Z�_�[��-�%���"�c |�Oعx��G��'�]��B*�<Jʙ����+���FIW�0�@���c,��.ne��_#�f5���qa�x�7&C��Xb���@V
��*�M����U�$*W��WX
q{�د�È���6c���,��_�Z|��LS�3m@%m�e9��hu��$*�fG���Y��� �	�apU�09rR��W�Njs�[Nu+z���Gy$���"�X¥�C���kv���*����s��I��)c�u�x�`��v����hWh�<��g�^��)-t�A�^��2�ljiq��?�E5ΰ��;�|�a�m��7��kT��U�LxA� �����,�kJ�1ʙm_��������kN}�H�d���x����:^O��%⼿���Gk��6*6?ȡ����K-gmC`W� ��6��a��U��%�f��Q��R�y^&�V	�+�꿢��֛2�6�s~y�����D��K�?����ɇˤfs��(��n��箙�w��"��	5�b�8E���`�;����\�C���T���w?А�/�����Xզ"2���f��p��nd!F$[4�C�p�f0*OL/���\�6�^�fAu^�a��������}���Y)�Q5�MB���� �a]2 �Wq��R͚<~W$s�Ms��n�y$�t�A"�����^l"1��:�A���3m�v�<�{�����!i��{觓F��|��:h��q_�r+��2���ǜ}��DDV���n�G.� �(/hE�w'���g���B�ܮ�&�*seG�H���漢k����D��ʃ-�� ݴ8�0�)΢\m{#�v�J�̷��~���%#=L�x�0��V ����r|ɔx�8�v�w��i��m�A��#�D����S�e��7��ػ^�����	���ǖX6�g�[�C��ű7c�<�:����FV�V>�۠��CYM��,�gE������-�,��̓���o�<Zz'���2�=�-��͵��Æ%��B�r�
��k~��z�I�W�A{W��a"���w��9+����۶�4�@=�� �wv�k�&L,��f�C�kԪ_�G����|����0v�S�L�-�)����b�ަg'��R�I[�b��b��H~����.䍫�	Nl�em�)1l�#�	������i[��Ǽ����9Lz}�����오�^�<j�h�������9T�tx�3Z�S�^'7M4sC��Vz���u�� k$b�+�#0_{
���W�/����9h�
�Kt���s6~�_��4&�݋$���e�G���t�ى�� \g���~_֫�yi.�ӊ�L���'�D�FR��� L�2ճ��f�7����R�{܈�u*~Њ���<yr��H���|�@�E�������n9 6m�͔� �,t�y�����?A�Maƒ6�W�c#�N����(7ք��̧���.��q���{�3'[�uY�x�	������O��+�OjIEp?�����XW	R�j%����Gs��x���gݍ�X^�,��JR�mCGI�T@o�+據�4�J}�̵��VN�o�M��?�k��BiŜ��}'�� �E'p"X&暔IoD*PUFы}��ID�r#��=��s��g�-랂J��h�[�¬� �δ��!^]fqT����G�r܋Z4%�_�٫�,�0!_X�w�H��SH=���K�"�*o��O�V�(�!��+ �ٶ
�h_�Fs�ř�d)h���Mu�Zd� �(�� t��U�io�¿Z
ν� 5:��S�[�3�O�̠~$�ܢ��Җ4s�����}[������_5+��o	4z@F�B�B�[h�Y�P^��k�h�&� ��i�Tg����~>,F(����K2����j,��CY�3O.�+�_�46����q�ʭ'�A�����_��b7�k�I��Q?�E?��.;/^��ʈ��d�N�K�a���4�B'���K6��CE_1 ʤ��ٛ{��߃�d�`�M��B&Bʸ!iKO¤,	Ē��>IjHEk>�yk�q����e-I|���a ɠ\�?����H�sW-S:�F:t�2vIp��'f���g��.�nI�a��y  !@6~s�%X�yk�K�,r(BW�1{���������� �-h%���DFj�?c#Vc-�+���kU� �}�^Ǉ����'}����=Ä������T���5$S�Ώ) ���WNOnura�Zz)KrIˋR��L��~�b~H|\������{�h�r��T��Su	D3����y�����{U zp@NY�8��F[$+L��?!��B;,��n/g�ē��gm�W�M��-�-Vu��)O��4oLl��"^�����D�%��߫�����TXH��p��n��'V����a%b'>�S߰׶���̮,!c|aTG����:�敲t�md_͇�4��_h�u]dھ�c�զ�/2T[��?��2@����[���?G*H�D~�For�kNw	�A;'��������r6P8�Т�\0���4{����5fG��=��_vE'�ʽ+�M������d�GKN�Zy��C�&��j�f��|Dʥ��W����ٲ=� �.|�r�Q�F���k/�X�8�Vg��6�y�� c;k/
��̉>�,�(�~3�^ݝ�������Z�TP�l {���r�ο?���q��Y���[5�Lp%�N��1�O�4����M1����90 I+3�az1�p��eCS=�I�=@��GǗK	�,��5K�!IÞ#����v-k4��!N�҂�\�{��<Gܤ��kz�x��oG�d����֝����b�dv^��'oX+�P�^[5�s�o8[����]���Wɓ(D�|�I`�l��~�$N<�d�%�T{O�S����.6p���{��������2$!�_�2�Z&Hs���u�]/���۫g�=��GGa�l.�ɖb����4�߹�P��a�S�LM
ȵ�}����R'�l�Tޥ��e�f�#'�z��e"t�+59��	�fA�����b��u�''�a���]tPdپ�z0R��4k�����7�;��y�T�F��ɬ[J��[4�>���$����sQi6�a��VZ�=��XǺS��>��_��6���8{��nB��ހ�jbxb@+�� �.�ԿY�N7�����o 4QTC�=�*��%rH㔹��T|��e��~��@9��H�J���2�d���~�䁟��	�ƌ�:��"C����6!;��9`�^�?�x��r@�0�B?�ĩE�w3,�G�/{b�$�@����N����G`^E}�?�]O����'l'E��HȰ(��o�X�v�>Ee���e��ۥ��������uV el㌊��5�k�Iml��2�q����KX�{^� ���n\=y�}8+3��s"�<�����h��g��/����E�����\kvQ��"o~��9�(�T��$|x֋�ܲ�R1���T́a��+wpMV�O�%��%fz'(��3��؄��
�<�iLB�ă���G��8F�x�O��X�g������n��ϥm����:��Tz��r]-g��eB���@J��7����t]�@�-&��J�FUR�m��"֧� >�T�M����cQRH{�|�+�x�׻�j#��3��m]
��'Z�� I��1r����ov��s�ܝ;nF��M�	R�wnt��[E������U`xEZ�]D�\��>��j!{�{�%������??�BV7��,�́�nWCԇ?�&Ǝr�A��ݚ3o�<v��K~s�T������W+� qf�&�� սF��&F��킂;0��h{/���P{v��*訛)P�]>6�-�Gؤ2Kk%n���?����H�Ù����U�Vӵ�H�JO-/l3e�n`�T5�B�.wm�6#a�$	<xNΒd�<���%�N�V6K~�Ybu����B�ćqQ�;g�תj��M
�n6���yսf�-�`��"���P[�I`����96�������w��:2����π�
�n�{��K>��d}L<}@zj�-m���K���
�x�N�W���'�"���I��T��&�f0Vؤ�X��"ߵ%��^�|CK㽸c�H5>`��u�:���й�\},\I���+�E#Z'6���4`�MqZ��T�oO���c�:_���|�e�OUd,sg�m�S��We�����V�N�C'Yw���T-e�����u��FU���w<��wz�Ŏ2�*��9!�č_��7a�a<�+�K
4��<~43k�ye3>�.`pt�2��HW���;�e�u�,��x�_���iG�+
��F���E�Ɨ;���^
E'�ѹT#w%� ��O�����C��f�c(欈�lX��&!��7��ײ�,�Q��gp�u�/�|�E�$�?Oԏ��^�7�q��� �X8�٬��3)�k��nzZ��ٲE(�,=6J�Ni�9�[�Z`+�NHof���݈���Y�A�����YVv����I�>d�^�gº~��>v�>��ch� ��	������5����W�tL������;�R �K� E_ ����I8Z���Z����®^B�)r�����)W�K8i�P���.?�K��N��u�A�ܟjLu���-r��H���oڿ���f(����ǽCL/�5y�v?yp�V��;j��@���`�4�"�����K�']�����_�	0�4�����W2.)�)��Մ��&���
�G��}?��=��.��*���o���o�/����|6
Lr�x�`z�u�R��c�RA�L�#r��H��2��ng!�ձc�� g#mj�� ��g:Γ
�%�NS�:�6��t���j5Q�ЀݑkP�x�=����X�VǗn6ˁ������4�#�$.*��
�$�D��0⭕�����;]��.�!!�I#x�@���j�P�@�\�UB[U��ۼa<`������]��,�;��S�1kѥr}K�Do�Z����Ԅ�&��({p����N���Fb��u�2��Ӎ��ڳ�I�6�)%:%.�;:G�� ���De����Xf�2�d�k`C��#�U�$�1�j��c�oem�A�lُ�}3��dK�Bi�1���p���g;Amj�L�oe���(Ry���=E����t9�2.WK�a��co�Z�~K�޶�3#�nA
�vc3�ɪۖ�Q�L���Q�Z�HzGYtM7u�f(n�������>�����'y]K#Jj'U��%�Sm�:���Pv_�3-����J��L�����|ڦy�i����QZ>A�xz��[K��e��^:��4/�my;�6'�[F��e��(\�