��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��XXո�S���%Х6��_�����7ONH7��}��� <a��7R�w-*�T-.I�h�]n��[�7ddVOOE���f�*�B�?�o����@L����|�b��=��EBx���}㝱�o�OEY�׋�S�#yI�v���l4����/�������R��$��������W�_-�{*O��W�E���D�'@�qvQ�Y"9����J_&���x�jo�����@:bP@dx�Y�i����刞�QYി�R�fʾ�������sE��$s���x�4�.4�l���!O����i&n�R�x���u�8=,�-I�W�̴ȹٝV�Ֆ�F��}�
�sJV/_k���,�9���9��%�G�5v�9G�&��Ty���uU��+�I��|��&6�%��Z�iXL�[K>�0����{rr�d����oRkIØ[�n��X")V٪�$���ٝ ���|�gDy�ޱ��wgr�q�^�t�U�;)\Js8�Qq@,%�=mFL����dLf+i�Ly��Dm�j���'��Eo��Ԅ$���d�h�ۀ�$���/����k�lG@�`�������m��_	*;Z��?��r�vpɈ�'�?f���k�G���o���[̤B���3����i�úpk�n�de�F�!���M�K���p�o���[B���hĽ���K�����w�ZH��k)Q��*���e���K��?�уӯ��;lř@ ��ِ��nS�6S��7iP�\9�g@�� p{�7œtu�M,��px1��P��W���+Z��9m���MkѴ^�Dko0��S���b��g�ǡ1�#]`����S�_����p$���0_y\W�N���j3��21b{)F�d��C������	�Z��X��l�������i�R�3�L6FΚR�a+�⻇7����x)R��uh��*�\xo)Ks�v��L�#B��|�Aԁ�pC�ˉ�~�u���$.�e��e
L��9D�m��_̡4�52���;��"Z4���?��܋��D���讽��!�~Ѓ���Q)V��&�8��샻{�-j�ND���>��)�̥s��f)/�6��j~�͊@�9u��~�.����:�E����׿ܪ]F����:�{Vsbs��؃��;A�E<��N��5�P���"4,��9�H0S���Z(�{���?�V�5+�	81.��e�X�I��c�-��L#:�(_����pCEy��?���]�j��rH���zD�	�^:K�A�u_8˖�X�#YϷJ8 �C\J�[�m��g	��r9���M��P�Q�.�������Lߨ���k�bv�p�e4,^���ґ?h�5�-Z����s��w-Qx쩀�3y��
g0k]k�������������e��`��l&���|T����{�@�OQND��hUC�@LX�C��!��%�n��c[@`���6J��/��9���ŧ�,/S[ۚ��@�wo�X��H� 2���_s�烟7�Q��i�~�!'xZL��sl|��O(�W�?0��I�����׷͜L1��L��.b�E��4��O��C���KY���2J{qǧ'婳-O��w��3/,}J:���1���	��8l|A���hxZ4�0}��U����r�`�'�����c3I�}�ֆ#Tz_2��.�R-�U�/S� V3m���jL��>3X_;R�Lj(��F\1��6����ٴ�P-���c�2n�Bn�:LC������	��s��-�C�ҁ�n|C��1x[�p�=���+¤�0<t_�Kx=Si��;Ǭ�uFNأ��\�h��^1s6�!i�#Ű�����t��N����s��?dm���r�S��e�qm��,�̶v����B�n_�ͪmi��+|2v�KE-�$Y.8N�BZ��!l��
re�`�K�1��R��n	^Q���X����;�����C��/�� �:(d�����B�&�t3ok;��H$���� Cz�����|�(�j��m���t�h����2"��9�e$5#�p� �$-��Ψ��F�Bv�Y���Ĥ0ޤ�$�<xL�|H���]M$��l~2�y�U�+h�g�p`DA��^�cX~ܥ�(~>���`�)�m�a�KSy�W3E�ie>�ӚΙ�ߏ.Ȃ�O�\*y����Q�����߽�Cf����w�2XK���)l�P7�6�اn�r�
Z�?�����Ug��qQ"�\:y��G�,A!�L�"�����w��;� D$"�oǰe�4`���?�\&�,��f��3�9>	�ʚ�-���p�Ρ�G�F������rß̮2����7�$to�#��l��̡*���͵0�����m��DI#�ᗡ�;�&ל���TW!�ɘ����C�[��.�ư���1D�7�M�u�6z���V��"Q�i���\�PC5'�x����Q�(��P����w�+_��zq�_. �fq�ɚ M�VG��C�����3�x�i�=Z0"��5��xv��]�ѷ�/��}<��� ���ؚ��kzЄe���o�M��ϓ�� �g�Mp�K��_�eW�F�t	��XԷ!���IާW��4�4;͓���fj%��g!�"�@���kt��b�]z�g����M�:�[���s��{I%Wg;��s���-l��l�h�:�� ��#l ��0E��"��qF�1ja��P�}�����r�t�f�	 P��!*g��4�+e�"����N�2��0��f���Ҏ<{�̬U�S�0yA ��}xѣ���-��F���wlѼ�L�&�9d`�g�U��b����?C	��֦]Ϥ�H}z����?[�(�[rt���gC��+?���nI���I9$�.M*$��"xvJ��G�ǳ��`C�&�H߆�P�!��4�BAT�7�/5�@�'��Z�ُ�;7ja��'��l�ktIl���&Yux�3�����J�J�];���VNN���@ܲ�u6
-�p姗��l��.�p$�"��j��_ݔ#�(�d �R� e�%����r)s�O����o�Hn�'��ơ.��us��<�)�m����HM�Z����+�݊k��h{k�=����QU����������St�	,����"8�=hC��_N�)���*$E�z�_�d�U���DL�Yhh�I��j9|жZ�H��4��,�Z�{��'{�@���Q�tR�d)� �}>ul#2�4=�U0Le7q�`��qK��}��-xC3ź!�d�O��	F8	���M�n�w��N��\W�K$�m��p��f4*����'�������;M���>��Y�އ��M!��<I��_ekJvMU��x��Bg�{�D���֬i,�5F� ��>
���t!Fw��ϫ�|E�DT|.Q:vt'��»�������^��ܺڸ�/�]
�Eh.Б�v�{�C�j�|ƨԷ!�^06Dc=�.ŭ��7�>��f�E�7�f���B\��-����1��>O�+=�6X�	�f\��ꆱ!G5�)�P����f�����슧=��uY�;�z�^���6�Of�������b�'h�Y�ѩOBk�1���d����h�M&�.	Tڨ���-m
;��$�� [�����cݚ�����9��F_�޳8)�Z*֢�˿%B� �r9צg��9����{��bʤib�@#
,�'���t[���넷��iʜ�v�4z��CB;T�H��:u�XS���S��ϼ� .��_#������
v��2�$�����_�tZ/��
�Sy�c��|�U�7�$:���S�d�r�O�����.�P����FИjz��)�#�b�С(���y���c�%����a�,���p� E|��p@��e�'���8�<=U�'8`��t$��~��ka��_c������γoHH�/,];;���;�#Z������t���g�Ҥ8]��Y(�����P��p�d�3���Y���+"&���|���.�$�.@�9�b �!��r�(��`왵��8��cP'����� F;�j����ek�� ������*V?x�x��A.$q��z�w���/�;�Z�0�w[�O�7�R�em�CP���M:71��&*�3܋�(��㊢a&��,̸$̘��n�!"�۰�z��������-�/Q�����6z�����a[a�R%Q)`$B��Qe��ޡ8i��{�DpMƢ�{��ԸP`������QL$���])�\�5����|��̇�ҁj�]Ѥ4����GnA�8�|~��f�'��)~�;'<%�Eb���C���Ý��!�>>���u�����| _A�j�w:����p�P��aƧ����m'JZ212h�����Xoݤ�?��}v�8�h76��s�����n�*r����D��*�\\�v'�����\r�B�Wu�u����c�n0�WN
��V@�
�PzaI5@M�|����p0���e�R��J��ֆg�:��Ɔ�
A6��Ї����"��]h�{D�_]&��;�4��'�i�C�P+~ ���:�$�탫ae d`�*,�:�(9,�s�y�(!��۱4�<����� �K�M�L�r�Iq_s�rgkw��K�����_wf�u�0�iXAUDK�=\Z�ޒx�衵���eCQO/a�����2=��O�u��1?��Oh������0���]��(�g��N�Pr�OѴq��|�+�,B"��^�Y}���^��#�S}U�����"��A��U�u��Ub*��`2����	�X�gi��@��	�i��t�s��ӷHƳq�{�K/��	Ҥ&�d|&��Kk{�����a|K���֡��`�گ��C�v8G�[���U^�����5w@Xܬx�q�'3(Sj�1��OW.&6<�Qu偶0�m��� �PI/���-��BէB"
��r�̘Dũ����m��N̸P��W1��>�M�b���3��=h�V�?8���Z��p�jH��ɺT<8��̦uV��Ŷ̚n�[+�QtMH�&l	6�qS���s(r�O���$<GDK4�/e�:7!˗2F���k�?%3P��P`��L8 ܫ@�V����䜬�Z�x.s�1���4{��� Π��$�3
���b6n����m!ǈ�yx���gl�$�{M��|��������o�=+��o~�Nq���~ي�6[d�Bo9(�k.M�<�Ћ7.���Ǽ��r|f�� ������_�bw�얿�1�����!�oH�4��ï��� ��qאq��.4�r�$�h^�Ǌv�<h=�����X(�V�j���/��k��,���e�ǣv�2s��R5&q��u�i��"0j�-p$!�j?�o7������6�\�Nj�9rK�ԛ��@�άb�$��7�I �L�
��'v
��w��m�m�t�ƎH6�E
pᨀ�d�{�}�:ՃC��=���2e��7���:�4�bڠ��PM^hߠ 4bz<R�N%�V`�6�Uon�&��]�5�5k]��� j�B3�\D���5B��{s�����Z���f�F����x�uIa�_]*̥^�r�/���#I�zE�P��≆��NZn;1'&X0�� ��}_���U1����<n���GDZ�Q�z޸�����Y�z��eԅ��cܪf���������$�;(V��A�+O��I����[��RQ[�[g|L�9����N�[�H����^Á�x���ԮW�1�3Ɍ���|[ڨ�'�XG=#��x�p(����]�y�@�c�5W����8���W�]���j��hA�v�h�X�.�6��k�Y���o��;���*#��N��Ws��%7����`��1�r3��'�����,��v���g@�[v:�o��G>ê��p O��U�G���Kr�'��Y��T_�92��H|P��{��Cl��<���<���ё̪��^d��.��m�l�y�_�_of:ɼM�z�k��3��࣮�1�=ցk�EF��҄�~Fxk�����>х4B��\�q2ٷ�`��"����Ls|�ب�r5���s/
U��\��
Md%���������^�������X1RC�����uWӄe���^��<��-0hã�G�E��XUn}⑩B/���3"�,����4z�MZ�̓�������a��|&ߵ�TV�j���8��Ԟ�r�A21VJ��P���^
�adY5r�>((�����e �Dѱۭ�uR�p�!���Pt�Xbd ��R���k׋����ZܚEQ�����3U񁭾�d|�պ�U������G����]������ݿ�I��F��f�Xp1��)E���0�"�sQG��-;��X�Ɲ&��(�b���]ėe�A���Z�d�=]���ˮ,{P�D��Iٕo ��y��lH����tRM��-��v�Y���KA�cW)ݱ5�gF�K�
�ƹH-��t�|��R�MGB�3gf���8�c'ua��]B��\4����.���Y��4�é(���wޢ�c����|3��g/(�8���T:��,��#h�*�����G1u��sK�
�)�&�p�.��,Z*!�`�
(�����EݹHUY#�b
\�#�,"E���I� �7����z��f3�^�i,D@f�-[��9�I�#��s�N5�����g|p�����D
����V`p�� �8!�^��jy�;����/�he}��B�{�Q!�u�Q���@��7pm�lb�ق$�����������R�F��e*;�V�V�3Kn9��, ����`'�T�t{��`N-��!�N��V
��� 	��6���]	���ֽ�����B�|B^�+��)z�R����6���I,~~��Q�:7&C�:��{DpG���S_'��+W*C_O����d���.�PP(<�c�ļ^)B������G��H(�u�W~��~J�#B��~e��Xa����c�Ta�|�q�+-�@ʣ4�
�ܩ:�Β
ojUm�~�0�Zr%��5'b͑e��t�cK��HtC!s��r.ִ�z�X	X�h�s<�p.��[�i�dͪK���>��gt>\��N��!I ��y�S����t7G['��k��}�<���@<L���X8"eP��S�g�v��Tdlp���PcV����$JE7Oib���e�!�NI�5���DƒY�鳽��d=� �sKo�LV{��˿�x)]����7�5�L�sC�#�]6�胙mW_�.��p������k�2A�թ��ӆ?y���%�b!_���l����6.�ns��5	�>�" (�������ts)���"�\�{�{��Y��B�S�R#�/;���/-Z�z�"��N�\����i�{9�\,�p+pq��P�0�����o��חIz�N3n\z��+�\��ॡ��)���=�)@��O�{-�v�Y���H0^5�~ߒLD�|�y���ݹ����;����9n�T.��23
pٯ��Z�\�x�
K2.b팕7�ß�Tx[�RT����^b�=m�򗮥3H�.�6��Y�˒T�2*�����T}x�+�.����V�_�F����1�6�@w,&`c�Ɠ��e,�<�q�ѡ�ա�W��M@����#X���l3��W��o�`R,�� G~���6b�+�����$��j$#Vw��-�>RCrΠ�j:CP��3��4�>�Ff��3W �� ����L����U]z�ްf$��(�+�Ѥ�5�u�C���ǋ=lN�0��'������{�C/�1~q��p� W��x|Tͽ-��sZ=�I	>��C���)����aJy5X��zD_%h)g|�le�7�,���KS����H��m�]a�!�q���a���K�=�Dl®�&v�yPމl0;q�x����rz#7ق��MS�D��e^��m���͕��`�l_J�ۅ,,�}�.Fi^�A�L%DK�b��|3�q<!8�bBp�{�g��BsK����B~w��)�Z��p�ϛi�Ϣ�I 8|���Kg
���b��QV9,�O�!���RH������ 1w�O6�\3��J3�j9�o�R��"bx��������)e�I�������Q��_9� J�����;*�V��`x��`7^Pr����hH�F�2@_�;'�0~��b�[�O�
���e��Z��NA�����Zk�m�)g� �|
2�M �~�I�7�VX ��@D� �W�W6�fC��{�a�q�3����$��h�u��Nqs��@ɂ	�Y���}�J�JM�� ��,�PNQ�Vp��`C���>iZ�L�]���C�����`\�5�d���r+�59���XaDX�"�{��h�ѐq4�r�pe�T0�:K�C�Ga��1��j�:˘>�lO0lo���O�����.�;�H�����2�7���>�5�ұ�-�#�~���;��8�,��`���*��������)(p�O�����=n��A�8�೬T�D�0�����T�n�P?�;M��+�����|�t��bL�2�<K��8���e�����N��m�X��Vq� )y-Q3.Ef��-Vы;��<�g�v�]���5
%�Z��ŘCv	�	)�}�K�&AS��]�[(�mqM�@�U�
�z(���>�#~����ɴ�i��)b..��»�:�LV�(�� T`\�s��!:�;G��[��؄{4}��u3�H⺪���V8o�ů���y�h�����M� ���Rԏq�)M�@i����	�~�6؝p�:�I�Z{���r��7Z?���NA��D70Qs�;�zZ�&�'���.�i�����6bCEp�K�Oza@�K;x�����I����Q��\ˁ�hoC�EOI	��>��Ū-%���f�eud��-������*O�xg�VX�q/���8+ΘA^��>c��_@���d|�	R���CJ��K���Px�"��2�D\�~6D��O�ӷu��	S������"0�-��{ƣ�D(��[p�H�Ba?��f��Iln�Ӿ� ��zs��7����j �X<uzDۛ
p��X"Żs��G���9�QhU=� �������]2�Q�齪%���� � �$S���*|l��w ~X����q��q�򜵐�KkX��#-G���m�Q� V3�Ċ�L}�g������0G,�����B�!y�}�����]�i�Β�Ш��n��i�uzK{Ւl�ޝ��	ћ�u���K�S��^7:�l^.ퟌX��15�FR��]���1rQ��&��6��1ߜ�\HG�m%��cS'�m�d��Oͩ��R@p��q��* ܳ>j��r��{�*A�뭚w5t�(�R�C��2�[W�"}���k]���V3n	e�D">�'�Vs�����e���,���l�]�Kr朹"m�;=@��I��l+�.1�1Vl�N��K$=ۖn��V��9������Rҽ��(,��C�4�C��up(�-�wOQ��ѭbq���$ӑ��3b�+�Uɛ X���\k��KF)�Zޥ�Hܨ��, m� զy�P�,��9'1�L����O����C���:��r%Êu��������%��wN�8]�-Б�y�	EO��W�髆o����*�rPV�`�b�$�xL�~�������h���v\.���Ϟ�")mչ����UFP��nzƄ�2�o���iۡ�Cw�a�F4�qHN����_@��:�;m�:g�bx&e��2�|PkT��X����$_QOTo�S�-�Nn���A_���d�P�U1��2����C���̙�޳im��X���~nn:�]*�����v_��u�]��s8�&:;1�
��_�EUO#ݔI�ٕh�~�[xق����Pҩ:�oDXH�����\rZ�� �h��{����< �q�`-���=���k��%��@�#�p·��%�Z;�Vdb��^'��2���_O� �s7�L�d~�)`��Վ�B�ǚ��	F%m쬎˛*�rOG?,�����1y���0��'��/]�ԯd��Y�e0�(��Yx��P��[hǉ�N�>z����"i��:È�FT�#���5��ʑ-�-w{��������R�D�>���{�古[�34RwBI���I�Qw�40�� ���j���^����C��Ş���Z0E8���S��4E82�\�EL1X(���DϼT��+�Sy �(����a���n~�2�A�U��3~�/��{����6�u]W-UXcsk=���:!��`v�o����ǒv�}�nk�-0��~�z�f�
#F�ޘBږ����pY6�K��jW�:1�O��%-�_����G#��ڥ����|�*��R�!�5)���x9|ч	MD�����A˸�Q��g+��
�L��<��Z���[��E�sUj�ڵos�.��*%E`���n��$�{�͋�]�(�E����+e�W1���U��?ڨf��;潰��7��s�W�X��*��k�嶠[#yÖ����\�49$������2,�ӆ`�@�f��nf�����R���iy�*�=J��pR#�S��22����4+����lQ�X�'JG�R�����k�C�0[`A��.a��,�g����ɮ�"��RK�i������G�[�R[���L�PZ�%�J8=Z^�z�f���u+�_��/���2�e���Өj�6�V\��WU�L;�R�Y��>"�ܒ{|-1�"�����[B��-�A!Ƙ��� �g����/�y�v�؏b���P�yZ�z�0�_;G��_��i�@몰�:ܷ��%��P���g��q�TE��� WԔ �����C����B9yǒֻ�]/���ăv�Q簫��������tuv�њ��M�9ഛS��$\����ab�г�����a�R��ާ�yE�>�?ۣkt��E�'K0#��d䈞�^���gV8�⺢.�����#����]�ٷ��
��ȃ9;�����*��!+5�+�-��G�xr��1�Ӌ������$���'u�J�o|,2A�������竈V?��^��ŀ��L �X�=?֍�9
�'��Q��\��{�U�&���15��i�n�7o����ݥ�Vz��`�]��Q$���E�٬7hji��6��tD���H�>��A�b<tDO?���Ph�>�&b�����=�쭜;����]�H)��8�<Yb����!����T�C��U�)h�x�r��=-;��Q�&B��YwjnE�c};�L�N��Ь�����JE|н�KJ�>��K����sI*�:�!�}�cٕ�/�4�E���9^ M�ȑj����?=�O��nx����2�]����j	$��-XGi���n�L@�f��/^��M��z�S$����BTQ���3�S!���e
�n1�p\M�����D���M4�����O�GU���uI�Ք0N����{�;�ٕŎ���xfz��tΐ��IsMJ�|mm��}nz�TB<�&e(��Z&�7�5B\Qr�A�)֘�եpБ�ov:)���?���S��|(]^I�q:���$W|,�X�<�Fw�p���G]��6ҎJ�����.� 崷�wc9���H��E1 ��U�YR���!�*��+]I�G�&r�qV5�9R�_�4��>����|�m ���3!e�$7W�5�H.�6;)�T�͈�t�S3&����}i��DG�r]	Z��U�0B�)�b�@o��uX �u��ȀbQ��bD!����]�q,�d�%H�m��R�ɈR�'Y�z��$Q�ޝ$Y?a�og��#��S�G/�r�Wlw#n��c�PD'���'�aG��lv]J�LBo����dKU`aϹ/"{V�`cрb�7���6��B,%����y1#M�B{=���M3�fH���{gJ��`�<	`�f�4��i}�����V�|d�V��g�N�+X���7�b*@�����	o[{��ڪ/T���;k�����J<:�:�{��X�֑�bdo�O;>�JɩqA�ߜg����.wTWen��fG�I�G��3��H����"丕�����H�r�{����!�^`e廃��ݓD\X��$�k�q�>7���q2�N~Emƻ�8��bq�[�<������RW�5�'���%�;/$OF9k|s�B^��~i���v����.`����[v��
�H����EV��݈?�k$6Q��gjV;������Rd���(�c茧?p��k�o���s�� SX���W�}{d�:�,�B�sGM(��p�:�e����~&?�P@���,r�q�|�0�������G^K) ���'��q�C_��_]�����=��	��\���HEMZ#w����@�j-P��'L
<C�:a/�,3#�P7�ҋx	f� ES79���{�[@P/�f����x<�8�ì]�)�J�j��q��H�j[\r��Ϙ�ߨQm��I
��;T6$2[���m�2Fb�x�9�5��]�"V!ϸ{̒<g�A&N�F�qС��Ns���i�����r�v�*��%���E��hc{W�*���̯ķ�K >`0=�)�s����>ÉOB���c�$%�E�Kᦳdu���ss�Z�Õ\�0���ӯb�o��݌�)r�� �Sw� j���0V��8���{O �'a87����}�:���=�R�EƸ�|Z��Ӡ�ဤ"e�^�9g�''�ZE	u��ȋ�LBN��:<�k(7��E��|�8b�0��W=^�t�]�C�I��jNJ�7ʅ&�襉�2U$��h{�$L�@�E��.��Ʒ�1�D����d�H�#�1��j2�5������$��^��vo�&�y�:W7��蹄�z����#��W0#�V:<����a@�.���
��b�u����7���u��l5�(���f���=H��1Ȼ�8��C���V����Q���u����Sh�9����\	M���
ퟮ3�����@<:�Q�������ܤ��ц�x����]�b���SnDΫH'hҘ��6��'s��-���eW��@q��I����5�	(z��"	����Տ(��}A6�Z�����cղ@�΅h�d�p�R�N��+�W����5�ɒ�_gF��U�A�{�yɲ�yN�~��`B���y�"l�������������,���w/m���3�[�J��ݞ��k�j����ӧ�Ͻ订�	.3Q�ؼ}��|>l<r?�!r�q�	m��b�?SpI����eT����#C5��dl�H4���$�oLZ�M����J\e�_v��Vk�Ҩ�f�o����u��W���� �N]u���� �%����Gd����8���=��2��J�O�ž-ۀ4ؘ��|��->�8CXDE���A&|�a�����#��;ݸ��Ku�ٜ�y��N��Iץf�vKb 2(h��^W�\3.��U�+Sâ������T����d^]Bp�u�0:��݁U��ΟUf ��-\	*���SX�42n����%1�'�0��Ѓ�1ھ԰�nn�.k��~T��u�Z�Ј�f0Z	��J�2d㙅:"LA���|X�#�����t��+�P�quT���Yo�d����}�@l?p�6��󏖄��1�g�[Ѷ�oHX*6�y#2��W��R`>���Pe�eg��3;u#�Iy���M9=0�GXm=���t(��xl�;��e����n��ye�$��v�1���IzRG3�/���F[���?~6��E����}�9[cl���2���]����ز����k�c]M�Մ-o� -��!#��i���6[p������=S�g=}[���������W�]?Za�������T��
��]�7C����,>R�)<�8v�t~�k=�Ԩb��֫|��J�"�%R-���C:h�S/�3��*kf�.!|��}FK�y�J8b��(�>�,��>Z�����'>��f#�m�c�4����gZ��6�V��uy��1'��I�@����8��ˋ��-~���yC��P�c�v�jW��Ǜd�(�īK��GK�*�"\[׫��bI�KC����-ߵù��S:C�ؗ���0r�����*Z���y���Г�D�t̏�K#3��˭}�#�e����5��,��Ș���*���Ot��c_"�AqN��@;)�����.�llh��~�Z������+B�wP��*7O��Mc蕃�`[!v�����F��M���9�޿��a�b����P�b �g{y>$���Wi�m�{��}9
YJ]B���
,�F��t\��0��i�����լ��\��1V֍�������C�ӢW!j��/9���.�9Fx�^�U?-N��r��4��V棈��y=���t0>��/F�������Ph��r��l�MP�XB�MI�+�S��f���CKC�K0}����.�U�T��3��5,�yP��,��;B!�S`��
O%J*��`�j(����Y�^�h��g�+y���7�&Xd���F����5'>W\�=�e|̌�Ol����>]�IH�'|4��?��|�;�/F�/E@[�Q����$�&��ge���:�Y�1T׼��'G��&R
�(�?�:�7Q��9\��lf����vkA�F��[�n�٩���V 	���- պ?���oz�TU14���f���|�\�I�*�X��Xn����ظ�ds���|w�;tRx���-$�)�W� ������e� �L.�4ma �B���گE_(��L[�Ξ_6&�I5�_n��	��J�A�������꯴�I(�-�\X���xӍ�J�-��uq1u6WNOi��4�(��5�(>�Z��j�;���C@e����=�	8Wy���U",��=D�JNm�'����/��fKO3����j�-��
�,X�&�h���V�=�S�Y�y�������\Y�д}vr�1�����>�X���"m�<k���k'����8P7�+�*f�N��y�>�4�>��@n�V��J��Kko�m������u�ݑ�X�#*@y�I��Ӄ94�m��� r<}q{���f̴�� ��Y�Ȣ��	H�����~�J���^w3C@.j'݀"D��&eL���6���|M?a�D�(�õ��Hj���;ꊦ����e�R4��ӗ��xIԴff����I�x	��_��ۓB�["�լO�\�-�-�����[v�.; �/��I;S��Pe=_y=�����$�C�����A,Q�Ӊ������uv��%x=���Q#�"<;��%�5��&���o�7�Dt�g�[�Y���9��m&F-鈭�IM���t��$S���L��s��
1Y�Z�Nf�T��1��#���-��䐃*31W�4rt�y��`�c�n��&��L��Vq�~�g�y8�V	2�R��%�Y:��;�=�8Sj�b��ȳU��J-����D��N;>{�|S�oﲱ�v0�aq�壶���+�!�j��b�k�3�o�����ż�@��d*�X=�Ņ�MT��!���͆4��.5�V��Z1���!��3� 6r���t�-acmv�$�54�����P��1Z�
Q}�(M�1c0���G
�i��8�6�.�>}cF���P'�.�%  V����'�n�wH��F\,�i�eYgs�x�������f3Hp1����G��р� >���VQf2�$�\@��V�ť̕��y�3^X��L�7��rf/���i>�v�����RYt�U��V���Ý�����#À��3þ������Tyb�����.9|��U�՚5�~���\��D%9�N��/�t�x�!��XK�ɯ�����p/4(�F��s"5�C���u�]�8���~�E~���^:]@~E9&�/�7�𘟀�T�
����q����G^�D�}�6���%<���``T��3Ύ�sM�u;����;�F�zH"<v�S�Y��kC�Qt�g'�@���*��Z%v�h���
@˪����*֖����BT^E#vwY�X�J�V���0��3�d���2���x�-�a/���V��ORXV��LX���� ��`A!]v�ݝf���;<��PP'6Y�x�r]��?���P��1s��S�4�ģ�:ݔ)�x�#]� F���`����-0�w�~h�Y�#�V��0�ݤ ��+��S�)�9����#ѡ���XZ��Z;ΎO?j茶�;9?�����r�GN�JJ�&R���z��iH����b;nZ|�l[/�#.��D���s�F��� Ov��� 8H�����-��f�.t��m���!�U$� ��?J�ek�צ|PI��ҙR�#�K�
m�;؟kV��#6P�Q!��n�����`�Tո)�/�F�s(��m�K����+-Ңa�������Q?52�|X}n
(}��-c�"�8��&/6�-�hHHq���c���}X��A�tIC�ɤQ������Vi������D�ERu��w�,�F�#�]�͐{~5:�2& J����.6�=^�"�J�X�L� �8M��'���r���)�h�w��EX�tf��АRFgK��%�P��bS��h�V�Gd[��o�Nl�f-��Rl8�1J����n	���+�ؚD {8�@{եS�!���4��@�^�^V�s�ը�-m83���%E�ؓ�km�u}��Z�o|�hw�'>H&+�v��h�1�n���R�Ʊ�]T�r�L9��Z" #bH��
V ����.,ژ5�!d�Hߍ�|g����f8�H>�eP��HoΓSҘD'����|�]�Ăv^D%^Zop/�`~����d���X��J����ہx�=�Q���Iw�V\Q?�5>|�ZYU' �����r�����:}I�8�A��h1؉^���z�UP3�H���%GM{��Rpb��%��8>d��$:.��������3O���R2��Õ�.M�t�*>l��I_�t�Vd���W�������&E��}�����ۋ�Hվ������2�$�Iݸ��LlÕUV�2%o����/۠��A�P(��C��
��rA�9�d'�l�{�4}��%���#	��v��\��bZf�@�S���&VR�UnCY[:���m����f@u��b�ǙnY\N����O��W�>��}���ݧ���U,W;�o�>1��%��f�C�"�o���v�as��\����+>�Vt�O/sa��yb��e��@Um%
�Oz�c<�՘%�;���@�g�z)�T=�y
�z*�O]{z�a�,(���~ϵ3bw�ͬ>gs���Y�
�&]ۥc�Ԗ;ˍYi�,la��B�.��_�nեq��N��	sU��9�H_3�[�b��P�+��0UY��U��D%üj��Z>�ٍ�!���ÕڴrˊwȻ5.��=S�HH"�����*8�R2� ����#�t#�
�Sg���v$?)���ndn�,��t4;��hu)�|/< D=����[L�00I���@��J131:�҄���;��'7��e� ����6��L���?���k��$:!�+6�p�Zxݛ߉�m�UG��q�� �2����)�d�c]�`_��=*_n�|�������K�� �RvIq��7�(.3�hg�X���Z,]gsBna��`j��{u�rT��9��~�k��8�m"e��^�c`\�ix���,��X��z���8Un��o⢮���a����y&��`��fv�K
t�X��wM�ϭ��ŶH
�k�B3�SG�7a"�b}!��(p{� �r�̱��KJ�{�R%"����;����X�+�K��=������X�K�:���8e��3��/i��h0�.Ds}������!_<�Z���ߕ(�	Ň����c�Z�7�7�9\2P�q�!��Bl���$�p��KT/�������D�'��*4}L���y_�*�{k���$�[dD�E����:�h�Їxs2�J�x�������)�޿�_v6��rr�+��IO��~ʜ�7@0�������Щ`���FJ~#���{6��U��a�)2�3���P}��7�*p[�1[PpNU����a#"y�zb��"X�Rj�`�K�"����x׶�=�܈*Ix�t�*�+A���W�L)J����m�}��͚�A�����~Q캱J�5K�[p&8���F���i�tP̸�: �\���gf��,�3q�j��4�iU��P�����\Q�z����>6�K�����QL1(��cY��1<O�EYJ�������r��&C]I~�%��y�L`�+qٗ-�;>�Q�*1�`zv�2/�d �� l	ɐ�F8�j�g'ISj�j��ך~+l� 3&�\�Gg�O+���;o��}ݰ�e�B+�q�O~L5��V���>��Z`���{D�N<nH��N����I�u7a����
�{%a�/�B�����hP_ц��$g$TJ�J!�HV)��j�Č����g����X#����Қ�h1n���_���XF�} �\�7_$ܡ"^�y����r�e�8�x�_�#o_�wo��o��ɮ�����(,ڊOBauB?�e����o�B\��� ���`�
	c�e-���>�D�Sgu�q��ѽk�Ћxщ�Nq	��&��ߓ	ئ�������q��ۺ&9df�e	��1k;I�E��m��^�Mf��(}�A��Ѡ�^ ���?V�+ʖ=����潻C�P!@�+����g���ڇ\����C2W����"�KӬ��8��$ɞI����S����+]��ؾ>��"3�9T�����dd���a͞�>�θ<�2B��;	�hA��̨u������*��M��'�����3C+6�.����#���1(��D��!�[��'���A�
`������� ��Jeb�[y�Ƚ�[~Z]u�	���֡�_s��v�$��ޥ����K����?ɣ\����и�l�U���ֻ̺��KkC�/�ݫ�,��\%��3z:*,f�9���p ����p#�0O%^�,���Y���@�nr_�	1������8��3|�7�~KN���w�y;��^�o����ϲ�$��z�����({1��#��U��\(�DM�W�Ƌ`݃�V�L�G�6O���N�l����S4>s��
��X��C��0���ͫ]N*A��J���Gwf�V��,~np���%)v���;�g�>h]��38�ȤN,�a`-�%[���Ρ&�&K&c6P'!��Ve7��hy|���S��+�i�ᣈf0ɭ��u�|X�y�+n�����1�̱�h��d�d��;�N� /3��x�8@>Jb�(U#�Պ0��_u1Sg����-x��c��W��}����DI��fo6PD�
����c�TƘ]��=��1w���ʮI�7�3�LZ?�f~@9�a���;X�9 m]�{��u��o���~�ɔ1���ǯ�hdN,�;�<[LzK�1d1��9�Ƈ'�kC��K}�A�~(����@5q{�w~~�ڠ��J�zr�RT�Fm�zV�YO`�IW�S�mX��5R�S�U�T�Y5��J"<ҽ*gFʵ+��^oWk��{���D`}�5�pD:?�)\pǪ�,,��O!�c�9Q_~�i���>���:M�H�d�Q�d�����R�g�D|Tr_���l��U�����f���7��hɭHů?�U�U��Ko��x�G�L3/h�<CWr>����б��Gn4aϕ�$�S��d��^u���;RO �v��0f��v�0O��A�㸺 �uݫ�FI/ХP�dA���Z��62���ApmF	f@�Xܰ���Lx�t/b����P�_�CYy���a��n�PM�B����9���,pj�P.%��e"mk��k�X��{�脙�~C>Rd)ܞ�9�zE��ts���^�0�O���9���pX��Z���';ۓ�~|h�hh��J�0nT�:3����c�����WR�+��!й�0@9��U�g�ђ;����2^c�8^F�#25Dio.L Z�� �z��D,JJwx��5�=��?�
�ÆE���Q�A�[��tߟ�� ߜ��e��Ck�i�� �f�R���J
��_���LU'ܢ�~j��}�p�MF��3{{��Č��#܄�V��C��q5�L
8~�
�MT�d��n�N%-�.��hS���ߛS�uAOYz\u���w������,7�"ِ�^q����OȆDn���h����S)��%�wE���F|U��+��^�dl�F��~���u���:��@��0��)��Q<�F�;��t|�=K�ؕ�%I���H���R.j�6g����n��wk6n濧1���<��0���$z�qE�����y�1� ��4z����Wy�>r�5��U�ڡF��V
��&�D�4�K=69R�X�E��Z�#`x3�A��娸�>_��!�n���T��{�=��ۃ��+�%�]����� �K7����d�5Ԧ�1�����P��]L��!�%�������v.zd�{�{}���u�c��$�D��P�DV��MH���QU�A���`b������4P��� ��/��-)m�#���l���a܁����z0�[��e��A�f�f؎�s�1L*�G�`��� s�
<��Z��@a�.�h*'�C'�)����;��ig�P�����.Oo�P�dx>�`���%��-����iG̭v���(��p�S�do�lC�,xd	�.�i�s��$AH�g��q�9��6֙qi!�O�����ƚ9򑘇��?����3��m��[��e����}ķ!�����<�(�<�Mɥ��r��=ڕ�,&����� -Q,+U�l��fs�g�,3�$�tsgaY<l��'�tz���m҃��ǦsM�2���ӎ_����m�v�@D�9����m�SV����G���.�\c�(K^�H�	
O�"�oxÝ#�8��������4>�P�A(��8̂�w�R��
���ˤ�f�"d㩃��Q��0��ۥ^����+_\�b���חVU
~[:M9���n�Y�	&�s��B�>~n죪&����ů�Ĳ^�A��kN��>j�*�9�JsB�d?�p���(\�,7+aD{/~g��#�-��閥�k��<�n����:4�5�e�X'B���%rd oF�}J��t� <d�f؞�8���ezW������F���C�4���b����Y�:�����7�k�W�x�dаZ��/ˢ"���Ln��=F���eW4��Ƃ&O���Qu|�,�����6Y�����NW-z�T�<���l��DCaD
Ko�m��T���u�H��M|�!a{��Ʒ�A��c�p�ѡ��g-,�p-�@*�B(�0��n۟�Y���?��.�)!u7Q��D�+�V�����q���+J� �A ���wFQ���in�m���}�pw�A��=8�_�]�v�nYƆ�EH⪐��{|'�h�E's�Y�*���6��_�����@��c�`��|�bf;��(�H0��؆L'BK�|L����q
4�)*�Ҭ�pKbc0O/bKxu���][28�`���C n��4����[F����R����>�*��v%�AMB�	��L�A	*�3Tw��~jZ��k�Ӹ�4*���s�,�hk�u�6�v�V�Ͼ��Ĝ�G�����vk
�sW8�Nd������� ������YMV�M���5r�G�L�ŦA�iA�3b��d�� c� �\�_|n�'��H5'��!�Ü��7ۭ��6�c��i�bY/�-!�P�C[M0E���!dʊ#G�Y��0I�%�+zcDN��f���G��!DS����#)k�8}�a�ݧ�S]=��n���n@LM�����.���(�Ma���L��/H��Bow�o�IO4�Q�ښNO�C{@�lj-�et$~B�l<�%.�1N����+����]a���u^��K���� o�kl���w%p�"[CA�Mw3�="P2 �Q��Hig?�����,�H���B0���2����L��M�*D�"ڌ� �JP4k�~cSI
4�6^$"��&�,���n�^]�|�$<��H�"�Q��iK�&�?B+�jP���Ҧ��L�C��1�p�VFH�Iy��F��ٶS��b��X�/�c9v��"��}��4��C�j���0��W�9��~D���r��
U���EZ�e05F�2~L=��1�"�I��rb�+�X���K�=�&ߧiZRq�����y��\K}ȝ1[4���	��Z�e�VJw���i�;�M�O����fz��;��+s�64aPA����������Pu�5�-�7yU_�g����5N���G9h�s��]z�)�Od����\��S%�>�\{�w��<υb�r���< ��+�"9N$����^Q�[޽��� F���Wv.x��G���5�<t�K��uîpC��w�u*Of�?)�O��ĜZZ
M�!�Ϣ�W_)X�}��dvˠ�]2k�M�@K2ha5,7�6�	�8v-��fQ�Q�����%�et(غ �����=D��)��7A���cV'��95��@��m�>g�MNaa&v�������lU~oںjh�PA��|9b?9gW�����J�#�
j���T.�r-"�lG�ڧ����S`C�_���F`8C��'�cŤ.����G��K�a�µؗn{��ħ�A���w)�9��os.|g��t8�C?N�xe��%"��p�Uԍ�B�:sKO8t�9�ʯ,��>k^�h����t�.ew$������;iʷ��[�2a�*�	�XN��f.-��i�/S��^v>k�˚�[z!��aEyF�����a7ס�UfGx_ޑk[4���%�J�Uy*!��&�K�fpv�Ԟ&�1���t����B^�u�Z���A}�z�Ӌ;�7���)8i�	93��'1�[f�]�dVv�s:��W�)������"a�y�?��i`��S
�������_������ѱ�ұ*)L�.��))����Q�h����f�?!q��1�5�� �*e�H�Z@�o �)���o�?�e� �Qe
���D���'�,^��bR�$��D�-��+ ���@�z��z��s7!m����k�T�%�v�N�p���?�Ÿ[�
th��b{	S�f�xs-����R(���Q���P4{{)�5XTP��f-�8�����4~�q�Ƣ�+t�������`�+� ]c��S����Y��KF��s.K�c�֏9Q���SDb�lF�!{a7�0]�-@��:��yR��ޕ|�A����uƏ"�J�=��y�R���󶜯w%�y�T�H�Pe�u��c|z7k�W���N��9�կ6ͬz��Ї(��#Y��it��ǐw5پT�������d�B�x����y_WL	���%#!{I�����0�E�B���S������=�����UX����ā�ȢL��!����Ew����s��zRG&X��!��G�#��?�!6w��[;K������K��O���Ϫ�c��=6D��8�,,7�#]1��@w�;om���:R;��<E�&;�N�):R V���ss���1����|���ɜ;�q��z�~z���D�_Q�|����1���\F>�6����z�u���_?��0�n	�z.�2]�|:&�yG��S�����R�q��Pa�1�4l��@������"@�9������n�,Վ�VE�Jߡ*�G&�)$�<5�獖ڣ@k&l�����O(����S���	�qi��ژB��-�ϥ�s�1�|h��]��0n���W��l�!ְ�K���PG��$����7�}`�:���c]�n���KW�z;5��u�6��G��|AU�N\���������O���sL�G9�A��6V�r�q[�C`�?Wd)����q���W:,I�s�������� D�m�q&t~�9㦕�,7H^3����f0c�������0��k�v���l/�H,yO���P�'�H���XԐ7g�s\�o�u�h�thX����@�R���֜����a�},w_�Is��Yrz�m��ג��࣪�����O�^$���l��/�:�
R!s�������ȩ�[��DS[��Ra�_��炃�RbR.P�'�ǂI�8�a�������kO-�rmo�)M8���~��Y�ciڬ6�R��wS��
%��A2�v�h<�Z��m�*߰)+�aQ#8?�m��.w�r��dp~M�@q�� $�]F�#�������^���7q��L)�D��ڥ��Y��V��Q��|�mP���k�|uy�@��]n��E�z������Ki:���US2\vD�<4h�+L�u��C��DESG&�Ѐ�N%�<�����ux�2\�����d��ڡ5���*O-��e��h�T*�g-�f{������ur"�≅u9v�\�U�,���"�D"�Ċ�D?uf�c]�_P�vS�-1���{'�$��S��q��("���9I�LI�x�B��ñRV��Ԩ��7�.�E�`A��7';�|$��X�l�0�eߦ�MrN��`��隷�H6��6��<J�yH5/��%�e
#H��4{2���Ne���O6ߺΜ�_o� mr��D�N�=�˲��u�w�T��$
��a���^�.�E������2��nP��&�m$�X��`�"C�C����o����zxx�)�C��Xo�jf�{���i�'�8�Ltq��f��[S�5T���f��v]zy����?/;�\uO�C0~���@����h����z(	�����̫b�����LU���{8H� �P��>�M';[H�M�4��*2W�o'ah�,kN��͖��I3�>V�I7c:e�e=*���8�&8���[+����Fym��q�G2�E.����xf��^:�.�[�u�?r]n�HG~������@Zn��B}����	&��a�r�g���/aU���j��m�%}�cԺ$�J��LH��w[��n`?.��'��L�泧���n�+���Z��xؕH:����.\������Ȯ��QH
�����l=��	�8������U>�r JG��Z��Z��3�UY�دo�e1gt0���cT����`Q
���
&1&�-�*��]�����-3�MJUc�X(�����*�H��X��V0�n��X�z����&��ش+Ȯ�m���ם����GT�&Ňg�'��.R��
֊�H\t�k�닪��������@J���3���c �UuE�B:�����j����'W�$y��,c(5��߇�md[ŵ�:��ށ&*����P~#,n���,�4y���vɆ j}.�|G��9��������i��|g�K��E�0��h|"H.1=�}Uqb��C�d��Bv����A�t���z��s1�g��M��Nm2���ք��=k��CH �P"P�N���ku��g+���	Kvh���KY��@��Nl/��:b��?��_,5!���>8�@S���#���3M�o�,���z�y�Guc���e��!�Mzd@QD��J��P�3�ol$%!��&[�����9=�:k��R�Y��M Y��d8�<�Y�6⚵��X>I.���%HB���G�%V��+�t|5QW���k�� ��$��1нn�i�X�/C��]1~��b�-�aG>��-�W(��kUGS�&�r���<h�#�d��(�-��Z�g���thO����;�ʝr���9bs�,�oS�Xv嬡�N��26�1,�ܤX�u�<2��^쯻����N�=�_xf6�$��AL@��@H��8����C�+�<Bx��'e+���Ng�)?������hA+�N
*+�>��9}��r�v>V�D�V�7��5ފ^t���i���憛������_:�uO����!��P	�,+��#ԏ�}�[	�s�1�s�%�t2"�?�W��hX����e�����Ju��GN|[>&gۛBw`�Q�Aw,y6IK�z9�`����޳^��D k�IX�����\�̗�|�7��g���`�y!kDԘo���Ft�O#�S���|����\�u�h_Q�a��
G� gG�@�ܔC����y��X��u�Pތ����I��(�P9)Z�~�}�3��z��'~!8�e|j�kȶW�vl��}�Ğ�bD�TE'��|*�<�ݺ�#Չs�+'�Y�� ����"�W����m�� ��(�g 9��v{RŔ�
�j#���]�1�<�ca��j�Z&�vсKk����M���.׵9�)��Ƅ\r=��o�M��pry*62[�L���L-ؿNo�R���%Hy�nx��/��t�k�{���S�ޱ8�V�-�9�`��{#��^Z/2���(*���O � pMh������pk:�:��s���j�θe�8�*��:��e����Kݽk�i��w����N,{�F��c�'Q�U����ګEPb�ѫA��N���(f,�r�NP�mW��w��*J/�'���C�(Z�h�)���]�,������h�)8o�af'��n�ԫ�-��N�Ji1�EO�RA 8�7+���W�=���k�8+���1���P}3��b/�J������ա��ȎP��~���|�:��ôo9��U^VD�v�x�e�1{����=�myf;����NW�)rc�5+�]'�5ܮ��RnGZ�:m>F%��`�i����O��B����k|���R2�)\��n[�*9��Qy%��=�v�Z?{���H��P�����!^��H뺺�S�x�9k�>Z����`1n��eS�"�a�������@�0�t��a:�����$�e�`���ңsi�̥�Ȫ#U�S���fӫ�����-����<��������3���g�u��ڷ�K&ʾt>��8�U�Aa���xvf�#�y�d��wyH�p��?�]���g�q���~�7�_�|�T�n��r3�Z>�Yx5�ɀ�ؓosD�/�P8!#��K�in�ț�ۇJ�� Yb��h8�J<�)�`頁,��U�����m�%����[�E\�ew>0��ưD�������/I}h)������O���Waksvex��ơ6�K�bP�i�-�":�c�R��g(�_�62Ӌ�y� �:������w�����m]��I}�_/�xMU�*��<D��)?.l���In(�J}$Xw�!�`2UG]�:�J� �nô޾�B�
�p¢����˂o�y
�?��yK�,m���%w
lt���=xU& ����a��(g�W�:�?	�Bu��;w�7M��MQ�������H��N`���%v٧�p���O��!$+��3s%E�VəԻ��ؿ�l��FW@�E��t���j����T@K�e��T�K�F �#�j,��(��8�~����?m�f�#S�U��?=�S�J�����+T��6�ap�z����ub@���n�D|O�7R�ȺY������e���*/���xpB����2���+��Ov����MQ������1��;��2o�9�Zj�/�C�Qv�5қ�SZ+\���/n�հ�C�ܰ��#�BO3�yHs�.�������Ș��s推�}!�e�*���^�E�����L�:�^}8�E��j'�b<7$P��+1ֿZ�Ǖ�t\����A���ļ�~��#�g���g��R���턪���9�!��,�ۉ��#�Rq4ORɿ����(O�c���Iz�m�r�bqX��9�z�z%OA���Ց{�T�	��O�k���T1����.�� 7e�����Ž퓧,#t�\�/�h�Wu�7l�c��}��>T�����Y�]8������p`j9Y���Z�-�GS�/]����g��0��u/.(oGѳ�,ifv��q&�J����g�M��b�<�˱=�>mbm�S�j%ǧI�������0>S�U��';�Vi⡝W$sM7�սy/�`��b��l)���&~�1�N_ئ��P<���,�҈)�ćUyl�h{�������6�a�D�S��]u�`��}l\����/կ;��2.�	Ki�M����Y�� h���+y�~ꉓ�P��m����{褟Ц��^U�n��˅w+�m����,��6f��oi��5C�UH�>Xi�9�(auʚ�����0k����Ur~��|���ЮMg(׊ƹ�zVɈ<���~�d���j978����S����cPRJ�o3Q?~���s�f|���_� W�����Jjo�+��,>������S�����e�Y)ؖ�� ɲ˵b��r ��wn����#k��DY���!�������|�%r�\�����o�k߀U�EɗH-C��ݣ
n�>���s,�6h�"6�/
�21����D��1ys�Ti^����P�S��~�h����9��Fi�瀆<ρJ(z��7�Uu� �A�VPn�2;v�tw6�	����_)$�L�˺i0+ٷw���xI�R	��w���A'ט����������X'N�h�� "�!��g/�?�ǜ���xj7s�R�~��7*7{o�F�� \.R������e|�x�_i�,4��kt-��><�0K]�������dh��q��~9�xl��d��J#
��$d�u���}Q��rР�6Q��i%>S}�r΂#�;zc���K�8ɿ��j�V'IeY(� ��(ō��<�~8���s�у�6���*W��Z�X��D"f���X}�߈#�g8�B��g%c;����ݙ���"�?:�{�� 5"�'/ǜT�Yx%��,�%����N��z���W�˛��;Cz��aV��^���U���* �gUm-]���U���P�|X���Ϊ�e�*��m���Վ��a�/*�GUjW'I����Z#��CY�-��w����:��~�y��d��I�v�
Z��-^ª�h�����Dl$v��Z��׬��N���z��������i.ӿ"L&
���Z�hB�N���i�1̜B�Z����yd�.P}������V{�V�j��&F|���PD^C����Z�`'%�������.q-ԉ�Ė�.�Z�F�@���X�{�¸�����P^	ऱǤ�zW��qt;1�S{��������6U�����퉢�W�����9�G��& �bt޼�gWŽ��(����Z�@�`Hp�ΔG��+7\���K�Uq��\��-�h6�f`,�z\?��d�c�������[�c�yn��D��V����c|ag��ݫ��r2ۤ�Cg�a��w%ldv�La�SY1��J	��1q�gQ�:�-����?�w*�U�˱S�&����'q�X=Ƀ��+B���r�������4���wg��L��aH���FP �����T�������!6�L���S��� ���p�lm0�u��y �?�����ﴟX���6�,��EϔȤKZ��8U59��<��3Kz囙- ���`���'�S�↴T<��X�Z�34��|�<�`�b�N���;K���ܟc��t�`�&l`a#Kg7�}��}��nyK{ '�Ug�/:gB��� �k����u�t�w�}(�9Z�k��6rj^ԕ��ɂ�K���'��mטI�m&B�+}���N�b�)Mh�WLZ%�󪳰:*���1qi��� ��H����[��&r�B�FN�9)۩��Qh��E�a?&&�`�vy����]5���,��D1\�fW����O��t�0{����_���L�L(��q.ױ�9I%�4��i�,�{�W\��w^�\���+IB�Ͷ>y�����s����yo��"���BC!�pڈ!���2��Pd��C��7i(ZC��Yq�N�ad���NA)b ��(��$�����O�w�̪���B�y�m�ȉH5�����3�3��"��ؾ�I)dg�y�������f���Tނf�IL�3��y[PV���U�ͦQur���l����P�+vCsc0ys����)�[Ӣ��ڱ�z4�7ɲ~�(�K�8��t��K�#����{@��	�H���uR� �S9�V�2��yuQK����*&x`<��|�_eK���h69��P�J¹<�6�v��?qz�~�p`�2߼���JT)�CN�Bvs1��x���Knu��h� ��О]d#����OH��h�}bC���z\l�h�n*��;�h魮��V���)a�u^u@v����2s�W��% ���T�|��B�R G��9��҃ˮ�LV{A�	A�3͖��]#6�Gl.�-}�aEi���"˪�' 5Z=P��z�I����5a3��t�T1kg����r���� 
J��q��Zl]\�r-}�XaIu�5u(ӕ$��?%��p��&��W�Dl�>S!�!/|�s������&��}��$?-��7`�#�Ы��HYR����QgVS�����2a+��c����b���S_�c�"j���G�����hEvD��k�S����3I׼",B�+Q���̵7B]X�����T���K$��Rϝt�s.7��~6]R�'y���&P���@�ހHB�뎱��"b޵�x�:�K]��Wa��0d���鼏�p����?�>n�	��#1����޵ .>Nnp��o�Ö�h����cR���+���@�����W�q6U~a�?�f������q�1>q��_�����ˍJrվw�ڑ�j�'��X�[.����ާ�致�}�������k���Ȏ�S�
�9٬���s����t�@�d�&�^��.�Y�H_�V�����b��e5W}��R+&,=���@���2��m3I��L��;5��2]�i������U��1��"��L�@ے���O��[ܰ5��l�+���еNG��rr3�k+�6�]+=sA5=�v��N|2nm*�;�0ɠZj֔���e��A���~g�7�Sw<�k��@���VE�3���w�<�:3 �0��3�Z�AB�UYs���t=H�1W��P(%�Z�
!��o���u�f`ɞ=��+��!4�8V���%1�OfB6���ފY_�o�Ή�kB�w�c�È�;����o!�?:���8�I�y����3d���ո;f���`�O���g��2��[B�N��Y���/R�M|�=��Ti8�6(�O��g�
s�Ut��X��H~[E��&w�(�6+��:�7Hڸ�7����T�h��{��հ�pNu^�7��3MǑ�^n~�����0���;ln|t�!ӣi\pb�{�I\��Q�	�ܤa�E-.�`���V�B���ŃABp����DP��}���-��Ob�n�����r
����d�ܾ�������:#$�w�Tyg�f�V����R��%���`2�%� ^F�4�ׅ�)*Kb����`��2��_��6�SL��H&�6F�AfȌ^Q���P�I7����'��G�j=<�����"�z�+���Mc����;l(��#�!ҽ�+�q�v��ԓN���1�˿F�����qlW���Go�{ߞ�<�n�N�>�l����X:��_=:�ɱua#9!,�Z͑�'�u�.X�)��ɨ�&A��g�c\	�l�|�!aw4(�4]$����-��>���J��A�N�y����?wbꦌb�>�«v�}��W�ɱ���.�x�c	mȩBl�~�U�H����zu���E�Cۺ1�ϥ�9��~E�$��hԑbf4 ��1f��Р9Sd]kAX������'�2yn�$����L�%k�u�|�DQ�;�}����VG�l�7�:;��Ś��$��2����Ǯ`����UF�0���J0�מ.'듽�u�m�zM��M<�E��J��"�����͛����w���d��m�vC���I��*	r��1(���E�ov��A�ph>E��L��vK�e8���2p���0qEx�2rb�G�p4�oq��ݧ��s�i�t.�L�N���^`�6�^��:#���nJ;�x���>P4�g>�����'Sy����˱��{@R���ݮ?Zܘ�'�G�s_鰎m(�H��_h�6�.���Pـ͈*�6�I��B�v���	-s�R�16�"��i�+���ɝi���u��xs���������!S�W��we޲АM^�l�㦁�δI�㞸���2�]�z�v{ˠJ��ޥԏ'c���Tl"��3�p@�>s~�����`k5�#(�ɶ�N���*>����8��E��U�M|w(�U��q�XNˋ��|LoH��-��8VeȈ4�<ݑ +ě���qDH�@@C��J����^����wѹ[аi��v\]J��C�Q�������b(>!�P��?��ڷ����ۈ�������H�fp�I.~M@<$[�O�T��ZAu����I���T������u�f}���7�\�_=��tND�\���6`����$�'��V�ِ������ Bd��.\�.O?H��	$��~JXA�����������z���1��G�g೛9I*���d8&!7���~S7�Q�_�◂���H��/��v�������i��Ap�WL�r�:�F������!�M�'`!�S.���-G�2���9m�����h��X�|N��:B�����#7R
I�ԍN�e\����D]��^ˏ���VZ2`V;sdz�lN5�@�f�N���Т>Zm/����~G̑.n�s��q�Զ����{���;B�yY�'�ᕤYU������#_/ �(dt}�`8?󁏆2䶥L����/�dp)�"q����B�B�Jdޕ�����C�`H��m�8Q��O>/1Z9 {aڶ��
u,�<�o�Kf0C}�r���w��m�M�������&�n#ٺBO^��U��c-iAV�\`��
!�V�_��jK!�����#��\0�i�pv*��SHvX��^n�uͲ�!�+���펁���ލ�`̤4�5��gD�=8m	�>nb�Q]wK�M*�ֆ6�I�9���q7�(�]hL\��Ю˩�y3�s�~~i����� �o�J���ga�Ѕt�k��:"�$�Ǵ������d@c$j�=b^��6
l3��m�&��/im]o��I��ʫ�υ�;<�Z�&,�f�p�Ӄ:J)��	��$��)��C�Zi~Rk�)�/��Gz���Xԇ�.�����wm橵�|�Q=q8�A��)�=޹�Z?uMۺ���+������Ҥy��[���F��܂�4��t���l�E�e�v�\ Y�s����ҵ��5]�I�]�͊���֔x��`�}�0��8����@^q��]�s3Z�ĴP�ʏ��eA���Λ�O)p�R˛$���6��a*<�_�2�W�DeK�w>yt�J��\�)v�7:NT�U�"(�s��$2J��E.�i��3\ŕ�i�`H^�{(�>�2��v�k>%>w�y�8*@g�7��TB�-<lAE��,ް\Z�w�pc�������՞��a��� ��{���:�bAD�E3ن��v�
m���G��c��Ͽ��UvԍO�^��(5_��=Jm���1f��e�u�Đ��P��2E �������?-��"=�v���z�?�Ƕk�ez���L@a��{zD��2Hw%rg�D��J��{����2V�Y���VV\��6���>�9{��UL�@e�A�6����W���S4ϭ�D��+(?���m�'�l��T�Y{��w��0�nSx��N�|� [q�ې,O��q`#s_~I���έw>aL���I$&��E���$��C�T�UA��(���J��  G�����b�aЁ�(�oBg���/�\����7���gMA	6�;q�T� GJ�_�kl�V?�f��"�[�ìu4���:���O4��0�C����t�Z�VM��ub`/�Z_�<���͑��M�uۈ{ ��0U�����J_w�l��>Ø�5o�s�$�5+���d*��/�hb��b?�y�,H ��,�i�%�S�M�z�u��N86�1�p6[ik4�Q+Gr�*`# ��ď�DGL��7��o�$�@E��Y�EkIG�e�[q�U]!WZR,�R��k@X���$,�7����V�/Tm��?޿&�<�_�pk�7!��EQkQfF��J�i����N��Y��?� CdK1SA�ѵO�[��*�זĴA+|U���s�j�19㖷ԶL�9�Gd%���83<	 Є����v��\EZ	^P���K�ǲ$t=����VO�с�1}ѧӦ��Yg_p�ܦ��x�@��#�2���fR"����v�\,2s�> �m��er���v��X �}����f����[%g���V�3�C�k+q�<!��_^��]���F��qt��ȿ�b��w��f�W���ɗ=U1聄��=���	lݷ�R�>f��#D�:���4���+����%��a. �n��
����~g˝U�	P�λ���aAl�!�xF�e$r�����,���e��Cמ#q�U(k2�4�]�|23���d���x�k�kI��v��+�|;�S�Fqܢ�!,���AL�!�|@M�����ۓS��b���k�����İ�mI��[�����a�M���y��oz���?Fho��l��JU������+:��͂���v���_hO��
.�(R>`+�h+�y��}��+-�t�`��h��^o�,��G���_}�l�$���x�����y�y��S��F[�:���XѰ^�z�L�B8=��m�VGO�j���{8o4h�a$R�}%�;d�n�
S 8Q��@�J������z�5)��{�������X���x����Y�Y��I�IA���d�z��
MNUN���
^H������j��gp�+ogu�4ȣ�OЙ�i;Z8�lZ����L �N7��<B���؍��X*���fk+�a+>�:�����0`��"��)aO�|�v{���P,d�Y������
"+�Vd��
0v{��.�f�DG��7�����-[�~����;�y����c���������i��]B2h�'Z�����Ч��bK%�vh����5�(�@y#����_�F�u}��G���bi�P�\Am*����_�%���&��_K�K�UU~�j��Q1��p��A�r�����V��Ym�	��+h���X.�-/4�B���"eK���X�[�������$��eg�w���}_�c4�(ց��p��
�e?�xW�:��ͪ��c�Q�l	/m�'�կe�� �d����E����vAv�3O��`s���ڮ�AR��3��"X*d�L#�aS�ڕHY�݆O�ǯ~v`����<D�7�;�b0_�j:�)/C�ܥ9j�������<�cAz����ŬIu���m�=ø��������:�;Qb'�c�&�_�=����{S�p���-�"�FY���Z������硥��� �Jrn��ɏ��eu'T4Z\1�4�k�\O�fMD�x� �7	ڥW.���;eo�e�Z䇛n����4R�]�=�X_YڝRuf�,>��a!�)�;:�2�5�-�-���9P�)uݨjX:ՍO0z�y>��JQ1�4�e�����ڑ7x��U������yK].+͔�2���%`H��H��q�RφW�$j@U��@F��6�:H�.������%s��5�J��h|SJ$��9�qc�+�T����5Գ7j%ʆ���G��XL�Y�k�������?t,\�,Ze2���{`�)�t}�[�
��.�U�kU�i��0!��¥�q��%��C�i���r��o�o��� �޻��^@��^�E�1��@���-.�-���Rz�w�r�t}�`����cw�rv_��3��5if���j�|������|m2���緂t{��Ρ���z��X����p�K0QC��G/�d&�&�����Ɇ�h.3f@������N�[�%�(ň;��ze!�̤�R�@9�}�9T�xY�B�i'27���͐[�j+��:�Lcu{³U4S�U��팄BKbE��o�T�L��t��c��4�t�@I�� �f�`N�J�"�~��w�f.����3?��2��x|3ؤ2�^�2��K���r�eB�x$�:��V�k':E)��r��gυ�&d���y�^ٲ$}�S@�:%K&�E<��X����V�-�,�J�!�'�Q���4�t�^��[sJ%��("�����k���>�a�-��	�`��P.]�WU��(�&G"�XP(�I�k"�INBD�V����i�rܐ�NI���M�4B֪�Y�f� �)Q��ѳ$��c�^Yeݚ:�y������n?n؛z�����mf�D�U�q�`a��Q�Z�ȣ/.��NSgU�]� e�m�9��>�K@P~��b������Ռ)E%(2G��9�QfiX�s.�N��S:>�+%6��m�N�GI`�{�(a�����d�̓X���1���&SH���e@V�4�z��S�a����.���C�}��]v/�CT��f�%��a��zN)M:JHqz=п� ;�^5�a��7����Ҧ|f��8CR9��E��s�v.]W
�ӕ��x�'F?�%��,$��>�;�â������Ɩd5���12I���;'rKT��`��a��8:i� �-�����RP�z�P�CT��T%T�������$V�E2\���Ww�|<G"b�6��@̦��T�e�8�S����#~�[����D���NdEo�l""�pVq{Y�.�5I������hJ9�n:��э�QJ����6�| ���!I8���9��@�AH��[�P��B>·B�&�}����x
��f��:�]�F��OH�����u�j����>�x�`��G(�;f��f�~u��c��)z���R�b�E���<�~��!���k�f��/�;`E̠�V�� �>P4�#�ud��ӕ�@/�5
s�9Td�?�Ee=���H��]����dU|�LSv8�v4��x;Yv�F��/LO����BB.�H�\�$S�j!s�jZt$X�6��'v-d&�t�f?Ph�"�q�G�T��h��0C7��o(�ky�Z��x�?��,¶�,M\�lq������� � ��W=$� ����zs�F�W�=�#nj�UA*t�9@��=���r�r
�,�/o|�p���o;d�z�߈V�O9=y�|�E[�����o��
#�^�����;���"�ÉX[gV3��L���RT'���B�'n
�f2�*v'�<qpF=���O)G�W��Ur�z4������#�b�X�?,ٌ0��(�/W[F��U�%�?]h׾ ��aUx$�����2�xըa�ʲKJmv"w�7�ؕm�W�AyU�գ�����E�n�V��ٗ_w����b�
��`JM_�5Z!m�=�\�����o)o|q�5"� ���`�"�-�O ��ޮޥ5췐/�D�k����_���^mr�:C�T" ����|L_�r"�~�)�HV�S|�?�;��ʛ1yz��kړ/$>Sh�v�N�o�����e��N���̘S�jYm�W���yT&Y�\23ם����"k�q�An�~7zնß�:F�d� Hǝ�=�X�VΔm�1�V��QJ���V�={�<�t�ɾ~S@���^�e5�p���L��M�;���&�xZ��B�Lb���������#�B�_KW����MN/��|�
�'��������b�8�J����3�#���3CX����}&�9���E�8��3�)J�a��.x kp���i�q�,��	��x$Rޛ��$�Z�k�e(�n=��|W� �L'�I�K����ʬ˖���j�j�j����g_Cr������N����vW��2�jn|��;�+�Dc��x��9Ia�f��8�I��hz`���^U�]��(X
������m�#���i=y0s3_�.�dy������V��c8}0[�b9e�㙙���[�yV���vn��Ta���uj��#@A���\BЖT�n�B�8;�Il��5�vWI�ySd6,M�ͤ�[��u�m#j�K����1n1@���.���ϔ����}s3!0v�FL�:o��WMT��L���3�>�`�:�,���fd��J�i�4|��;%nJ/�j~��x!M*Ǔ��ۀ�=�A�uj�/���Ѿ�����Т�J�0�?ixg�X�h�	��2�I���G���l�b�}A�f7�k���J��T){=8ϰ�����(|᧏qD��.�/i��:z^�V���C�=W��P�$���w�}9��y�m�v������}��GYD����*�V�s>��������O1�6�F��VZ1����=u�u����7[�9�t~��l�s1����`�\��[B �YwO�]�/�L=8�{=f���n�����t��ڂ�۵H+F=����.r�
~�Kl~@�{���sps�]��Y@�/f�Z��3���%�o�ҔWPO��9)g8������$F���Q��Y��|�ܤ1�� ���n��d��Xm�`h�:(	��9j֑����j �����],�zÓT��s����$S���p%�G0h�v�j���ܲtJY�Қ���]~�d�jv�9�b�A��N��yT��c�).��.1\�^��u��S�:�N�vC0��فX�5�T���*��~,�y�\:OcO5��K��q��TnZ8^k3�8u�b������"#/Y#����}w<�K�B�3�� �&9�n3_Q�6Ni�6��ʌ�F�����xd ��\ѥT�tMʖ���_<�W�uֲ� M̕����������s��O�6����0V>�������H���c�%k� ���su���$��ͼ���C�*�r+������!:��L%:s��Ck���e)C[ع��L�ڶNn.�zS���_żR��D7�G��`���b�]�wE /"��H��&�=�HG V����GK��	E���v"Y���@���}`RU���Xh�Lu���(7B:4��&�����+:Aee!C�g1%9b�X�qL}��v��=�~��0^@6H�Z&H�/k:��axQ����A�ip�ʭ�e�ьg9�x��ܕxEG�(�}��`\���2�4W[���'��ю��D���2:d��uR~�7��)�}�e���N��VPFu�)U��<	R�\E&V�Q\Grec.G-���
��m-�ܜ�Z��H7 P��XTr���S6�q�H�SH&�W#XJ����?F��G��_'�E�\t<�S��Vtt'�7��Cy�a�Jq�
�������������[��o��ֺC"[�i
K�h�Cx��A���O�v?��m��ܰR��LZ��r��y�����>���Pw�5:�?"��^�D�L�M��EВ�r�يA;\������J�n�o��[����we��Ӗ��k�{��L8V1N�]]}E�U�_L�m�ٶn�,�f���!bY�tx׽�������S ��������j����0��Uh7�C���g��,��In��? ��h} �[=�
����.οp�7��x�0J���:q�K��'b�Ĭ�]�S�X@Uw��ooF�E��Ջ��P墙Y5�d�8�5����Q�߁eg�H4�`@褯��^�,��D+t�.���լ���#-Ezt�B��TZ(GH��M3+Tn��#C)�[6���!xB�Qu���nd���3��v�Voo�XC�n��<�sS�w8�ze�K�*�>��j��k[D�>� ���~��욻��L}�q�[{�V��M������yPSk�Y.p�3F�*�c��(�t��r8���U�+�h�%ײQ�T�~x�Gq홚E�q*��F��x�a��D"D~�u�$����0��k���0%�q��r�thڧ�t~�G�_u��ȳ-�In�c���*���+J�)�dO�j�T�s!"L�I�J��g����z�o
�T��A�|��x FG$k�ݐ��Np��hh��W鐯`>u��
��J9��.GN:k	����ƨ|�'�������`J+�v�Q@/.�n���a�+��@.�sV�2��ǲy(N�r�퀱�*��X�&�����#��Kj*�#r��)o�[1��?��� �c�]Q8��+t�ʧ��\@�my^�<�0�8���޼{A�!D�.�N��[��tS::�|�����;!LrR�F���5�)��9�}���7�s�>?�~�c�{Rڅ8����S�����\0��Ii�T��s5���5��3��*0B �"�!�|nթ��U���4�~/3R8�xG��/��V�ww��r�3?Q܇5:Z��Abt�u�@4T���G���k RhǨ�aݾ����S;����e!��d
�ad��j�����`��.Ϸ\	�uH$���:��l��7[���<�li���o��-6��Q�����Ȏy4�F��r�9�N�V��Y 
�[`J�/��tNDl[�`QAq�j�߳kȋ�tJX��h � ���y�&Y�كh�'Y/�7$�����w��%����5�u_�Q{s��������ֻ�1L!�M�U�t֒>�B�m��C�)r�aD��1Wݠ��-(C��${��m�kp�����sP��%��`E�]�y����QC�l &p���Y�q�5�jR�c"�[����s�~�
eഫ�;!�P��eW�GFZ;�.p�2V3��i�JET�h
��,���*���������b�Q��ϧL@~]��	���Q����k����1}����,��ή��j�WL��=�aa��Y����sL����pY��H�H�X~���;�E�%��t6h��}/a�)��a����k!O"�g<p��>�d�־�mWn��>�(<"R6����� �a����M;4=@?���m4��W�lZK3"����nR�L/bv���&nc����r?�p�z�N�E�~^�������YzbH�@�n!K�"b���T\l�D�â��/E`Ό�;�Z�D>��I"�n�7:��'�"��eE�
��:�R(9G��@���b|nM�8�� �YP@S][0����ز���M��:#6<���+b2�4��LD�Ne�)߱5.K�iX���O�@M��>�+A�a�w0]�}�]����p4Q�+���R�o�_����j9O+$<�����9@����G��n�Y$
�g��Q��0�{����l�mu�)P|�W|<�ψ�-�[!
���<[�±�6���_��Jֶ��S���tNat���q˧��P����H�\�B1)����̹���#o���N��9���}J�rڌ0U��3��mDi�@ǧ�z�;���UC�{'�)/�-�W������:�j+�8dS�"�B��:�-Íf4b�T�7،r�9ٌ+ʉ�[6I��6[kH�]�����o��XٳP2j��(%�cs�hx�.����Ⱦ�a�U�v��aEQnYq!��b�/�����8Z6�}G�Ҹ�J���Erw��ر�]6��U���+X����bz���T��,z�%�@e��B$�]�S���C�p1�[�=b�K�%>��l�"�]�w��-5	=e���r�kyeų�-�D[|�,d�k��*c���~uw=�c9z ��ϩ	��5�l.ό�Y%:��� s��j�$ڵ���Ȫ4���SO�A����I�i��89A�`�]����U4(�S�b�t,v�Jj+�2�_��i�[鏇�Wp�B�ܣ�D��.M뎾�ẑ}O�V�f$��{�;�[�#�+��{�F�e�h�Q�us�0�=&�9n�P�"��e�����$�86�gɮ�s-}���q!l��@j�F�.�-�xl�v�W��O����C�Ȩ�fU9�-�>dA�� ��O��<'�c��SG���1u["�!�sM�kc�`����NZM�ǭ�>D�⏏�V�ЈҐ�妕|=b����6F+H�-�C���E,Ä�+�1%Pn�Ͼ,���.  �ꗆ����*�<�-���IKx@_����ǧ���w)5�cE/>���p.7H#{�x�/�}�M�&�^�ʻ. �'��n���?�D�B1���%$dk)�l!r�R ���oÞf^�y!�&!�Od��KB�Ϙ�����<����/k�����	�����f�vC��)�!����#�J�i��nm;�B���3F$�� 8C��,�F
67w���-~�w̑�M������U�*����ُa��b�Q� &u�Iv$��E�=ER���Hl9�h���΁գ����sn��P���v��Iǋ#���pLl^;F~��\^*�#I��v�me��ii�q[���gQ[6����K��FP�<h���-��Y��2��n%�"N� x[��L� -��*���#q��b}��r�z�*���ZwC�P_��m��ʧ�MKo��8ɫ�S�(��~�奠��n����3 �� X�dI	�r�s^�u����֗��s#ruі�۫2�8�v�����w���%���\4�	�+�Ti^� n�]9�3��e�[��}�=�R���ϺQ|�w��ߕW�\����Voҁ��^#��xl���_�}8QzrTR<&X5BS�f��V*� ��T-�$��;D4�%BYV\�~瓖��ӑd�&?����)��hQ��۷��������O�������XPx��(��T0G��:����ڃ�Y�P��0�Rg�,�5;��³t*>i�q�� d%i�-A���i@\�r��]�R�����:u�)DK(@ݱD����A#[XRN�ovCW��Ɠq�[9AeŸ�ǟn����㎌6b(΁��l�{�g�nq0�-D����p��pز�7*�s��2���}�j���#������jpvî/�ŗ�^t%�U��Í�c�������WmP/�8T���H��'Wx��b����DܥzEh��f_�Q�4��Ƈ5w�z�l%��s�v]�X��D|ԃ�jۭY���d����Hv��JwLp�_�"M���iK�Z����x$���>��`БK����^��2�����˃�L�ʠ�j���A���iH���W�)��
r:&��x�#��"�OQ������HqJ�������;�uZݺ�� h�RI~кUWEM+4�v�JO�h�����Ec�?�K�wr����[�ݑǜѿ�
9��	:�������H�(�i|�O�ͽD�G�I��6Q!�8��K&,X|����Ǝ'�J���*£Ѵ��̮��L���BO{����@g�������'���XL'��6SpZ�)���RmmdГ����t9�[Z������!5=����N��D���"�բBy�.��"�|����GDXj��ƈ���2�4�5�.�Rf����6�.~�{|mΰ�F$�ܘ����g��t�}��N�~�	2�L�;��Y�,�-km����}&�,����l#��L���;���4l\$X�Պ��C�2dܚ�I�iJ�)�p B������דC0�4�i��h����8b�l�o��z��тI����WiD��lu���B�����!TW}X�Do�Ɵ8�P�3��s!�d����5����.pr�B)0�)s�o��]8׎��3�q�_�fk�TEפ�& �Zd�,�|��R�����_:j����Ds�~�v ���d��\)�$�S��V"�������B��o�\��Y��ip�V����0��J~���t�G���"+}���N�c�����
rZ�в�΋p�\��s�D�2Vq�cUBfޙ���\�����" �ƹ��y��r̆Y��w WLgO��6��T�� D*.u-�62d��d��l�K-CGÅ?;�����5hk7co�C�1O�+MQN;��B%+�(mL&ס9X�z�dxqG��<h�?��������!�oy�̽ԿN"���8F��hT'�IP��qq���E����C����`�1���df�<<���� �Ѓ$<���|q�*�����T ���� װ��v���\��#���tN��yY:(�������j�)eE�8�h��ϰ��4�����OO~c,\:R�u����(,(�rZ�;��HZ��TS��x��(=����'�12����GB�j$y��@z.�Cw���/l�E�F���gI�O� e���i�d��ʨ�-�B�	���_H(�9F]��a�_��׎��Mx,��Q?�"Nn� ���'/3⾓D��
��m���V����2���:`�5�"}�A�\,�C;6����U).7���p֊	l����~�h6!��=|;�������s+�Bg�\�t�����%UA���u�mՈy���s�}ɍ�`n2Z����W�U*Ar�-5�./vp�Y��mb'6l�����
|�����J'I�@��"�������]IT�5��B��P#Q�`R���~��jI[OS�������x�II�/κ��63RG���$�M`�t�'�Ȳy=�t!����nRb��
��%t�1��D������<�~RQ�ֹ�!�r`G�B��0��빗:0E7����?����~G*8�݌�0`�5l�0���K���&i�ct���|5���u^ά�Bx���Ys�ԕ���0�<��jV���=���u�$�����k�2�A��*�T�����I�e�����Y=���l��;GT�-~L!j㚽\�蚮d��YC���$�^(qd�+[!@z.-B��m��B4S���}��W���2�\ӊNMM`���|�N��y9,���>�ϑￃqg����<Հ�7�T��gA�X�����1s�����#�����܈"��܇���`
�m��`���c�<��+�y��}v���(�Gf1��G�Y��Lp0�3B(	a�̼�����|U�~�t��q$Phq$[��y�Gh��+�l�5�_��������y6\t% ��;�R�:Wm�W
B~b�l�#Gx^@m���'�f���G@���`�d���0~�4��č|�Ӳ�m�A0��y���f�Q��Y��X8���Z�Qgc't��ݨ����VD�����f��
̀/M1?乗ɷ�<Lz N=L�:��S����V������z/����u�N�P��sQ[����v!���>w��D�gʀ���Q`�EU�Tu"���=1��P_1֢���>Y��\z�5}���Y��Ǡ��Ǘz�k̫"������J0�]&�J��C��ƭln�F�
��:�B&�4
5�51��f��mК>+h:H:V1?�4��;��ג� ^t���z͆B8�r��-Nk����[p�k�H���Zd��<�HP��v���!h��/S���6O�Kn-p�ӼH��j^�v0M�u��������2�0?S�G`�Ҏ1��J�?�R�]�7�V�+{��Yݔ�^Z�!(9ooS�)�ӆ�֣�����U�"g��A�2�[t�7�;@�[�Oh�
�}c�XKw�M��hK���
���P�6�Δ�a��q�yIA�y��PDQ�H�cۣ�$,�����;�` ��UFG]9���v9��ʌ�Lϭ�-�������T��˅yd��)n���ʆ��w�	ӓ��~M�u��9����9z)���-)��F������B��`@�o�]���oI`�3M��?Lɚ�ۉOkJN�|��n]X�g|�LW�l�\y�as�2�E��-�M0��`;�&ߟ��8z���1)�t�E��ĥ���� Q��M$�B��F{�ݮb*�� ZL]h5f`�Vɝ"G�T/˂�D�y ���<��)�q`���l�J���4���'/�ԍ�zN�F�*
B�Dh.���~�����R���,�A���覊�.Uc��R/0,0��'���#]�KLd��({1~�2n����S�ɯwX�6:u�]�`�N��CJ�ӛ�4O��(��7�%���z�3�b|��,����z�U�|�n��]��Л�KCyN�ZBh�TE��:�D�a/�D�%|�~׾Q\9���ޤ��Z�ڇfHwXW˞�{����j��ˌf�R
װX�"&���Ԝ,Q�lzDi^7ȧ�L[;��G���\������ ���[��Ҁ�C�P}kL��$0y�`��n
��q�����H��ti2	��Ȟ28��Õ��X��̩6�{^���H�w�!��xĝ>���%�=��st�2��Å��D]:ޏ*4{V/A�;ɚ�5��~7ؤ<?x�NY�s^=�W���?V�T�t],�f�
����$dk[/�m�L֊�oN�r�	Z�0VmY,�n���J�o5�K M.]�CV�8�Q��������U2�V5�дA$���f��J��:&��q����@Z
'K����`��*������+3��d 5܂e��ɛ��kpǟ���n�y��8C�_�W�=��}S��Qnf��&��	F
�a3�n�|��<MJ���i����U�s���0 �jy�,`?����񋅥@U
>�F����Wn2�tƄ�bX�D�%l��X~J��h️0`wB3��X�H)�y9#�P��Du^W&f
��unR���ү�o�\'xr;o�?�����0�h�oI�	ӡd�âS��D����6�e&��e���1Ϗo�{�z7<��\�6{N4�Ѭ1E�W��y��F���՛�
rX�PSБ����g�F�%9��Q��7�e��FY7����ŀ_8j$5+q��`M'#YK8w+]�YM��h��)w��t��A8%]��NTP2�,֘��g�Ki��Q�
�q��Oh�C�gM��C��^,����pD���\S�!ݸ�����(����y�U�b��I�ύ 7�a-�E��W�kY�XpC-\,�/�ܐ;�N�^qF���Mf��3N$�L�f�fރ�a�&������7@G���R���Yű N	��)�`k�RE��	}�DCj�ܧ�MDǘ���C���'���곂��/�w���vq�[����6q��D�!�0��m�b���)��xЮά�������"���s�eG$�[�ZeC�4���m���6�Y)���$:���Q�o#Z�׊���|��}�*��i���<�F��������D�-{s��%���B��<$4���<�{83p�i�,#�o�y6�D��5/�l��wI�}?5g�>�ѳ�O���r�>C�b��J���k�/�G3/6�~�aYrɜ�N�	jRTг��hk��.I܁�o��$A|�ŖG9n+�x�q�+c�?��Q�EE5v�@����Ŷ��u����֨��.FJ#W���t�>���_�q\Ā�
lI����*%�-������2H|E��S��HU�r;��s>VdG���>�<.2�-�b�ɫ�]8� ��,��Q�JC��&��q6���ь4l���� ������|�:��#u��������s�]L�Yp�`!t �{�j��ntr�Y>��:	FI����#���Q��ι�Z�R�N�}���f�{�XK�#���绹��J_v1L��/�$ʟ�o|)���*G�	���[sq#B7Wb����;>�ZGtSV�zR�FȺ�nx{�ɭ�%��߱��:���*�b^H�p�Gf�
FB1��L�Cj3���4C�W�{��t�ԟ�R-5�s�sA�����׆�}�}��;}�����_��9h�h��c�B(�����`d��"`
Ծ؈_��Mtf��߫,��`}a�d��"��:[�Gȸi��C�qnKY��GO�_�)�5�I����j<�� ���H6�J�s�t��:!�v�P`�1��\�"��/&�8}qq��j��sa��I�iw�����g�h�֨)��|#�'8V��}���C��|�Ӗ�U�]���ۓQ{5�]�w��k����1����;��f�C��V��F�+�g�b ��U@�I*������Z6J�v��EEt���Zz0*u����Y�P�V]<h�q������<�Yxa_v,(��Gu;*[���&��;�R��h�?+����8h]}��Qr촄��
IO�p1��մ��IS�sa��+�)�G��H[P�����I�Ō�)+������8�����w��<��i�o��
i�,7�k����'96�b����=��!"�ύ>%D������V�A����x��F�\�O�ՙ�?�iCGo�<��}�@eyĪu(��
PZ��@._YO^�GNKF삤�I)D}}��t�e�F��&��D'ި �rڢ)�+>�n7��&�;}>�C=�{ێ���*VXdr7�4�Ңq���]Gu�_�D�j�6����*������~V�i7�5J�v�2���ݽ?r��{$n9F>�ɸ2���0W������MƟ�S��C�A�D2�q�!^L��L�1�))��W{d�t�-\�t��E�I����:�����(��,�|#�W��u�����G݋`�SC��^��0_=xql&��\�����p
Z�ʖ�©��"D)��+Ev�d����f�C�/���I�WCw��eJ��`�Vp�2��m�@�'��/�6 >�$ <@l���G�!C;?jH=f��;^p	(�c��/9�?K3FP�tK
ӂ3��lĄd���Q�����:)�$o�|E7:�O��v1��k�:��yE�����_8�B���Ŵ&�Ώ�C$���l�o$"�n.���<�]�t���bX$%��_7_�I�f?G&A3W0fN������p��8eua�qԃd�c"KJ�+�����%�
[6�~WeNN�"�d=��v��
���r!qE
�Ny���]H&��W ������Ȍ��<UnBC<2G�gv�p,��^$G?�����L)��m؄�&p��\�<m! �iw�T�	�s�T���k`�N����mg��Sr@z�JS�DI��Ƴ�����.�]L3ݹ�ؽ<�кj����5���kV�XL��L�:�7?�o,��D�v�V�B�`z����\a�\�Vo�6aq�=��X�_���c4tS���cB/��)qgyAGLG0}��n��	��H-_����z~b�W@Z.e���K�|��j��=mI-�\�0�WK��8�V	��k7�V�b��m0�"j��U���4 I����5� ���v�2NK�yL�NMoпy�٢�������oQ����>9~J��,/Y�o3���۟GX��t�٢��J��Ŝ�jQ4F3�h�襈��Q]%cu�-jp�u�,�X�QHi�.����������J��oMs \�w�6��ΐx�]j)�]�+j��>��c=�!%�!y���j\�p;f'�@ �W+yw���'��P*�0J��[�1�jA�<Q��u�Pz��!ui+�G�|�#��ީ��!��NK�Z�׼]w,�9����I�l�6,��x�����w~u��/��=��J&B8�;�����	SV�*�'�^������&@=�+8��׸�_�߄���إlAI���t���7�;3��A��:w�(����t��V+�2��1H�#��i���OB��	X�GF��	�>9����x��Cﾌ������aH�÷ Gǐ�u�<�4�9v����s�[���`4�ʀ�u�x
����)��l�b���*��SMߡ��L3�WJ/4E��2��M���?�{�_��lyBe�Շv�{�L�;W��` -܌h	��J���՘�#���^�z��<,�$ i)��V��s �KͰ�`v� ��R�*'$<��%�~��z:��4|�p3�����C��!%z9v;�����9{������:
@���GCyj�kuL��`��Md'�zXgǮY��G�vN��v��*�a�uF�а�F:�;ڞ�Dh���pi\b]K�]KX��DG�qbR�,؎�(I7�A�N��hV�]�Ap��0ڦw�a]!���b����%���~���XQ�2���	���]�)�)5�$M8��L�e����!� Q�zz���C��נ�_|6	*9�u\��,#�����v�*n���0x�b���'���|H8f�-����N���_����5�pLUX���g��@�l�@Y�/��>�>��*�T�59 � �ay?��-�. w�8�*ɵr/ϫ�c�����V�q)ػ��k �I̱⨷�-'��0m�F���D���mJ��x��(���<Gw�)�/�Tj�UyR�j���-������Ͼ(J0c��/�_c�t���(�u�4)c�^�%-N�SI������9�{�,�{O� D�O4W�Acf�T�S{����T��XV}�(����r�c��lՙv5��SY�&Mj!��#&�������Yb��'({H`�k/s���Ia��/�<u�~r�G����t ,�~]!]���勢Ɛ�1�p��#)������Oe|�w&�(��U�b�m3O��s�?_Q��L����i<Z�f�����%�@~�Ƒ�GeY:�;0s�#����Ԏ�����>�����5c"5
�����6ᇆ�آ�G��& 5��I�g�Ca~�:�~�OŠ
[.���uRB�Qs��k@�ZxP��JPPn>��u����l�Z=@І�W7zY��h�57���կb��	R��ǿr5��xx��g�S�~2�-���<p�����G	����{KB6�ޗ��{�োE{����U��X��:���h������ _�,���O�2��{M���`$=����&�i$���>@"�e��<�͡���"��
sm�<��P�~|��Qǌ�y`↴I�5�s�S�ƫ��镴K��Dıa`�� Y���e�豑��q�K��v5+�z1Ncid�"���)�7�S�#b(�4ʆ���כZu\E��FX8`��H��š�/D�ȎV� ��i"q�WfY��E]4��N��/���Ϟ� &ز��M&_x�.�x�f]|�>� �,�?��pIj��؄�c8�8e�Դ���>�g{��ǜ̈́�(���y��x!���V�4��U�:2�n��ζ�EU��P�ux�kOw�@��.l���4{C�ȗ�~{a)!�@e]M���I�j�#'����h��`���?g�F�	�����V��J���Cp�b��i%�#46sg���� Y#�� ���Og�6lÖ�������e��c8]���cs6C���j��1>�[k��%R��U"�w��A9��w�Tz��o�Q"ѧM��̂|����xHG+�?يE��`����=kdj[��\_����R<����ꈝ��a�iM	���9F�h�����'bB�a ���1d��6���9]�"�!���6��R ��+Bw�u��J�`aird���K4]��I�;�!����6p��z�}�����?�ŋ��.�*�$�QVHo̷�.]m�v�{�B:ׯ!b��cd�y��)�.�o�*�{q����C����{&r�;�9�s�;!�aE�er�]C6��`��%Q�+��Y8�ct�A=�ſc�[�`�[]��Nm���.�3�tD��Zٛ���, �������5���1�] �<�?c&wd\�㖡��CFu��褑�o��\��D'��>WwS�͏�v/�/��C�&x&�ۯ� T<1�tq�~�R�]�_C��2�ܨ<X,�D�L	�5/W��d��[��TB��]�ił�8�>�P�d���yXc�o%�o{'�o�C1��<+����?�6���釷�J��ۉ��f���L�8f�K�ŭ�����E�0@��)��RnM�]�u�2����������|MY������� &����L�I��  �Ѓz�t8���Ѯ���*�>�M˔�J��ľY��eR��*H���R�<����O���߬��\����%K'��|�~)ù�e�W0q>��I�#�b� n�wE�� 69�M��K/# �B�m�"�>:@aL9�(�����9�����V��cR���MK5�[�1ϯs;k^ge��4R��N��L���)V��;0v	뎜V��4�la�_!��'x��9A�%�L(�֒#Myb����oB��xr��wMR��X�
�q�2�r���>��#�����R�U�H�W�\�6c�sE�!�TYw���v�UxXu:`�49+S������R1�D����yv"�p�n��	�����u���3?A�\e�/S�cDIuT"SWrGz@�N�o�:IV���<�1B�^�)�[�p���2���u
՞��y�"�)xہ�#�=���͵�!}��������z*a�X�qNX�g�4�*5�c��/c1���c��G��/�s�Z�s���dߙˇQ��՛��GQQ��
v�6[η<����1t����Mq��-T��k0��Ԇ>�&3D�5��٣Ҩd�Z�#b��|w�Ѿ�G�#S5wE��;:yL���o+�'Q�|֔glND�2�0�\�{MS�R,W��o�:����"Z�̯x��סּ����ΩLܺ(G!e��.N�_�>��B����n��T�6�Vs��;x$&���a1d9�J�t_���ٙ:-�qT4�<���$����Le��F�ޗ����s�Í?AvJZ�G��-f/�VtK�&���!I�{L��������o����;��r�_�h��^#���O�ͬf���f�Z���=��ȲO
"[����,g��D��X���<;1�:3MPc�������Zp�l8�PwH
��*]�����NW�E`��1@�wd�$І��$ZG?�)�/��#��Pq���w��&?Dr��
������j�l-=��G�vI05i��W��W+�����p�BA��wð4�O�FʴR���Ta
�/��Y�Br5$�I�
�0V�<%�)g�a�ß�v��(��9`4�����9&Lt����Y;U��12�E����4�2Pƀ�+� �h��wl�e�BA1CyŠ��v�5E��2k�7�-<�
b�K_�_�l�<;��H�$Ӎm�A��;���"����@�A�_��9��fI�|(L�9����K�*�e��_@���%�W�&��b�sܧ0m��Ȅp����O].Q�d�.�t�~;f�E�h��Տ��@z���S;Q
�j;����c+9�U��5�W�b������< �����U���:D�I߀�s���
!�F�,�[Mŝ�����`��E!���n-�+��ʟ��z���=��r업J�=���9�s&���0�S��/g�hp�פF]�R��,���S��	�-���+���w��V���KG�g"��/V卑���e*��ē��[�v�qQ5�

W�U�;$qw1�e��?"�F�{f��jQ�x1z$�������֎u=[iֹl�*�`�I9�d��PRb��_�v�~���@�V`��f0^�����G}5�챷'S�_M�l�˙H8�o1�����֩�×޷
Y��=(�.^��B>���zX!u��y=ԋx���CG\�����Q�{�`د�x�?lI��hـx%��G
�1x���fOnԫ*ݱC��S��Eܕ�	�E�Rl�{^�|���D����Z[}B�bfQ�:��gǠ�mPf[�Vҩ���;��T��oT�����I��T�P�]�r{r^\���0�}NT��,>P�� �0q!�AI�d�Q�W��⒠V��M�Jc�;��Ny��>k���8}���/u3�����\�~|b1lG4�����eX���'SU/��[EF^ˤ�,j�"����p�k�;�D����K�!�����L|�%B I{=a�Ǉ�Or~/�s��U�7�ɒ�#�st�K/�;�f`h��n���sc0���*8׉��i�&��`��u7/��4�����V�j��4��z�{�Ù��Ձ��%�h��4�����9�o��%gN�꤂��D�L�I(�"h�˙�������X.M&:�E.̷�Y�k�?R
Y�Svq��	�Vepr+N�2u/�(s�*�h�Co#�_��j� )�Y�]#U��`1�@��i�5B��
��!ɦFY8h)n��8"���i*��r\\~��\>�#��=���04hѿ�0y�U�e��9ۃ�����ͅ&tB��ʞh`٪��|Ҟ��lu��1@&��tQ,��&AX!��{[��8]� ���&	1ϩ�q��.� C��`s#݌O��x����~1;^�;�P���g�f�� �Nf�m�6c?���7��]�>	�W�Λ�7mk�P�(ZP�h(�}�n%����_N�$U��_G��m��7I�y�a���K�O>`���	�8��|� �m��b+B\Om�W�:��Ί� X�+�$=�ʩ�z�-Ck����I��s4�@}�U�t���(��XG$�:�pP$���6
Y9���r��8��CyD_D��o�%���7й�xT��*��ǘ�R2��������G���,��`<1*
i�GEV�`�D�[қ����wW*��{��FC�=e�t����w٢>%�}�p
�~O˵w#�҉^�Xr��� �-� 7��L���ɬ�b{3hZG�~ kꡩ�[JH���:�����Q��yE�v7"5�қN��&���!���59���34:p���&�CX�48E�˹&���k���{?N��{{8=�qZn5*a6��6U�=�����vߢ���dgruf*��q^��pIv�) ����Ʒ\*KCg���܄�vA6�*SJ`7�S�x#�G|biO6��dN��:a�ߦ-μ�V��L�ۀ�	ɍ�^����θ����m�|;����8�(����7(��5T����D*��᭽�fⷽ@��rʪ��	$^Zt&������qZ�k���F�c �ػ�ȃ�U��`2㲺�:7P(��r�2���\�|�هt���@|�� �6�-�u�5�^�������0��?����6��/�q�$w��΃껽J5V�<���/���6�܋��;A϶ĭ�^����B�Ȑa~� {����
��ǎp��r
��Ͱ͹5؋�/���:�3�����B)���������Y�n?oZ�|de5����u��!��f�w���s7�|y��⛦���zR�P���/��Qc��m��p$c���x�lM��o-�>�����+�[����AA�D12l`��S�賴����i��� �m���J�Ϸ�.�I��F�/h`��;ʎlq��HY֓�p����3	�L���	�+���JX���3DX�s���e��5���r7���$_�$�%����}��sZR���@[��7{=&��,HN�g�6#�C�!�0���Sv1�/~�-6�X�1gќ~)�t�_W����~����5k�hȴ�P�ȏ{qU=9�$�3�*�B�ܶp��Dtr�$S�_�U�n��fr81;r��:�X%�d�enP�#������.�Sϖ_n0b䃃F�E���.�a�`E����M6�l!��\&5�ՙV#qu\*�	���w>��<��\�k�N�ב��E[@E>
=̉�)`�~c����*�A�,��س����4�e>P�r�3���k%��z�UD��W[s(;2K�*E��r�͚�>���cߪ;���70rƟu�`ֶ�3��E@$���D�}��Fu�W����-5K�51�8�V>��\�Ո$�E-n呣�wd���E���}�ڎ���3y��e�����_�?�@+�s5d��I�v6��6:�z��tϵz/Ea���8
��kc(����8�r>����HKE��B�0pzE �����=N��?�ڤ��9\UheLW/��{�`��@]�G�1��n�+Z����
�XU��e��},���jMx�S'���H�FGGǥ4)���NG��Łj��4g����K*s�Z'�N�Y?iҾ����J�	��̢��`�ίp����p�(y��4"���%ҍ�o�o�)$��7�i��#�m��"��td��p��{:�n�̣ך����P�R��:o$)q7�@�G�d\}k����� ;��()���ҧ����1K�2ԛ͸3)�y�� %�њ�C��e)h7�{���{�ëq*�h�&˒T�����#<}��#giI_;��
�$ <[���?W1,=06P��b��mؾ¾�L��L�JW�o���}_�#�߅�*9<�ț��Zrg�I;+�VL���<Qׯ@��9�%3�̾qн�z`�6Z�K��� ��c�����m��4�?��W9���כ�d,��hv9�-_>�ϯ��v	�c�`l@�C1����
}�E����exY����5>E�=p0�da(�S���4��"�!hf�;-�r���c�R�)�3Y'�i"w�Y>ݬ���ê�B{�"ΉMO��R�if��krNǅM�h/������e����)���ٳ7�m�c�=�h]r��!���shCk�7���7��`�q��̑!G�e��fv5Z��S+,1�$�h��&(o��<�Pk�{gSv�5_=���Vv�x�|/.c���{u�ui�>x3p�����z��FE6jW��8"�'�~d1���C��eur��FN�a�i����"� 2�X[��Y�rO���C-�T���j���1��
��,�g��T2�8�#�AD/������"*�p����VK���9�3 cqV�2��g��ے��أ9�z?��6��r��A}@�(�(K[@�B�K�J�
�	��nkpa�5&�p��)����J�=����/��[�ε}%�uI��J��Ȳ�ڐY�Y�2䎀Օ��r̈́��V�~��Q��F��W7J�a9 ��0�������{��R�~f��%q=S*
�"�"ώBl���GB�;��:g#"}��j։6�J
EOÕ`��% &?<�#�%��� �D	�:z��E��HUȺ�A+�!_N�;���(-�/@�6i�Nr�����ˡ�n�v�Kv }���ZR���r/�Xi�*��b��2k���^T=	���@�)�9�58�!W�iW��w�X��@|��	���Q�r���������=>�u��S�F��V �mC���F��~�2'����X���`�[����sC�=Dw\E�8��a�$ǻ��V ��=��"�A�L��7�vk[�{C�?��93��o�ck= y
�v>ݽ�H,�Zt�'��5����|Amu�V�p��W�n�d�D�ϫ����ɀ.�?II+�!�j�����9!�y�7�YA��L��So�C��2x�X|sE����Zo&|/:l�>��S�r��97_�����)P�@	bBwn��K��]�V��A��)��R'��4��%3z�S��ڏl:���{�i�
�2j�S�-s��"�a��A��c�!pGF�oD c��(�׭5��ҷ�T\kGQ/�y����xӭ�f��8K0�$`�e�<("��	��+ۢ�N�@���B�����\1M�W���e�'o�HF�6���c��1��K1��4~���
p�J�����)��k�%~�<�����y.�6.?K1�Ϩ����s�>���s�kf����ho�B]R��C0�-��L���m΅ꬫY��{�F�!3ŋ�Nu����:��E�����G��ܿ����әI� ��f�5륲IWO��z�v��0�Uq��o-�ԫ!��`r�b�X�-��ø���&�
�C����ze#h����h"`���
P�MVM[�um"�zN�L��o����˵z�u�cNw����S"zm��]���(+��B���6xe�i�RD���(#�~X�%��do���Y�05�*;k�o�g�t�L�vq��N3t�}� (��K����Ms�ئ�!U����т�-��J��X��Kwȶ{��	^��,S(� Ǆ�Y��u�HSL�<�?2p.0�>�Tt�(��=��R`�n�dop_����-�hP"�s$e!����0�N�e����wعOX�aP�p�Gb�b�G�u��Q�`{��3���~S?�޿��S&}個���g�[��ZI��[>�F_D̯��Ng���9��sP�����Ϛ2�w�-��ff�s?��=�����8g�j�q�)��/���V�Dތg�6m:V]J��Ɵ��UAf0ņ|3hK�I�����䛒���u+���2>�!Z݈ ��� ���4�x���-�6z�8�otdO��)����rP��-v���\#�}b�um����F��P �s:�e�i!��AȊ�v5t�o]^Q�f���R#p|Wȅ��2ص�������͈$�fU��3�3T7���05�w��J������圱8�x��]4$*��7�Å�����=���*XA)o��.��/�c�cR�	�
�3��-g�?�ͤ��0�"�Aˣ�fm��Uu�B�P���m���g�4O[[�1��S��],o���ҵ#�~��'���cB��U�- I�7�݀��|g��5ʠp�'+\�+_��g�@UBY�[��]���9;>�^����[��6!^}�p����NN?��,������D����Ew|����Ƶ�`2V.C0[��ZC��4����-���8GbQ���m��f���:��/�S����FǮ�W�%���c�GK1<(yd�� ���N~9�m���n�.��_������{���O�y���TG�$���_inE��q�ɋ�0���P��t���N�ԗ��A�V�{ʕ0�.�
f�ȇ��)<��hhբ�]6�{�a��V������{ő�O����F�@72ܾ��i��r)�t���"Eq��vr��u�$�˽�H&�d�<�}�e�3 �#j�/5���R1qc�Jm���56�#/��R�ǿ~�[�s'6�U8T�ޘU�����e�+�S�%i�q���+�_�^�X�ѻ_��\DS�Cw��U7�ޖ`mo������ß��q����y���Z�t�r��O"�j���z���-���daz�p����Oem�����K�a�����u�ߔ$x{K�-,ս��NJQMq� �|��="T����ئ��G��B����i=��τ�l���m�'o�Fͅ)La`�N�a�������L�I���M^�ťٱ�	 �$0b������3�N �92�g�@�����`g��jZo���ӲQVjc��e�8�g�OW�@d��s(��%w���p�ӹ&t�8Q�Sm���.o����Өn�`Y��?�7Q�UZLxY�~f#t$t�O[�C��{O$��#2-�C�< ʯ?����� ����I5*ܕMkwu�M�6�x\����-"sn�<=?{�5F!7X�#M�v�߃E�� ��r.�vo^�#�ћ�2��g��i�=�vRuU�W����?�p�1��O�z4D�G�Rf��%��)���R�>%h��qt��\� �l灁���>>�]I�>kb�����jn����Zn��~���Vб�@K���J�z���
f1T�~�d�İo��,_�Mަ|�ƘFKl�K�>����M��2Z������?��Z6�:j�4d��w6p]x��c�\�&�/{A>�>l2l�R�`��+:�O��)�#�&.�8��a�M���e�S/�"���L]���m���ڕS���몞��
���Pe��͈�_x''3b�vj�g��X��i�(��u瓑�0��}�FО�ф������L��H���7�M���r��SWI��B��Y�s����~, �ˎH�y���H�Nt�bW�h����;*;["�Jr��>�8�Cc��A޾1}P�At�"VӼ��<�ѽ�l�W=��g*�c���HN_5�F��U(q�X#�t)����4q$(}�yZx_�~�I��Ї ��\��c@;Seq��$���'�h��x�"���VMc�]��;�W�)���Ѣ��S��Ц�*2JR�p��	��x���o�Mո��PL�';�
�8^��`�}0���mO��n�"�\�=��g�P��xv�}a�& �zZc{c+&?m���i��ۭ�(�Lw-,&����^����3�1�zX-��0��I5���&Ā�SKu&?�YU,�O�ݞK�VN5i����m�ۤG}~�#�|�;�����J�^�݋��R\��b`[5AfH};y��5=(�Nt�ޣ~���t���B��m�}F��%0o��#����]'1���geS����ZȲ�?� ]NJZ�s�v��Y����*�#�]�3�T?I���ߓy���7_�����{;E����L+[��.f(��A��ΰ�5+��6�ە#M�����_~_�yIg�oe��6�WM��39��������m��F�,�o��ѷ����`p�-�a>j��'1���b1(:F��<��2�?�|OF@���NFb�E�+���̅��00����Y�O�Z��+������ �a����7I!ϪAPa�,� ��V����gBI���Z��ɖ����yP�Q��3�B�0�@��X�ꩂ,<�T�\ F"��T�H��3�ZS��CQ{�*�!�Sp+�'/,i1;x-�w����:�IU+T����F�1�7G��)M�v-k�d$`>��M5�
��hZu�L�����]���b�~�	��� ��o�[��!
��U�{�ҕ`��AA�plFD0�Z�;Iz��G�<kIL��oLӓϭހ��p�6\;PR�j�zu!���9!a��uj:	�����O���c�H"� ����s1�/�&��yA��5��]����I��s���aj`�����2�	�&�7Lv-�|Yb?܄h&_w�mp"PҙJ/S��'by�Z�S#�������4���pu�g��$�/lrB���̓d����Z����W��z�q�c`�7�b�=b��{���z��(G#i���ϲ��r���N��X�rYv�c�	#|oӅ�����#Y�>�{�;Ӂ�Ë��32��@K�1\ �3_�<�4u�d֬��Y���Ds��+�U4�/�����#���tځ����e0��쨾�+��\��Y�b]n-J�uz����
!<��ag�W|z�x��279����~�S�#P���<���
b���N�T!$Ol/F����tP�H��P�n��p
gY�Ât�����<Hy���b�)r]�f����r����H�!l�j�������NN>O�3�{=�A6w�C��A�E04L��9Ef��{Jkz��d� 츢��on���Ȩ��y�n���7��!ßLeP��*{��=(}SEi�mH���@y揋�5��p���8,��61A�����'y��/��XHł��>t��R65�j����E���d,4�R8뮱;"��ʘd�n~����s];��~���~c9������
ЈD5-�=<�8H(2���H��w������G��J�V�oI����C��w���H��4���zI5���p�^�A^�ƪY�yWƥ���sD�[n��Ҽ���+��B3[���S��N�7��1jAuY�w����*ŝ�o+M��D72!��dSB���.��WPʸ�$�u��Ψlm���`�=���C)r�n����@�Gx�2���˫����h������]��G(\Q�B���U:��O�i�H���m���,�(\��b�h��D@,���-'(�މ�V{b
�Y.������;�s��(^�"ޙ^��>��k�p�����`Gկx�(5ٶa��䛊ZL#��B8	�j�>h��zm��51	:6[$i��t�xfcC������M>Nڨ���K��$���R�9F��%���QBAq�C.�c�"��la�]��!w���4vP�oΗ�Q�2t��C�iO	 ���jIA
�V-��>�JC0I�4���E��[��!LSb��K�j�WQ"t��P�ޅ��|-o���P�E%:�pw~�)���Gkx��⪟#���	��G9$��u
%^���5)$C�:�]&J�ye�8ۊ�
WK�'-O�7c�nDA谁�9~y�|�[Av(W�����`�l3ȈQ�e�P�Z#�������6���T��w����,e�@�����N�������mتF�*s�N}+���a
��'�b|�����N�yg�M�m�t홻�4���_�93�8�6M�G���$"~�~��i�	Զt}�W�o��\���KzV�b	�mX����B�i=��n#�[�)e��7��=���^�R�q�d�����ï\��/I֦R��=�bQ3Z��LЪœ�A��7hW��3��0����El����^gE�c֫���qI�C��Rq�_�p{�b��T�A8��(u��G���X�c�0Q+��t#��#��=�1:td/:�lc��Fk:U����<|Y�R���D%>���h30w�jB$'�P����6,H���gkV6@�XH�<�*�)�Y&V[��r��W��:>h�x�~J/pMjdE�fKlK���'ط�g�[f��c���Ye�Fc��9��l,��T_mY[��!vi 8�=$���,�P�k	.������KC�Ɛ����A��@0�H@�C�n�fZ�^��#4EԈT�Q�y��4 �/�:�	v�[U<�%�,%q-��g��y���?�W7U��"��H�͓�-�F�f���(�: � 9�O*����x!Fz�2L� �%�w���:�{巴F�՛���3L�w����g)��v��ZY�l"Q#I��g�B���"��
7'��z쨼mK��g�d��)�n�M��A+�CkWS7l����2���t[3wܓ��-�����|Q_N'7��m���^/�&������a|L57��7�CĽ���!?��B#��P� h��$��U�y0� ��D��`ɧ��I�	6�?���g�$0����#FQ�w�gO3B����⚦��q�$a��v��7��͵�V�������l�7(q}����SҶ+of}���}B�-nݎq���_9�'�W.�%�\E��#(�3�������m��&Cc�vN]`�O?͊�ʾ���oԨ=O8�ECւ��+����j�i�&A hZ�� Y_j��&�8��(rrU�r����-M������� ��3��������:E��tH^�kD�QZ9 �:�ue����ˁK���."jA7��t`. ml5��}s�Uy0h�	(-э�,�V+?#�W"4+����s�I@|�8���BX�Ǎ|���"�1}_LX�@�v������M��'"�X�đ:�ʶ�;�-����-)��J:��Qջ�֞z�);ߡq���~��27^Ֆ���+��=�Cޛ�j"!>�V�=G ٤�X B��P�{�7��>V<���/obK��?p
�¥S�2��T��3mJ�_3R�gg���֏Ս.�B�������r`����r�q%M��y3Q1
�gcL,sx��C��bK�¹��A�_��t���2Q�BR$�>k���?��㰕 ��/�O7�w)��	��Yt� K�|X��)-]@��6#�0 �+�M��/�qn?B��
-�^�}�:|�J,W*���0�S�e	nd*y\�郜�X�勏�eM(s�1�.}��0��25�iJi�O�r��p��V4�&$ۿ���u^rBG�W��=v=��wk��-c����c`R` [���~���ǌ_0l���&��kƷ����j�Kt-%�����s�~&OD~�	�r�i� �������޸v�/��O���&�O�'Ǝ�ܜ�����06R
���&N�q�	�v�<>�Y�:��٘B�9U 
U����L%ܞm��WM��G��b��k:}��g&B4t"N/�`��Ի��7���tG�>�X8�R�A�ap�K y�#��9L����N%߬Y2<�N�sq�[�|U�F����˘7j\<�"�t��݉I�2�w�#��7l&�u����fsn�.�5@:"�����0w��8�&�犑Y(�.q�;0��\�%L*vM��딗�4�̴W ��z��-�ʿ��Ωe���܎��AoԂ!/�[K>b�1�|�Y�-�]��r2y9����6T<�=��wL]�oϫz�smO�Atuڞ�ٵ3Cnt�>~���E�a/=���L�H�����<V�0� �ud�}���K"�i� H`ǭ�V��4��J��1���E����0�Ty���7�۰��96u;)�����Q�u60��4%��S��"a��V޺c��2����dþ����}S����J��]�Y8/�㊪�O�D�ȹ�����+�P��D-.�kd�٢`�ML�z���E��.��ǁ�^T;� Y
EiAI��mf��G�i���?��A��
���T�TG3�W�(흹a���z�M�M�?��^)�����I�eo�-� �6��B_3pw��1A�O�5�ك(ٳ����x4�$~�k ���1��Z���`[mo,�n[����x:��_M����<�&)��pYo�c�ߔ��-��	��6xMfz2Fʣ���Gɑ<��Dˬ�z����&�qD������5��]v��!1#�FO����⊻���w6��ɆǛ%���y6Y�;&����,	�W#n~��ؖn /�Ǫ}H��)���o�?J���MŊ{�U�N�9�w�%������,�9�k��s�ѩ��l�gz���\F{�Wt*��m��}�$Ǚ.�$W5���,�A��?}7]0f�R(��A
���Z�gH�D�	?J�����CLِ�4�$���=�U��ˏE��w���g*�XE_ߠ�Ʉc_��.��+{�v���tt�xȉ�V�u��M�'�rI�9��� lf�Txҷ��ni���>�3�#L��0VA ��].��Xσ�x)O�,&կ���kvU�jQq��ΰ-?fD�n��:]?p(�E�W�R+nr%��w�7�@����V�!�Sf�ɉ�RR ���j����oWĵ*P)yV��!�]����U��w�^9�!r��d��H���(m{�\4T�}�F���-���n�u�� \L"h�4	���;#��/���Ȉ`�ۃ&,"y��X�Ez�ko��o��X	k��0qv�S�"F=�,x�5�����Z+����eO�\��oʄM(D��C�}u�P��a���5f��o��������;?
80�|:�/���7&c�^e{��8W ��.#�e�  ϵө�;�a�i�������c֌�Mu�"��(�}�p�s��S��8�Q��!H�~E"3ҩAJ%{CGΌ#�ҟ�9��=$^"�'">��H�����7B6S���S�_�<.�GΙ���]�-'|��^Z �V�5=�H�3�r�K��n�]1� w�����]�Vˡq�k�^��9+�S
z\q�迕��@�����#���蹻�u�k�5>�٧!���K�Q� .-���H�:p.|	�g��I��	�Z~y�h�m*H�K�5��V�1d��ʆAiC@0���1��D�q�|p��p���u�5=U�[e
ecڴ�<���O��Q�LeI]����vz־��>'�M���1Ch5�4����z�_.{Ƴe���2��3�Vu�GY��E����w�;D���\
��!2S^޺�z��	E�A�7��b��5g�k�0"u����랟�[��������?�o /���,�z��}f�Х`�� �U�����d�d(�UB�ͯhG��������<m�$������%�Y����0��s|���0��Ʈ�1y����H&��ZYO^�w��1�&����X���7���5is���w�6�ɬ`T�٢IRY�����a�[.Q�{lP`7}�2����b^X�ܖ§Z��%�X
p�(�M�|���Ϲ��h$fx4��GZ��m4�I?W/(1㌍��l/�x]�'��s;7W��[�LS�8r��S�{�;Ѳ�	D*����'���I� ��R<<IG`�N*��}*�}��<u��1�$5�5���`|)H�Y�vz���N���$������ǺW���i��5��\�yO�n~(J����sS�~Ɔ!�X-�
�ȵ>�)�Mn[��$z@l��R����+��&�����sl{��]��X��XP�� kM�o��q�Q������
�qU[ďgP�-����-x�f\�eY8�;�SD��X�B8p�f�J�#?�٠m�+�D��ө��+n�n{������3�B�iȶ�lC#���y��T=a_����[���]N��g@J3>��F�0]�k�8�!.�&ׄӋG߈��Z坹���n�7�v�xD�AsFF��Y�$�]M�e�Rqi�D+���v�g���T8��:�W{�Zr�^���6D����JMcF�m�o�Hh���(W1E/*s;��@�c�-�H���4(�RcT��+��c�ZV0����������C���T|���į��N��c
~j��@;�Q����C�����������O�R�5"`jnJ=]�z�^�
���N�yR����'fL��+��A/Y^���y͞s\�Yi�E#�\}>1��c�X0=[:�� �fe����ky�7)4y2��S��.g�j٧+8$"r�8��H��w��Xf�u7�zcl%�b�{Z��I�=|4(�jJ�A$���Q���ZD�U��K��4�z�	��G���ކ�гnvH��u�Z�Y�	,�7�d�~�[c�33/y ��H���h8�ƥܕ���w��(��/TB��D���Y5����n�kX��(�'u(L#�X�O$��B�� �g��؊�((�tG6js+��%�~�;	�yҧ~�QU����&@t�g����/q&Jz�A��mK��zBZ�(�!�����it`��ު	�E�ĳ�����{nK�#	8.�q�S\e�C�.��w ���I�	zf��/J�yYe�Z)�jv��T24iQ`[쬦gt�����Z�:aj��~�]����7�bxP� ?4��3���S����V��<i�0]�=1�".w(�Hh	�כ��H�%GO��;t��!�`6�6n?�]�<z�@���o��!�y%
֞{gx�յ���&���k2���D����0�2K�u	�~��Pf�a�U^5-��?g �b/�_�l3O��*���K'CANx@��:�H
�u-w���� ����.��q{�
%�솤)t�h�| Ib�;T��o�1l������*t��+�~�)`�㵻����Q!���|g���ʼᵨ�%�s���̻�^D"���ۢɿ��]��q�Be�+;<��0���3w欳A̍1�l�	�<�8��#@?��C(��!�M4t�Nh{�C��1X���1p�*��+�ή�oyZ~�V����Aޫ �h�BɵZYN�9��ψ�Q�����ɍk\�/����e@�z9̞z�4-��l�n��j�G�j
`Z�0�􀪈a���7,�{2d��`�0A��7�d��ظ�ңmT�9��I/�������?�ȅ��~�{�܁�!��՛O����������9o�l��iy��$��*�uخd���9�rd6�L�� b�w"���Y�H�D���pA�N-ߝ9�"�-���4 8a�j������g�]#���9��cu�p�qRߝ.�m@��iḺ��i��t�V�4���M�LGo�䯄ݫ��Et�K䫀��#Ux����������,�оH~L�����C�uo�|��r8z�ӭ.ܵ���2�Z;ζ�������~9,�T����u�%T~GM񮕷W����X!N8�X
��Kvh�t���d0����l�β�c���\	�K����)���Hb����UZ`s쉋�QYo�]�p�fD���'{��1�R��)$����n܀�2찋�]��+�ʅ�q�G�k݉��X�Z���g�A-�Z�u�Pd�xtx)�'�N�le1Z����^���z?��!H�f��l_��z�|�Gv���eG��C�GH���؋ϳ��n���Y��L���ꀠ��ȃ�E\_?'�#�ۖz�A� $�8Z?|�b���.���zH46���)���89p�N�H/��y��R��e^�:���(��˶�7�e�V��6�I�������M�kWQ�烌~��_3�	P2*s����n�>�ء6�Ѽ�1e�ʗ����좀L����g7*���D�RC/S?'��(lH��YLR�P�s[^VCn�TQ#������gNk5f�ރ��g(1g��0eo��-r�gSi�n��^�Pē�s��ܝ岐Ub���5�e4s�RâS�	8^ɾ�nv�1�!p��.pU�}�ߟ쩰=rc�e*�S�;�.������΂�ӎ�خ��'�O�T��mRW��.���9�{29ރ�V#@�Ь�̍����1��r/q]���ZRq�Onn��(��c!��'�(�pT�;�u���l�����k�!���f�e�/��t�����^!?5�5.��ӻ^c���T��e�9��-4��v�c�2�[6�G�{$���FYE�\��B����w��Q�C^�f��p�)#���O�G2AOe`F���mu�ʣ
��b��:s�Ӄ�UcQ�a�wyJ�]oj��ԝ_-��܄@^&��G�J)�^�:��#\Q�t�j��Kzv�]g�n�����	�3�� )�׉6fxK��#q�>פ����
��WQcIM�}�����x UnE�%����.��N���ĿJ�|z�r�����!�.�����*�<��7β�"���[N?�L�:q�a.M�S���V�sqR:�pF�/�@#�x��,3*'jg���X�Rj� l5]kק�U��F�ª����@�@���SM[o�{N��m��,��&��F��t�4#�w���A*���`��| h\`_�t��?�L�7MZ�I�62?^+��)U M��嫖$�+@�d=�']��bc�`w�P�R����8,C*0��[6�f�fG{d�m��݅�!Y�j�D��*��s?!�c�(�Vব�c@���m��S2:n�j')G�=*A&��B ���"O�-j�+��w�^���O)&�؟�tg�m���e� �D&H�����Q�2�7R�d�T�F-��ʢ��T���|u�\ ��,d��ce�fWz�?M~�Z0wơf���i��>�"�k&LO���,s��H%��<��D�V����� |m�7��i���p��6Tȯ1*ɘ9���]���dP��8~���g�h
]�>s�0V�.Q~��D�Ͻm��+�z�A�!�1�I�6��6~�pX�O�:a�*-�_LH,�ъQ�VRE�ok(��F�k5	\.� U8�f�_{���8�D�D�A��9Mş�iP�ZۇFܜ�|�٦�{lk���ZM�Q�Iצ��;]���R��w��{FE��UH��]Ⓧ�Yp O�z�Ii���d?��y�۸M�8�#�v��+���ϵ�Xe*��HK����R'�j�>���b��u��*��#,,|8��&��R�������|�Z��Y��7���>LZ�&~Ķ������Y���GV&��eO�H~���2�����K�n~�� %8�(�mJ�HqH�HU�7�LI�f\���_Y�X�}�ʩM�Y�1�_�_.=A�sX��z��uA���E �����%nڪ;|LGf���?�5�7������^��S�&�C5���:$7ނ��&���(�R��5�}�~�?��됖h�̡����^h)����*$���p������ǔK��X��
6��0��빸u��'	|E�ݼ�ź����_S_���nQ���K<��a��W����Mi��x�����L�8�5P�����i�3~��&���`!U-9#��{��ܵ�	��/&�����u�8�g��\I�\������y�ߤ���	��Tѯ]���(�~�kJw�LTmƌ��+� ���me�L~��e���Ý��B��v�������9��<v-�+ĺ�Rd��b�T�!�D���m�4c&��I+ى*���E}�&�H�A��&U.گ��L�b3�sµB��#������{�&V�Q���k>H<�5��:@O�#���;���"�xe�j�9����6�p�S��d:�&�Q���5U��ܶ�����ՅՋ`Ds+�,���S�D�Ѱ�j q�>��ޗ�ut�,�^ڞ��!�M^{���o��vH�8w�3�1K�u���/Cpn
<�D�(_�߆��`GN�=W��ƾIӔ����]�9�P��� N3� g�?�dt`��Є����+F!�o)�X����p��ap�0ކ�u�jA3<�%4�𸌐Hz�+"�,�͕�e#T�k�,yC.�`?�~i� �r�Ve� �� �`�}OaES  2BY��B�M'��oƵ*n~��H~�R�K�a�,tW9����a֐��bo�<'�G�-`,�Dw�))v6!�iع���Ώ�L���1�#�F��pS����$;��R�P�I�˳�Xe����|�ic��m�QSm�,h��4uK>D ���P�	�B+�E���-ϯ��hLK#��&:�f<�2���E�B�	h�Ӣf�T�݋��'�FՓ�ܶ��<�A���#�+�yE��;0�0��z�(H��Lr& WD�/��^@�Fٯ� �\�Fڥ��eo�oh��B�lTܩ��%4Z\^˪B�k�~Z�t���m6�S�����㽐)0v��~a��le��>i�?
"�n�$�]���oP�9ꋴWp���%��U[+���~���
�E�qm��*T1 o��iNY햨�������]��i�1c� ���v�~Ep��J��Y��⟰�eت8D#XĂ7
��P���6q"-��Zp�9vu�K�	*����ѷ���]d��5.G��7�LA������L��j�����[�����DB����5\�}���`�k�LW�x%��*O���5�(p2uwo��G��9$ako���Ҵ�,Nu���N���+rI���� ��DU����⺜�.��m>ic8�{*���w ��ATS(-P/j���\��ݱp�,��Ȧ�c��mY�A-�ޣ�t*�|��b��:`��~6(��?A3�F�Qar���c�=�%�R%�N:��z����i�HĪ��[\#��%�>0/����a��;6��^��a�J�f�(�*������6�et�C�6h>b��k��kh��x*��Qr[eYVN�Z�~;P�G\��y\$f2���ȏH�s|��+0m�m���P�@�o�e�!6��r���K�@tqF�d:���T=E1���A���Ґ��f��D^�d��9X����&��r�[8�䥶dJ��I	��9r�U�0���v�#��#�'ܲ␤fs4KC���,��
�K�{�Vʃ�����<���uM�%�a��ۀ�Qi��|�4�(�q��,}���?sq%�fH�M
�����Ⴇ���=BřZ��M����4Ќ�"i�+��bz�#x?(
B"��}�d�H3�����Z1���c���A���HT�"�:�H�-"mv"�ƞ��u���E�ho�U�i�J����O�ut��DW�����G4bB����@���%"UUan�i�@˖�)��C�>`�S�)����{EA1m����qW��t��$�1�)�M�e�N�]҃ͺ��y��訬}�r��-�OO�F-�.A]A�(�ϻ�.4Á	��w�b�gwE�|<�}��Q}c���#+V��#����u�o�۸�Ճ\��2� ���	� -���o� �/qp���$\�r[��l��M���&Lvm�xK_5�,6��W��?�^��υ�]NK�<���BK�LY�h��"{��A��t�h�y�3��1aP �ѧ��v�������e&��m�:��G���*�s�S�jO��A�3���}#���b�������P�NG�t��3h����q'E�&l��; �e��B���m�-���Ei䭿���[l��W> ��}�r�0|���)p�w%#��r�\w�醷{�S�Еƭa!�V1�.r��+��Qa��{ljC���._&��ˌI��75�����FD��23�.�F�蔀�p�uV����<ޕ!?F�W�
I�-ǀs%�X���O5U�r���ϣ��j�МP=����W>,����ZNP��'WƲy��q�op=|(�u7"��W��>�Z�3�Y�s�o;[N�G�3�C��l���7�L~�?ԧ�9V�.x[CgSu��w#lc{nG}6�5±F�c�az�&Y���D�>��U$��IS �dΛ�R>-$�ߺ�jn�ɺ��e�o������7�b��x`���sS?p�{Ƙ�Ѥr���lc�K8���D6Z�O^1�d�H�.�T�VR�p�i���C�5�������,��m�k�����	TƢ�F��%���q���t�#�G˂9 �@@�$��]�'o�H����'�-�?���}�(޻�⋀JG�)5�o�o��uo�0���U�De\l(e�|���äח3�lHBjD?|���u�i�m�4	ө�VV�8'�31	���i�&l%�0��9}�
��T;˭;K��7�/*m ���������^}�rCy0}K���$O?`��Xܶ����"Y5���aj��`骯�e�LUt�A��E� f+5U���]�vsy��8�7����D3�G���x�o��k�C�|�$���8���;t�s+#�'|�u�!���&�7)h�l��@�{ju����m.�1�o)'��mt�<sU=#Jk���Mĵ}.��c��s��ńv'�2�>I�INj�&�Pw�ב)��A�X�"z*��SCZ�y���N���~��#v{�m;1�w�0.�� �1�7�YH�Ν3f54�Rpɋ��#��%Պ�4���ގ��%�~*�~��.f��7B �ޓ	�y��QY>x X�����r׼����t3ȍ%o�����y��������mE>���"EI�ڿ|A�b,�er,o4�q���h��J�s��k3q�e��.��L�#y�
��$\@����}��`��?a�ɢy��C����
:-%ea�R����I�nN���(����I��V�m���0u�&f�z�9�#߇!��u��7ڏ�G��\b��В���
,ջ �-� �0����eK�NN�A�إ�o�"2�V�a�s�$O��G,��?�����!�&JG|�z�m<\۔����X��<�p�?��]�k�|~ށd�M&p�� {
)TJ,��syoG�M��]l:�N����-L��1E.��$ 3��6��?
�����A�<�e��,��U������9��z�>�F��!,&sǭ���l9�1{���<b'H��C���˄G�eZg��$�恅��;��Q�/�YYd�O�YQ;�*���oa$��8kiG�d񿺲ѓ��]��<�/|D,h�g=yc��j�Xb�*����R'�1���p��D�;�1��7{����|$���})^��맑�dN�D$�׊!l�(�1�||ZNg�di�BH��⏵+��4Ȼ�X�0W��ΰ��
�C0�d���@�0J�+��[�d�}��b��׎�Ż�D��x��g�4WN��hd��O�P�ě�(�����)sY;�D�d��5�ju|���#a�π��q���p��2)"K�)`7�v`]�D{gԹ����8���CO�T1Dt���Og�o�H�'?�� s�1����`��?�wX���6; NP2����5�r�{��g�# �7xz��oXn��Z{�I�ק��Ѭ��U�5�p���!�f��o2-���F�#���d�� �Ʒa���1ߌ�3s��0��OC����׈�x�+2�51S���Ui�H�Zӯ�H���:��DA�_푺�3�����0��:"��~ô��%G%���V=v�T���L�RM�����&��"�J��'�U�g�?��ߜG��$�k9sT�Uk(�M��mJ�:�k�y��~){�聬�����Ȕg_� ��R?�S����"��� �_�C��w��/������:D}ݢt0
;Uy:a��8Hl�X�:�X;��� ��`D	��z`ɢ�Gi=�L�:AO�z�>��TbY67_�j7(�C��ϔ����=Q@�i�h��KA0�DW��^��;A��i"E�8$S��[B���EՋ�`ك̵�R�2��;(���
�āow�����n�'���A#>�(�f� �4�/��V�p��j���nF�m��Hx���X�V�h�>�2�y���9v���<�B)Q�z�?�Wl�Q���;�4c&b�~2G]�3~�nսXWZȎ���㾣E(���(�R��w�k�ֈ�9�HO���7D���M�7�.`�E�8Lۤ^�y��y��娛�թ�W�tqwqƓ.{gv��h�I�..9PE��C���S��e+���&u�G�U�'���)��7�"j6Й�!	h�<	{�BT��;��>3����Oc%}@Y^��@�#���\?��{X9�A��c,��������ȿSO����R�zngC��;���a�Py
�/+�4���Ӻ$�L�	�hg�4��U�Ģ�3��7�R�s�Ki�>`��υ��`2�S ����i폺�E�ė�;W�-#SP��OF��,_V�'@Ym�k�!k����!Uq;����h�gd�����x�#B������XIi @ťځ��#%��e-s�3�K��W3�D����.`ݣ�词iH25�F�D1�����:�m�~^���
DH�K���1�ϖ��.
���'��g	��%b�_P���C��w��$�n�ڎ�Ǎ��P�
��[���)	�K(n��˲���$R���`����^�I�G�#4q��ä�C�`^��P�ZĴ:,��H���\IyN2��(ilDd��i<֟��V3�Se�I
��)����!�z=�m(���#����9"��N�3^@q@���ܔ�w� �uP�:��ĸ��q��ճx0�3�l�K
�sH�&N�ΐm��j]�/r^��EM���or���� �|���� ��Qebl���S���Y���u��G8�s,�O^�� ba�k����\s{��og�M9'bo��W��Z�ht�7�����jy��BNb�=o7.4�\J�nنT�ي�`���w_ ����G&Ђ5	�����l�0P��U���*tw�_�y�Z�x����"�>�p}���3�N�S�Eb8h�� /�`�u
A�~�4�:�!U�?�����%}���@6_�q�q�n���i�(�����>}Au�,%�$[�=J������WE��t�T�g\`��O�Ԯ_<`*n0*�(X!�!����d�x�����&~g/z�B�c�5(*�O�&4�4́�rY�-��^�[u{�j��2��,҄[p�R�Aq�х��b��e���Ӎ6e�j/m�Do�#F	{�w
ѵ�H�6YG���U����B����Y��Y�e�#ܾ��2N���»EG�eo���D8�])�_$G/IYu�Cʲ�GZ��K��ɠ�e��;�v��-`gW��ϑ3���,���}G
��W+p��͜JJ��y��?*yʞk	_H*o�������=����t��qْ���c�Q��Vs��#`������]���F�vOC�>�銊-���k����3r��y�g�x7�Ze>0�C(ף�Wl�~�>��[�[�(���2��4i��ԋ��(�����+F:��.e�M?<���S6�N �_��$��7���O�Z��J����ho�UR��G�+��Ah���Y�y�=B$>n�#�|���0��e-pT6i����CJ#VVL��g�קx+�z���ϊ���\v�~~�2x���IU
��Fk�~��Iv�`�.qI��}�[��-Z�Z]|��
��Y��b�[ X�^լ�s��a����,�,M����"�����6�i��
�o����_����hg��th��\��/�ј��i1��X��j�-�����N8�_[Yq�Ё�O����6�ި	s�Wm����U>��5G�v��K�堨��7���o�/'+�ảrUZ��W������ڭ^�V%�@)R�bA�ܔU��Ey��ͪd��7<�Qd�Ӿ3�pg-�/y>3g���@�]:�S	�ˠ�t$6��zpZb�
��ՋZµ+�T�c����.U FTZ�gM����`s��3�����y��,�N��r������g�������)Ft�U�@ȟ��[r�ꙛ�?d���M�*1�C�4
������Ki=hb�䉾{����SnTe����f �I*���������܉�t\��X%E�A#ml���T�H4���������?D��}Џ>s>ls%t�C�u�GN�*0�?<�E���М�J�#�z�Z�3�H����2k���&P;C��_��%�<$pin��1:㣑���|.A��=�._q��]$y�(�A���9�0��@����R��rB�2�o;od5�~gk[���%��x{L�s��"D��6�RBgMn�S�{!����|0aFEk�G�V
��o-��q:��������r��*H{����(-iH�t��jأ@_m�v,��[h7$\
sƍ`cDS�����N~ɴa5�v��]Q��"����.�OK������V���
H�&�Y?�a�����]E䘂.A�˥�1O�C�H�"G6w�g�|�G7<����=M��+��J��6[�-��7��r؀�_�ą��/h0o���Tk�x��
���B�O�g�<�W���v���)vTN?�(K��?�����r���� \]�A�DY�B[˷��Pt��w<o�<����ḾH�w!e8D�}�p�3^�����T�̺ٜB�_2�䶽�_a�}~�	�!~�Z<�E��µ��6/ቸ�>� �T,�n+>d�v��7�"KUA�e�Z����O��?'�*z�߬��9r_G����(��>�+J���`:Jv/:g�b�����W��z�L�6,GUZ�@�a����>� ��i2�E�)iit��ΜEUTxp�O�>_̎}G�dg}�"=���Bz@����\2^x�e(������*��Jc5��1j%k���cO��=_�y�͏��P����h*U��[)B��r�h�[-\��4�c^<���.�A��S[�����������f�˲|�n��ӫ��k0��3���}L�[y"��3S'v���jJ���0Ç��Ә@� {���uCJa� �HVW������ Y�c�,$��`
D��#�r�M'�Cf褗�h��띥����.�ګc1 ��B|]��"_���q�����[$\�o�*>1�R���Y�1�}�[�?����pj١�m��]�⣙�9&����L==/ѿ���[��q;����G!�D=�-�b�:Zx\b0H>5�늖�>m����^�,��*�L�>�r.�E�N4�����"Q�Y����өQK�o��)�XR}��.����H���P�����r5a�y+�FI��]
2[&I.��^ڈ��o,�����k7�ۏ�}�&�iq-�}�n�aBJD����܃~�5wN�u�r�ׇ�Z� �Nx��&��O�Fj��L�/�љ����~#1�X-h����!o}�(Y�]F9ω���'�t�H�B����7�u�n��6� G���撇r��@�9R��-����I]� ��� �t�r��Mj��9g�tI�Ѷ�*asL��F�RO�f;��.���^@�溶��w9��x@��B�Al	�f���%�����͍�g��@x���b�}Њ��3"�ϐ����ON���n���{e&�~%���˂͘	Sz�f�/�#]�@K5�@���Ob�X�Gi���G�D��[=-K_�{@�ꬣ�0��4N�Ƃ����r��{u��C.G��ؔ7�R�&��|��ֶ�{��ǭ,�|�5JW\ʗ�Oj�6�5��kN���u��9ߦړY^�"[V;6;�j�4�\�͒,�j�)O�7��_R��� e��!�gk�,{��
���i�� a�1��s�~�K�6]o��\z��#(���|��%��更����>�;GT:�LRdO)@U�m{}h,m���i+i��d����W
�d��o�J��J�J������Ԇ/
�c��)��a�T��
�Ry��vF��b�`�1z�|sj��ܘ�ި��~^���3���Ym	nxVc��d:��8�1!
���*u<aa��vrLt"4I���𳋣��}�Qt��:���#Є2��/������2����#���h4�寮l��2��a^$�m;�Ɵp�f-�}�r:��@��%��ʀ �oy~��}ͅ3�L	d��G��^R�~[�O��^\�Nfb���[��vYv���z�2�REal�V5�u��fh��VKrq�����D�2_�(I�hX$����� �b�͵$P�+U�����sc��̂\�ջ�J����d͝��nZqQ�[
D��K]7{�إ�t��"��u1�%����]�,<,������������p���lt�����@��� ��a��_�x!�K�>��:�H�|�w��/��h���H�N�:(ǌ!�qP�� ����7s��^mǢ����S�����w���q���SX ��N����C�#&�����+��u�p��I�7���s�o=k���t!�E�.�@p���qC��LG6H�B/k�	=���4>3��u���av�p�~\���Y���[]����v��C��R�dm�G�x�!'��n5������ŕ`��g/W ��_�Ɲ��j}�&[e��]�)�����8���D�wg2K�?�@b�(}��>�.I�����@�	[�oU�]���,��t7� �����j�:TQ&�G���,]��Z,A��� ��v�_ʳ�7�<����n	�E%��f��&��\k��YLj�wa���}q�ژ���� f�[��&�NS2�
����>��$���
�����[��|�au=�V9k����7S?�5Ec/�Oh�#^vN�0��s*�q�WG8餥���u�3]5H�!�Fo�l��l@�$�X��F'�_��9(C�m�m��]�S�9/�/�u=r8IN�>w~Ԛ�����S�����U�ޟ9���Y�y����Cq2K��;���ú�ͻe�	e���}��H�8Ei�8Ҫ�a��ɞ��Bk�������/f:xˊ�nl�cS����c.XX��;�P4jt�Z#�zS�{��j"Zz�A�2
"�0�~��:�%$��x�=V�,+t�T��aVS�d�Srd���r��#��I�t�>���R�c.����N��1Z��e[+8b����,�q�L�|=��Ϊ3Ր�b���N���~Y���W������H�[��j���PC񜔹�%��4�b�b���Y�������/sEr��z�۪�T��ya�̭��'�����V)'xpba��Q۱<��E%���t��y�����p�0��Ӻ���O9EU��� �k��bV�Uw�#6���(�Q"e"u}E�ҏރ4��Ϩ�O�Z/<��<��n����P?�2�*�Sf�P^��4�~y��+�����/�E��!�~��1U���4��U�8���}O��v@�Tܞ��Y#�s��V	|x� ��$[G�27+��� jU����g)���}�Е�#�pl3^s�3]\>�3��z�7��Al|ͽܪ���D���!�X$���ƕ1	P���G!��0n3���Vh�st
�,��-M����h�8�з[�>��8q��>`X��8�Ã�4W�3�u/M;aY���� ������.YO�0փ+߄(�W��n��e��m>���z�!����1�[d�&�u��� ��o��i�2��*���^��i�Y��R	d 2P�?�DW�X�ؒ�:@2AQ�+m|*F��4(8����@��ll�bFz�EIPKwh=��X;,���̥���!sp�S�P��4�~��@p=X��Zox܂�4k�l��(W��+?{J2O����ot���ʿ��N^w7�s!���~;���s�Fy�.�d�u#8���1��rd@&О+�D�r#݁�n{���f�rG��}�E;)A�ߏ���Od��T�3�ݙ��[�y��L��F�y��GP8@�21�'�ĩΊ�� 2�]�ZnkDp!I��O�%JYg� ��b�NfO�pS<$����&�Q�J[�y�{{�W�^�O�\��hW��IR�d������V���, �>�Fq|Z�l�ZBhא� 	z�ީ�Bt^������&C���(����]����l=U����~73��S��゚\�*����^P98կ�.""��G�k��Q�T�¹]���y�6��
pC8�Q��Cxɂ��.��kԇJ���Ym��=�쎢]��>K��=�Do���wp�a�w%e1���(�`�͆���	Q8Jr�`kIc Jp���B 
'�>��գa�gP����6_�����Uƍ�їQ���#���2�I��kԔ�� 5,mWK�4�;%��@#��$B_5�ihu6�Nͷ�]�G%p�L8j��
��/�Q*��ôT�R�c�v�˥��8;�����E��o�FL@�%�*���S�����\k��a��NKB.�9䦙�dě(���E�:��������]~0�/+9T�0���vb˹��c��&��)Ѱ|�>2�9P<O���0�A��o�.�d��t��@�9��=km�|>d�{R�V�m�tcQ��y�m�c�.{x�H�kQ-^yd���]ov�,f�N�����J~<�Rq#{;��y�����H����N� 趙ʪ-�0<�ˁT�m����X�$u�1�A���� ����yw����/=�[��x�����@2�l]�YOm8#L���"D�����	��u�}�b�9�M�f(3կj���37�tfF�=����䫋3Jl]��)
�"���X�����A�+��ӖP(
��/�QWu=�(���7�^Öq�{D���޾�&kr~�n��%��O��s�6ۙ�|��d��n�FtZq������ o��@ �a�|�	����"(GG���y|�h��%�ܲ�f��%:�ż9.�rB!IV�J8����/ ��*��cL�6yO�o�һ/S{�j$԰w䞕Q�נ�Iڅ��t ZӸ9�͛��u�&���C�c��{�zM�����|��#["�lVUW�������"��xl(���[p�X�DS\V�4fJG�>�)��~�(�'�dR��a�l�D�Z6|�-��ྒྷ��;���p�i�Ԋ;'��m�1�(m�G	0�y�h]z�I\�Q4�ɤt��JD#�p�oLKd�|ag5q�݄>�[�;>�ʽ��¡Pl�Xа����}1�"�&�
z2W��X5��ik�/��G�I������Z澐�\,)1p���8]���;�^ɳ;���7
/b�Е�X����p	hKx���V���
����]��DL��s�������f<�v��s�/�LU0��n�5\]C*C�>x"ֹ1;�g�4&iY�&3UF �R���������^���E��,�L�+�E�N�R$Y��<�5i��� ��gy�8�p��t��ݟ��h���V��m�pT@��\?���תa��1��;����S����n�v4"���*���zP�a��`:��Y�u� ��+�#�l*�RP���#��r��9aԽa��~�`-�!&2D<4�"� e��<<�Ax�`����IyLI�-l�;*�x"�������t��A�h�[V�����!^��(O����^�L+�9�a�C�$�
�U�ۖ�U�;mDnd���~��Ø&��z�Ӳ�ƨ����v�o���G`_��w�r|�$�j���j�qFh����G�?z�1T�Y��_Ne-]F�P{���Z����1��d
�뼉b[�(i���i�ɰ��Qv��h���!ގ�#�Q���7��E'-.p\d�����s

 �]�7�Q�iL^H���Z�`*�!�D�z5�i�W#�P"g`'��
�K��YW���Et�.!�`�ro��Zi���sʗpa�mV#�i�Cg�p�A��`Ҡ�p��
���K�lx_�F7�fwEy��sg	��	�	B�F��;.8�M�q�Z3UҶ��uc�/��� Q"B`96sМ^64��xb�����0�m��I0�j�=J^!�+��e���yy���ɧ)n��8�D�پ��jϛa��_l|]l�3���Egf��|H녀k��2*i����̄o��"����+/��Y�F�.�e���%�u�R�8yfz����Дn#���)~hM�zy��T&T�(V&:O����
p�	&-E�%�]:Κ���A�O��5�D��k~Ǒ� Kv^%�NB?Lxo���N����.Dג��~�cOE�[�k��y)G��ΌŤ��\�CW,�����~@�ߥx ��z=I��j�D����U�X/��ʷHb���-���D�Z��u��.=��
V*����F�b�/���S�u{X;��IG��~#��#�;N{ ;� >$��yi�p�������Sr}^�Bv�V���bE�ԣ�t{�we9a�v J���CP~�����1Q�� ��N�&�6��KZ��l�Exa��&�,>t>J,�\�q���l]�hPmj�M m��~3*���->_x�M��_��E9b����i{!��?��5��o��t����'�ñ�i���S��77T�B��X#���w���A���C)H��ƅ;骼` ��/I8���YC7����t��*[�`-عMn�:ֻ����k��D#�R��%\�Q;l�B�{�1�࢏��g�j&�ڝ�1s{
���f�#������㕒Uԁ�S��Vn�&�+�X�J�^��s� �SnkW0.��'�6�6�@&1�	�nC�8���&��ǉ���XH��j4G�^"U6��J.s�i-�K!ޯ@H�l�4��;{���O��3|�܈3��)�ѦѝPC�&�C����^���Hˁ�(�� �0���AQ���.�=g4�<�� �����x�4�k���"��Gn5� �Sst��B^�x�(йmc#OZ9�#��4l$`j)ՈȀ(�c�7��~���c3�v%�jA�?�v:Ci�S}�5ᠶ��#؅28���)�	�g"�߄3��US����r	4�"�)�U7�ͮB1�:1���3V5�r ����5�"ݍi	f4>3?��).2d�F�/���
r�=���R�7��T�k�x�}�� ���g���|YcأњYY� _N���znѽr��7�x�.�˂H[Y����jܐ�EQn!
;���v�����P�ha3��\�)��:����c��������Z�S����;b�ۤ�����B�?�����V2��y��v��鲹g ��ܲN��m�`���Tc�[�~w�VH7�m%��'��f��r1�.��������I�I�(	H�˶h���S��$�ܢ�I�R*��h;�
�ڲ]��C ���q]u�O���`�s��=*=~}�8�o��d[$u������X��ig����H�����tP��[^���c	]��OU���׮g9��G9��A�ppJ1ٟ-)��_q��þ��u�D�W.)������qF�i��	p�zլ��^��A�I��|y$%�[@��8p�,���Z��Q+d0�N+�W+��<��e-K�?�晃2���� �9Flvi!���'x�ZΡa���SJJ;N4[�`,/�٠��m(R�����]�f`��8�3��;�ID������5�"�I�C����6��M#Sd���/�'Ho�Z��f��w�н�l�Q�:�bK��i���K�E�r���FtV�rIěg��>Br(��a�� �3�.?�@����'��,��i��w,#�ZI"�V�|!��4�BL���̛��zj���ձL�,�hb�+�z��%Y��z�L���Y��&-Ø	x�R#���f?��K2�ѽ!�t����;͕0�� =���!ۍ����;�,��@EoG����"�Acg2{�Q���/��I1W�^�̻7"6AbT�MCwZ�TA�o:��ۡ��4�����cίC��j\s�9�-�����|�ztXK2�\��kb+��u,��^4/<Zi@h��q�xC}�d�Z����ͅ���D��|�I���hë�^��7$s"5Eß�aS��Ɩ��#�j�n:Kߠ��(V��8 9�4�^�X���d_h)p�G��n��4����bs�l<�;1<�u������%;4X1s��A+�QTܐAc��N	����#�2�"��fZ�e7�ͮ��7ݍ2����}�@c�����݌��)m��P��<b�qgdT�׹_ZQǚ�A�
��h�^b���\	��׈H��B#$y���e�i�^�=ҡ\�e1Ns�8�X��g08|��e�q�+�׻׉�M��w`���61ܹ$⠂��Y�4[�b�BZ:���9��9���q�LK�](FM$5�"�^3�u���R&����o�w�^��y~6�6��~жpRѻ,�NZ��i�X�!+���7�R(����ܴ�����b�vq����>ZԵ`�`%���dw2�#dFM��}qQ%W_C��Ҽٹ��\���C�bL?H2/U��0������#am�o?>�¡�`���\և��R3COd���%��4��B�^i����Kr���(y������а��Hz�����J�r4�&мx7�S�:�>��p%ȅ�?�,����$�+w� ��lZ���tR�כG��"a9���}�a>N��q����7�@0��f򃲵�����)*�dP|�5������{��uȽ��,���	���_��vW���Z���><z��ho���Z�i�����$�t��Sg"�ǃ&z��u>�O��M�fY��S���-��Ԣ��J7�3���7?
%��m�%6��~T������ʕ�L��$�[����(>1<-j���|���U@^'��������)ߊ�5�x�H�
1�mӚt3}�*TF�?��ôӇ���0)e�7vQ��@�瀃W�Ks�{q�mZ�-Q� y};Ex�mC������]��v���$�2�$�$Q�ϾK���.���b�ZcZsWM�2��TZ�A��cxQ��~m�F}'��'��nv���Z�J1u�R�dA���yiĐ�bT����u�{�~pwm�@�d,�[��,­�[����D�+*�4���1�fee8�Z�7V�m(��Ӎ{���ɀ����eC\-E��l��㘲yX�\�Ŏ�R�\��g"��Ƶ'5j�Ρ�D�g-ۈ�1�Uu��V֬d� ���LQ�鏥��T�G�>(���~ź�V�	��⤵P}�&~M k��dX�0��j�Ƌ����{dK��]>)���j�Ů"_�d��<vF������=�{�bO�	�c٠!ȶ&��F@4�<����ނK�Jx�.k��<����s�����f���Dc_;(%�5'�,b�������3{��,"� 8u�H>#������AŠAk���WtNnZ��!rf�,jm��<�=ܜ�0r���$��7�E..s�PņN:,^����L8�	<��+0�S8Lj70$�q�ë����n�ڮ�,R�D���Ɯ��>�&�Dt�R܀{5y^�|���0<-�x�ҥR|�}f��m�i������<a��Ӛ���|�T�Թ�&G*�J�O�%����u`IAW	=�֔�I�ZMI2>���C�%������	]�m�3�ڡ�5^��WL�ካap�lQN�oю����t��յ�|� #ɫ��պ�%��.��n��'筅.>�`�E�W3|�Nl�@$�ϓy�845���5��P�u�o��n�&�V�;T�����c.��`�7[���ʮE��<(|�����2]��*Rǲoa�A���,��
�.D�b�"�L󜉂ZĈV@�g����$5ՆuD�[_���1�p�|ޥ�;4F�@&�OY��/�����b�TSs��̰�K��228���pgh��=W~ȥ��~���%��-Cΐu�圴+x������K���Z�*�*qAfO,�,�����S,�GЊ�D�����xfP����d�  ���M��!���ʩ�o�����uUn䖗&5�H:� AB�|diڦMYS�5
����;� m�{�����i��[H�"��*Yis����1*�V2Y�2hf��d�ς=����\:�͘���^�.W��b�xO�UO��_��u��ڑM���=��HE4R�.�)�6X���0�%�̦�;K?!�������T:jg?_c����R��P�&�_�D����A�Vbg�@ٌ�فd�򯪇d�ݟ\���,�<f���^3��A6��ضA|xX��撁�x�3�b>]�|��P]D��s/Z�D�a�_���>��=�+���)+$����p�ڗ��DjÝ��~�KH�{"=4�����w���(��@���r��~�>\�����cD� ��>�H"t�c}�� ����m!�X�
cKw�O�������ȗ�$�&��̦�F��]`Z�w^�~����aC]%n����Y8{<l�����t��(=�ץ/�*�~S��w��O�X��$zP��}mIR��n;�J�	h�F����o���
q�I��ۿ;�b��	��]�x�m��e�O<KDH�*��տ����S��gR�2��M�1�c<L�y�\��ڦw�<��t��D�}JE::/;ý8V���/I���4:jnB���YG�f�C	6C�C;���7��zC�(��l�i;����V����=?~>��S{���*lH��}P-z����k%�z$�5����E����hwq���y�Uy����xv/!��BmD9�|W/ʒW�b���b�3�mF��R �@�UE?��C��:��J��7#�ڊ��PѣN洖�8������k���ƣC乻�lߝߺH���GΜ�E�m�t�gّ���p�`� Z���d�̽#e�T�4`1/���}����0FraH��f���QjSX̀
n�q��u��{�Ƿ���k$M�D"���A�H ag ��\'ΰ�f���i�K7�p�R}�u&S��ғ�~��2����C0�4�B��1#��x�nb��`�P�݃T���v��9Բ���C���E$iB�f~�&��*e��^� @�U�����,i3Z��V����ExJ���pjB�X��������U�\���d5�dF��,��2EF�y�g-��ê$J}R#OK+Tn�mY
,E�nZE�a�&���E�����u}�܌�ui��|+�������YF�>�XH 5x�fv���nK�5>=�V��4w�����
+�`���6=�aAlB�B���5}#!?N�񆐊U��9A^����M;��S�1[��:��>�M�:m�2��C(7�L�$�<&>�44�O�|��{-��T��v�::� �L��̙��z��Y�Ū�=R]fP!���}9ͼ {Ȱ�~�g
�g�:FZ����� <JC;�O~ˍ�� ���Y�2��#�x�����`U)>VC��u��� !����q���8�R�rP.���`�T���=����C��١�A�_�jG��P���ɔؾ���J��C;$�6tLF�S6:�Tu��mih2"sm^�&��Ui�zeTX�����_�뿳�y�0$�c�= me��}�~�5�Kp�����e�Km�`B�F�ݓ�n���)㤃�@G�1Q�	�\ױ�5z&���h~���6�Aq6:˟�'�β��@�1�꿱ー�p��X��K���t&VPCp$�}��'L>z�mʜb�����4��Z�$O�qO%�.+����9�����Ǯ��Kǩ:�c�Hg> ���$�/{�g�~I��g	�u2[�GԮS�L�a�|��P���U��-"�s���7Ҍ�dh�w˂S�5�6|��tr$o���,
SoO��ur����~`�.J���l��v��<AM7x=��b���X'��\V�A�R�f��7�̺ �2�-壇S��e�M��EJz�B|�v��GRJ̽�`6�ν�Z��D+9�8�F�"�,`��N��TuHPa@��	���cQ��_gY���@�����q��
����n�����R�-{γ�g�~J�=�����K�����8[��oE�2��^�\�*xቤ��.v[䩤��#^u[P�2=N�7W>�%:|�e���1�Tȱ]K�q*�i�אP>hW���Z�B߭Eש`���:����(j�_�]e[�� �_�//Vi���~��Es�>*�������,$�����5��1uZ�#�� �n	D�#r��%_��OѼ3Ӽ(a��O��񾉤&Ծ�TQ�v����MU'	ioT�t蠚8��$���V�5�t�pAқ#mu�ʶJ/ۍ�T�J��3�es�w�g��ʛe.Î����Dq2ei�����d%:K{ū!2!_i�����@�7<Z�:g�����V���uf�Wh׆�0x��ExW��ǫ)3���kH�����rR�)����l%O%P)�ɼJRo,����P���+�SF�%4�:#��\��~�u������_���Jj����qÔ�xdΫ��h*��Mk�{:|�ؔX���c�z�D�H�q�O���	e��!��"��_�L��[��Q����k�I���I{��y��@{���Ti�6�=f���[(�"��3�82좇>Eu��"o�C.�%�D����@��8yǷ��9TUADu�8~j�a~�G��d l��QU�ҫ�N��&��3}����T�zL��N_Z� ��i���(�p�Ce��x[.ɏb�6�k��WH�.�'�W�ś��qT Z�v��m{�+����.K����@���#V�	B�}�w"���:{ ��V�P��|e�@Ky��*n��S��6W۱�!0�R�J���+�|�mZ����,RMy�4��t��T_��ȸ��Z*d}�z^����ڮ��h�	te�&���ER�	~b{3�L�X�k[@+_p��J�+-X`dE���H�|'�ǩ���1��������x^�1V��i*����+nB���MV�����B����enm#�'�
���-!��(4XP� -iӒhW:�+~pS6K�ǿ`(:Z�JUe��3sz�\uM���G�"�R�S��s@}҃�~��UU�;�(���lK�h���n��]�)�Rp��X��௎,	��>�|�`o���ί�=�����Z����St�>/���K$.��r�48�~�Z58�2k�/,�'Hx7��g��{���c�b{79��?kOBG�Z_��j���S|1�JV/�H�ii��Ga���gQG�����%�̩<3�̩����d�-0NR�(Rs26-.�P44<q��h5c襝#n} �. �E�kw�%�]���*���xn�!�lW	xg$�g1�5���g��3q뱐M�v@�3���s��]3F������0�ƶ�'�b��FJH6�/���*ǈ��l�O4bQ�~�L�W>aY�y஡Io��	�T�R�A_�Kx��e���͒��v����
x�_���iT|~<�|*!v����v�M���sy��:��L�Ϟ�'��\zLt���ϧ��f�a"i�G�9�r�z)�^*��рg����.�[�1�Y�?{��)�6�r4��+��G��"�� �p��l��8/�Zrl��zD�z/�Ddf�6 e��b�;�Y��$�SHRE:#f7.]X��G���U�7����?$g����eA���4d�ؗa�W�}��h���A�8K.���!+m�s�0ޠ;�FLX���ɢ��7=Z!�"aߐq�h?��BTOf�-�jH������0�Mbz��Z6��R��3�7y��������2�c!J��T�Qe�"��a�^1����F��G��]�rۢ�2T�>:���JY�F�k.[}��@s` =C w��=8KD\�"M���8�t>,+@�rQ�a������0l��?��Z�~r���C�w����Ƕ)�=����7����ɂ�1���:7�>�;��e���m�m�S�'ŉ?|���4�R�y�Б����n��۶`�����0'�>$�^��8�T4X��ɺ�94����f�P��@�*/��0���7�8��54hZ���2�=vι,��ٻ�� � tI;P�<�c�av�-J{|�����A�yDbA�-�,%���ui�7��#]����.v�cT}T����A$o�X2ߋM��@��|�f��������ȑmV|��) ��:Ppt�"��,��V�NȷG�kQ��Nˇ�*����@�i�X����2s8�t�C����mP�'�m���<�������ں�0D�)�z�#
m�fiY��|��VH���]����6<3z�)�K�|��}�YQۦSk���@�<�~$?�;ı��@�B���f�^u�f�a�N��h�DF�)�3��|�$(�Ŀ$�U�ZR�����d ���n�Q��iJZ a�TS˒�/�e!�/9T���+L��ʣx�ص��#�>��%�:�<4e�i	ˢLm�d����ؑ�f
��4��z�6'���wCp9mCR�)��Id4G��}�ue���l�dl3&��Z܍cV��窢Ɗ�n�ղ��F���"U2��H�Q���s�����0�g�K_\>c>!|%V�[椅��&�8�kޡ�e@��|2�����u�Cx��	�D3�7YqN@ߒu��[������Uk�|%�K�"u��Ufiw��.��A)�W%%�iy��=%�������q'-�dO����_�������ۛx��)p�.�I~ٝ��&�Q`e�n�����k�(k�D�<.-��r𡩥�l�����uzRᣳ�q��Bk�}!�S�Q��̭�B ��ciy�9������@�P����4p�\�55G�#|�{��� l�A=�	�F� �V�+��z�Zs��2�,����D(�\:������O�p �ȟ�����n�7���L;���b��ن��
wH����uxP#j��Np�����<c|ױ����EC���?4��c��a��N�����Y�3�%�ŌS����W�9���Z�w�ž����d���՟J vU�� �?㾻e�2�1�Q!z��-��p��¹�V1��iՊ��wf}a���g%;�Ne�8Mҝ��}*�Z�)l>��&L�e�	�4�7mE���T��*�pG���&��`F�3��=��T4�v��PE�{�,�ҡ�n�^�Zu�(���(8d֛�%����Ϗ�w����� �ϻ����Ф�b�a��E �O�����������Q�<�>��Y�4�� �M���po�h��{��X���׋�i�.4��&��b�V�}�M?�ȣS��������o��1���
3����(9eo��}�s��Y�;��	;`R�f{ݦC���|��WEh
I��>ht��W��k���ڍ��%G 
}���j��4)���Zhuu�u�o���n=:��Q&�Уi#8�~�W������/���O����-�3�kɪ3GL�`�U	�<����(0lz�T}��y�G���(#$��>r̮WVX���a`��P[xO�������+��'�~�q�wb|�o3����Y�O��Z-���TI����7��ym�avgN�B��Z+k!%��������(���ݺ'��]�O�p9��\�?Xe+��Cř�~��"6�������K�o2��v���G�u(E
'�x��͂�^�|��x #����!���:�z(��
�exH�`iMv�iNzK�騉���d5ٙД�(�Io�I{�:3�i����T3��O8 '�f���Ӓ��חl,-?
X̚�]�%R6̚����q	�AMɸ��=f �P�dCڀ�*f���Xo��/	�&��M�!F8��"���ɑ�f]����:OL�ـ\Q]��֛�/j�b���*��g/UVB~�^�=&9��МҎ����H���У�)Q���%.C�Lm���u��y/6eq]���x��=mM��"1$�Qb䰫�i�3h/��t\�hQ��w�G0���3�k�(H�5S�p���T���������$���8E獨G��~(7�ͽ���D���
�+sp=�VяI�]�`���;��������	_7\�}��j�>�����_+��{k=!���j �a)�u������c�qg��.;�=�����u�q���#�ǳ�� b��=\�\5��:*��XM�5Y��P�2�`[bS·���x�M�u��#��� =+V'#ќ��kߕpR�n�/.yC�5<�vQ�oV"�Y$s��i�5�Ɲ�$��Y���&^���qլ�0����SO����Wf����+�	���ƌ7�IJ���H�K�p�,ɻêjq�8dzo缾�
KR����v��w�M:�^�ɨg(ܨ�����̕"M~�R1<Y3���-�s0��֘S��o
?L�i1X�q�
E18�3w�x�>Ғ*̛����)��e�K|D�9�g8Ls|gb�W׬)�T\E��w�~x7:|�a�jB�������Y�v_�g.2�̈́�d艊 eX��54��M���?2źٍ�"�[�x�Ȃq���m(������P��Щ��e�Dsv�@�g�!�:�W8��$i�{���zZ������šM��7LTE�%�Ĉe�lt�dj��^�U�O��h��rԆuu���wYj�`k�#nB6���VZL7B���G�u�<[$�Ծ�+{�dn��������(Z�b'�@�\xt�[7�tVwS(�S��{ &��'KB�:��(�Mi+�F3���+m��W��t8�Ǽ�G�j������Oon�_��[�1c�d�6�j�^��械v�̱�v�Ҿ�!��EʇSG(��C����b��4�Y�O�)�p�'�׹�g_�v{"{yϲ��h�k:[�7Le�1�FH��+Q��9& ��N1^���\���A��y��WOo@"�9Y�R�}Q�������8��WǙ��:ঋ��Z�&���r�G��T/jA��3��FA�_C���k���r���"2��nMU��ىj>��EM�S1���~���* ��N�N>��#xo�	#�tѨ�Sj���5���d��|�ÞO�t��c��xV��:����*[��F<���%\G�3��[�ؠ^�* -P���o>���FvZ	*858g�J񯼴������ug����B%r�/s�<��Ѡw5"�2�n�C�� ��l}^rZ�G��E�@�-����,�]�
a�<S�E����b�xl�qu���r��W�Q$���Ř>����
- �� �0��������@����-a�����#���@�x6m�b�� �ӣ�a�|R(����q�D�U��]��B�8D�c�8�LO� ^��j��Ď�H$�}O�h
�[�>6���7��,A�;���Jy�>-Ix$���z2�T�R��QN��C,^k
��I��~�-�,�F�$��ڃ����{Sa�A_񧖘/�f�6��%�!{���v�zl�\��)K���Z�/�b; ��W��As8��a6�Sg�d�q|Ye�!�h�À�����R�3��]�td��B�A���9�(��!���m�ìqE��p��;��1���$��#���D��ȴ��d�V�������3��+�g$^6$�b}�����������M���+SEe96۴`�8/����٧�@|�K4	Ķ�7�F��"��gH�{����� �b�9��cꅍ�jZ�u�1�څ?(��a���y`*�t���_���	]S��s*K�<^�Rtz���1mNZ"��Q��F�B�x`T���_躙i ������о�:_c�2FBƆ�W^\��Nk��#N' �𯀴p��:&/t���=L�ǔ�ǩ^��*���"�"�L�e�,���D��r�eG�芈L�&�=�T'o�c�ZI+I�`�!c�l��4;;'h͎:y����і��V�����j��	=zD����QJ��M���WǓ����u��,�)֘��^B:�_�x]�}:~��h���bª�����N�]aM���U��F�(���|BT]	�^��V��Η���=�o��d�����Yw�"��M��c��e����ҁ1j�A"P��,�� ��~��]��o4�~��=j|��U5Iu=T�zխ)s�:�8L� ���:��a��8O{�p�����#vɲYM���м�r��W�-!�m=��{�أXP�M��}x����b���C�]FeV݉���{�mO�������p�� {�J�k؈fՠ�Yq��!�1	5\�K��R�T���<&���x��/7�2�����;:��Z[�"�CjW6��z���f��{9p-6�.�� ��̣�g��b߻�V:_�j2{����b�(����c��g��zGy����J��=oo?� �|����:��ֹ�<�$a^�W�������ť�|)�Ѷ�x�_)�ykb��n#�cž��Am@�����m�l�u�������n��W�cì���{-��~���ɂ~&���]
M&ղ��o�٨���1���3�X�x7���º����@c�l�pX�T`�<��ː'@DbJ^{ޚ1�@��#/bn��7��4lo[�z�s�ߤ��bq_5���k��u�Z�犝�G뺮%dE�P���D(9c�܇���K��'�!�:~�gҀ��g�6�W�����W^W���_�:g4�Ak7HV�50V��9H�kBfv�>�� �34�,������`�ou���c&�+	j��`Z��t,����= Nq��	����c����[s�⑎��"e�>�չfC觥�Tج����<PV�n�k6Up��0���͑{�^�7`b��J��*�8��	l~��V�e%�[�N��=�se��\���OH*�s���z��?j<O��N�-�D7��H��J��F_J$>My��.p�/���GІ> ����|��ە�Afn�̚z����Ob�	#�l0��Z�Hi{�p�d����N���/Ι	ߧ¯�rn2�����
�^% ���.l��2U���~[�A�	��\�G��TR�R�/����:d=M��[�����o<����wʛ]б�F�;(��Ҩ6���%m����o�7��Dv��ũ߉���j`��j�OU@�*�D��
4i�<��!F^�X3��l<���q�Ȁ��,]��i���BA�c|�*b|����nG�2�?i�A���WԷ!\
��2	R��Y���(�x��A�^�:���9���8&��7�:�d^ҋg��bR�`ܱ����چ~��3�#���m�Ľ���8��9��ߪK<����z�u54�7A�k6������J2S�]�c��At���	X 
��ɑ7'2P�:�'F������<�����
_C(���T<325�=����.yYu8�3"��t�گ�L0F��X����\s�#{�S��e��k�m0��� �:�����Qk04$ �Gݱ'@@?��W�K����	���م���,� ��1#��U�kO�B��wu��̔H��Oc��'���_�ڧ�d�1Zc����q�T��9n�^���fϠ�󰞍%�P�KW3��c�|�^V�<�'����rf�Q�b�NC_�p%dC�� #]���@��;�X������O�$O�EpEϵP�yљi�V#,�E"j*�P�k�����B���Ag�6	nqyY�ߛ�&/���S��i�l7�.��`3��/Qs�0Ysf�
Ӿ����A����O{�,����g��f��:��<���GΒ*nw�*LôcH��[4�_r�()�d�A�Y��#��H�uj;�������$�4�71h����+�)Z?K��aL=#��OP�(`5��yMM�H��֮xr��">l�t*�ƕ���L���#��n��s���C	8Z�h���a�i����dv����c�,�i��)"�h��-ZG4Tqh
��2�3�.��r�����3@��o_��y�3~�a��r9��D/���SQ&Ӱ��x�JnSR��v�*G���
�͋��f�g=�4��v1y�x#S�-��J۰�%�7G[F�.e���2
�3'!P�B�Q�&;�b*\�O d_X�a! F��mɥ��Ϡ���~
��@V4��(�1��Z!�\'[�U<3���g��\�\�(�~<�N%�n��w�>�4�Ii��e�`����
W�iCP|��l�z$:����@�{Vhk#�b,\�R�l20;��I8�g� 	}�D�B��UU9l�/�	�c-PB ��M�vtGg#�)Ǹ�6�H�-�'Կ�LzZ��Հ7f�V�&׉�H�w��э�k��� ��^m� �Ev��������g�U�� ��.%��o+WJ ��U�/�J����7wcY��.U��<����v��/mo���,� u ��ѣ̗����5(0;�� �Ax��$u��az+cx�h'�����t��?��U9L� ;oTzXga�Z3���o�d
�{�N��ܯ��яr��Y7By@IrN��,S"�Cɶ$��CU ��n���Gj�I��i~��єJ�'�Y˛T���R�l�qf�WP%(o������Tf�^6�"�)n ɝN؁i�kj�T�~�����_���A���i1fxQ�����}�z�'p�_�v
��YV�v�[�Ѝk=�/>�ɛ�x����T�K�/$��Ļ�m��l�l+�$�\��)tDhK��a5�`6���^'$���ح�el�b�SO��+.N��bd+�˚4zyv
��dx���Ak�n�-�U�/
�#%RT�ć��i����o[�h��"�!=MW�1Hj���B���,�:Z�R��Ⱦ�i	�A� QQT̨�W��Z��i�B1�a�tk4�I�q�^1�+�>k��˫;��9V�,G���vI�B��ijI�8�k����@�ԺYπ?p����]��f����d� *�.����c�UB2�=#מG��Nء8-盓j��+���n��k����*2�l�����;��pAUi���B��e�^L�(+/ٞLq�p>��Va8G(��YW
x�<Ť.h�*A�'���
X�6� �8�,ɟ[��,>l���e^���AV]�b����:!�U��m���Ӝ��B��h*iɝs0���X��a��K����5��:�d���\S��R����V�:�?�3f�BZ)A���V�݇����ɕ�480������مϸY����CKi�2�p�ɶ�aJ"�l�9�SU��T�l�.��f�O`��Ŧ&�g���뢓iT����N0���F�k�;�-��)���AX)sY�3����OEd�kt䘈+�)�B���m'����¥I�H��NJIQ����\2p�Nzɞ�wq`TD'�=�G�t|.�3�IC卑1E�:��(%\-Փ������/z}1Z�.#��=�����P5|�W>:�:�Np��*�����8R��~e�XD�N�.�: {��pֵ��t��PIs���^�T�n�r`1�!�Ck���e��A
��.�BL��k��{A��q��4��RM���A-�q7����?8���˴j�ʁ�$�d��?\��Y��10��H{{?�M*3��������~b����1xr*�Zv;�3oT�r򽐊���U>ak�F]�����d�Eg!
Zw��+���]���9��><�Υ�e&�x�0��z�1u�t~<�}������8|�aD�%�uOl�xBkA�&��(����/�b,��6	����ȫ��Kcz-!���_}lt�o�d{D���wL�`��rZ̳�/�}���z!�]����ڭ�	aX���Rט�����>�I1��F���f�''/ƙ�9�f�,��5_0���X�)h�}��#jͤ�x�G�;�zd@�X�S~}�h�!���4�0N�7{Le1O�&[π�Gtp���Z��o��0�%��GU���J��������¹�]��ݜ�O͢�[�7����e����y|��I����L��y��l�/q��	{�%@�[�7>�zƴ�R����p�m+ܬ�����k�U{���f۾��d/2HϿ<���7�����^�?����7�:�6���U���9r+]�S���i�H�S�I�e� #��]��iJ�&���[%&PEO���5ҷ�<�:�ߵ�t�{�KͨC�`G��[)�s掠�hsZw�X����xH1� �Z�#W���K�������l�剪�Ob�f�Z�Z��7�0|e�9(v#�=�nG��%Pfn�L��){�*�h5F�Y�'���WFc@����!B���:nC$E�Q��?Q~
����@Jݶ�?��X� `�) .����A\c���A�瘬�L�Sϓ�����7 �"�է�U��*�q�d�8DĚ3{�b	����?d�����ς�<�ac��z��YR�Pjsǩ�q���]?kJfM���Qj�X�g�֎�+�ׯ�w2:=C)?����^���W�ɽ1w̲'dʲ��J�K���;׫��B�������:6��7,C�o��u�x�9	>����[�:���j$I�ʔ�)ʞ�:�H�x�L��m�CR�
�'��S]��by���:�`��g�����7Y��L��w3�ډ��Uԇ������k�ş�1C�y�7a�7]��9�#� ͤ:�}��N(k�=�O�`���[��ˎ�T������G�����`��O�0� �?�GZ̭L\�J�P��DW�C��_y+RԵ��<&�qV��kaM����;E��i���Z�Q�{E��B y�C�Z?�mv�~�?m,�c:FH��M'�`�j�9���F�')�<��xɧA?L�m�R��ԅ���Ȃ�:�c�4;�z"���-,���ِ�	ʝ2-��q$]+��//���y��(ȱ�yEP�� _�o����ݶIz9U۷��#���;w(��.zn��'"5��ԩ#���=+/�10<� u�5�%���Yv}X�a$O�2B�2Ap�_�:�"�5b|�k��P�N�K�����FW�\M_R�ց�4���l!�����8�ҳr�j�-�x:�[.֙/�m��%����o����"�UD��Q�܆��������o�yˋHx�������/M)ν�A_q��?��b}�����vj#�966�Lz�q�z�3`m�j�=W�z����r�����9��(�"��O�^����{Nţ��ɷY�]*������]����Haf��1�d!�[N�a�B;��=
x��3�Zv�*l@Q\�L ��c��g	:�V(h1���J�\d�*��c��~�<^�׋�U�⑻1l�<��
``�����E,Pɭ�5�NsQ��e�g��v�Q�`�q�1�P��W] AM�@��T�
��Rc.���V���O���̹%��;3�X�}�^����.U�+�A�e�{�s����k�x�:��{;ї�G�=��jê�ys�������2��C�+�n�샆��8�2mn�鮴�5M��f�[􇯩��"�22x�9כ�d!g8s���S�b�00G�� `EF>^O�S��-r��P��r���,��$%L%腏�!3�|{����B��	��v�l+ �4q�X�o�b�I�̞�H�b�e&`��s��(G?����R�tf�vX>q (/S�Ćqy�+�:���9"S��T��+W���i�U��a�:\rK�XZ��v}��U���z�/��zQzd�ĸt�1����˸w,R�p��&Y�_Z�$i��	�2
�`WHC-,�)� F?hY��$ВCzϷ32K�U넺kH�KU��%d��Wl�nDR����>�aWP����",1��ھV,��*RC�*���$4M�~i8y����|���@��d��$9������`���{�b�������φ64M#9*�f�jO�?}�T�IȺɦ)2�93�v�2�{$Z�r}��8���+랊���tY9�yV�7���X�rF��r�U��ug �ҡN�:�+"���;�QI@�b`����;�s9K�M7hg|x_X��O�JV�I�L��b��*������Sh�)��P������hIa�H��~��{�����j�֎�B��?�D3.�H��g�ɿϣ}�w0�]���d��G��E����b�=眖� �Rh��q��q��j�Do�p����W�*V1�_#�<尞0�5m��^8�u{�^rI����33���T�&�J��%��C��Zr1Tq6ʺ���aO�*	5b]4��5p�!]�}�u�H��@�Fi'R4Z~E
Dӂ��[���m�91���-��x����-·����}�i_�s��%2����i�:�P�>	�5�&�Z@@�T� ŭ<��!�9�	���0Y�=8q������]5��1�c��-���W%)�����iA����	d�s[�&n�W"��;硴gɴA��k,0���@�S2�] 	�V>�tr���[Z/^�����y	�U.�	4���p��Y�F�C�ܬ�]@�I��몕)_
�E+�(�mڼ�Z�ç<����".l��{��bgz�����g��7l�$��(ꏪWճ�����L��oTnaO��d�Nwj*��S}�:X��_H(���tPUs�Ń�� �$��)�{ú�)	V�`3�s�D��= ǲ6�d��orvM�J)��٨#�7����J���yIsd� ��l76��ӊ��H<�ڕ�c�zǢ�(�g}���)S|gd��[8�^	`�t!Y��R�.��]=Lb'S�P��?v{(#�M@&s�Sm*���o�1b������&6Q���D���^���a���Z�>�����;q%���3��Oo|@KQ}ͱ�@��=��n1h �3��\9y��\����ja�G����#���(�|ܹwB��H�5�S���רRRa7&�� �9ҩ! .*O4��a.+Ĵ�HB'�_�ea����r� ���V������.t3k�z ����A�9nf�m����,J����-(
҈���4�j������W�p�Z|���2ܯ-�'��K�*B����S>�Q���S��~�W�`nU.Z�N��\���W7�O��>ڗMvR�=�ҒQ�sJ��"ri��mY�C;%��Ch�<>X���>
 Ɵ�],��A!B�JOP���������gٶ�
b~�S֞-mU�}����(޽U�I�@n*�sz!��/HF�;~ٙ���z���E�Hb~D�J���>֪�aS�vg��C�zQ��m�d�.�GC%)7{<sk����x��!qtE)�ť�δC�y��˨�
���(a~ҹ�v=�f�@��Xvb�i�Wάb�e��'�WL%_6�eD�5�wŮ��l�{`�6/0:E�7@��L�4���M�!�h�Uoh"a�79v�KY�I�۷ BIS�����8-?�w��`~�*I�5��Dl�B@z`J���xI���:�!�|�{vW�X���y�?��l�]���u������&u�ZO���zfUG��/���!�����H,�h�����mj��5dK�2�:"��a�����Zl ��@�M�)cCC�`$E~�[^չMpG��Rt�hz�s�nc�9>ƞ�#&ҫ֡?�u�6�(2��Fh���,�+G��+e{��JD	^�B�	�6W�"%8�yD�qL7
��רqY7�d�.K��x�T���'?�I�p�a�Y�����'��_G�J ��I"�R�t�[��i�����]�u�܏��|����Kb�)7^2�� >j�h���(u��y?">��;8�Ivmu��{.�Wu�8�.��vՕ����������m�G0�]f�Jk	�Rчsꃢ4=���z�0Ȱ�}k�~=1$聆�\�G_�r���<��^!��Y�i���������.��k��z�@�{�Y]�&Ves���=($�PD�z�IY��͛(�4(��Q#e�`�E���A���W'�#��<sI	ZN��l��������&Z�j�R�C�(����1�"��*���"��H^�G&�pU�V�1v��Dc4�0��t��{�O�B�,J��m��؃�1�F^a��,�{��Uw��;����&�Q���������zr� 2��W_�o�B1m?>��d4�4�>���U*�2�(|������ľ�<��y]�.e��aNջ!��W�.�e�;y�K6M�/�	D#8��HA���8�bH;�s��������.tL��!c�]c�~t�z&����-�0�>,�h�֡e�od,]?�$�X��d��_׊���N5=!_ᵾj"����Y�ᗫ�� 	�^�Ƽc~�`歸v�2�@�&E��Β��~#��_h��7�Q��@�����_��=�;1졽�7���M�]KX	��cs�4�e"��ڛܰ3�cZ��"�V�����b����W�2�p<���/S����&m�ޭrf�$t�w����X� F(�L�ʛѷ�]o�T;�`u&�U��(�|b@�{*/��5w���"y��_u5���K���6���w,��іH���R��;���*��q�����>/���F����&�=Ή�:��-�
s��Cj��#&D�Pz��]�4���?����걊wj�8��c����\�V�\�Յ�DfW ��@����E�jM���A���z6�z���"����l$H����`l;��V��z�
����.R�e���{�?^%Ouf�ok�;^��~������}
׮������]�T˽ԱE?cq5��d�
-�?B#��y_��7/��C�
4 �c�`*HGg��.z\��߃i޿~Qdg9�kΟ����l�0��@/�����4��h+C̧�%��%���&��g�m�����1d�n}����deػk@s���H��;�����#�!�;���S�~MT�g���z��q�_f�{A�����(�;alO2�H��r1��(��� ���"�b�w?�p&Vx�&�}��S�f�vu_7��:�\}(I��Ƴ7�=#���V_��1�h���6�,����I�Q�Lԡ��?��7�~��VS��:�3$,1�x�\�SgV�w�N���o�X��%�6S3ОH�UW�9�N�[1���%U�����֟��M�#6�j��S K&m� �����v`�|�*�*b�8�G�0���t��tNJG񬀋
�ƞ�l��r��/:�T)�����2��+@��5�n�����z1�Ԅ.e�9�YYgE�7��M����)=� �;җ�2�jg�_cAgy�+|M��iJ�|Do:��B����!A����eޡd7�F�sY�((�1�c�#;_|vT�~�f@SN��@�����z�\6�3c�|���jO�K����\��אKĦ��y4ؕ����g�|�}�?�(U �T��-k�zwS�)��!�h g �A9�n�g��Q�0{�z�lڕ��mC`nk3�zc���8�:���7�@wa�|�}
��f"R�:Y�=��:��z����b�:�@���U��2�Vy�	�ڍ/|P'� 6ޕt`�w�د Y-�����5j�I�sh�Rmk�~�u�'3��f&EҌ��Z�9�_?�6�Ә�d��"/]Vx$9�Tm�U
�9��S��
��Y-V��j��E�SR6X�g;8��?�z���r싟�Z�C����0�{���-�:?v�S���m�H�i��Jq�q��$��O��	�-G1)AX�� ��aWv��"+�Q������,�9���יhׄ��E?ϳj:�� ��O��u�C����w����w�������A�X�0�8�� \z�t�0�̒�D:�8�Fc4)��̉k0�����5�0��������҆�(G�Âr��%@ī#^(T%�P���[<?��jʪ,�(���+�g��:�+���~�]�����C>\>�V�/!*�wM4v���]�[l� :^�)c���OZ
0�vɆY���S@~�y����l0�9Va�А.�r�m�^����Gi��,�)0��K`�̛��
��v
�9��:��/�L�������P �O����t:��j�������Ʈ|�$;�G%}��h�����K����)&%`3�~죹q��S��^�-��u�J<b��S�쁼f#���ɴ֝�iH�>�4�hV�Px�y�ne�c�Ro�fnB�r0�~k#�{���l����T}�����a�gvx�N�g�aoE����k����#Ho��P⒅7�MKQ��	�.v���C0	���I����V�o$�fU���nGK����q�IFmv��Xb�+(�V�.VA#G�Ec�(��o.�b^?'c2�dy��mR^+�VH��^ębN<�'�ksÉ��̜L-q�\��q�����o�֨�W��q�]�����︟��cQ��<ژ)%���W��3A�2�qͶ���u��E����������{n��k��W&�H2��z�
6G?�R�\>�G�©�+��(UM�������(��l��B	� ���?d�1���)��
��\���ZO��? c��]7���h���
ٓ恵n�0�� ��H�I�-��^���Ԓ3 %?0^Q�	J�X���=�v�@�3�ǆ�YЖ�k�����lGM� �j�F�~*e�K�Z%j���P\��/ʀ,���;�� ��Vct5�kZ��Y�L:ޢOrg ��ݩ`ѧb E���_Lr�����m��)*��}'٦,v��2Y�ZZU��(�)%���ٲ��3�-���=ѢI����M��y�o0�.��m�&� )��h�`��`ڭ֣�8*�%$q��F�2�2]����;��V�@�o�?aב��n�hA-uQ7�A�5`�?�hسJ'y��I�%#����wI�Yw����k��*��y|�b.I墿ЄR%��=��ԵQ���~ن�u��&6�	�^�\?]Ò݆1:�2z$��;<}��+p��ܭD�I���i�Od:��Ɩ��9�6o>��,%�v�ߟv۹h���x��ӰƑ!�f<b��MN�|�{IFm_6��.Y�������C�<�<��+��
:��Ԩ�=:�e�jl�Q���|�r�W�*p䬔'
�bT�~S��kIæ%.���ר��Fl$���m�����Z�]�u!�������GęZ�
���^��b�$��6�v�#��ӓ�\�v���Ȫ@D���_(�/�%�S���FҀ�?l�q\�]��l����<�eR��P��x�۹���l��?�=��UK�}4(갘*��A���ǲ�n�;��v�kٚ�ŵp	P��qzW�3+f*��&��E��E��&(&�@ꅇ`;+�cN7�KJ��K;�=I��(BcE��܄���\e����h��ؽ$*��`��NHҞ�<ȿ���(Nך{j�9^)T9B���)Qf��p���Չ��2��.�Y�I�`���V9�ݺ-��e�e����"D��{�����f��9?+5ޕ�7m���kH��@Վ���\�Tc�m����T�p}ƙ��֚o�&s�Z�����]�V#hJ���IS��pi����Zo��g�x�������S`d���[""��!�Z�rRE%�����(�H��M>���{�)�b���s��V����\��ɒj���o&I� f������Z�d�N���(��d�m�Hٿ6�s�F�/����#2��v��2�r�#���\aͽ߳A��7�Įu�*q��Tf�2V������h�C)�>6k�v�w�`��,:�$a�-Ip^�oK�}����4S�����Ҷ.�o6R�̼��5jƆf�-�'�=N���<�(�f5z��M������"�˼$�OY\�2�Ix,O\��7;(/>-��f�F��X�[������d���:~n)�����T��[�� >�J8�nȋ��1�O<>�k�.kt�Mht�H�N��B5�H)T��7�!d:s��:�C��B��f�JE/�n� :>.f(
dQن�	Tz)�V� ����(�Q
��~E�RK��.��?���9X_�����vm�����O���\!��	7��x�Xz����ۦH�����'�b�m�1��o-��WvN��p=�IP���$�����@�" eݍ��0T���9:}~�S[YH����õT$��?�A��tE�Q�%������}��w{��5z�mF�t�h�-�:ɵåo��z�t�b������.��Fm��l��s����K��5�������+���ͨOu���h��^��A·��S&��\��:HJ������y�o��Yw�����-�4�m�[�R�ȭ4y>24k�V�a5m*H�?���
�L�ѨjyIߡ!�o�w^��Ue$fk������c��1����'!��W��P�0jH�E]צ뇒Ԩ�tBJ8>��AJg�)���_�,"�oɰ������N��{���rA7����+��qZc�?���V��c	YX/�P=��d}���[�PTL�����cX�����Bc�N�X���'X�L����j�#_cQ���7\��{�t�WpX&B�Jț=e�O#궴ͤ�JP�0˨�Z0��� �y�6�uME��a�O�,���%��ԇ(c������V)���*�j�W�+J-�é[���������V�0�~�fc�~��:t�M �t�k�z�\�1��Er�m�:!*��Jߖ�h�K�GR�&�3�6%�È��_���,�ߥ����]�B�k�"#s Ѭ�{F�D��t�TSj�Nt+2r���M�ڂ$NO�=��B!0�Tv�~ǐO�I���-n��Zfū^�)+�8qq*p�^�0��L���8����t:_,EX�f����7��)��8�-�X��c�]o~dձ�0��zsc�flu��лs�Omy��+3;�uFx�~(��B`H���5?�,��",e^Bo����ɭsU�e�k	Z��R��PyF�� �<$��d���$�u����Z-���#)A"�P�F���C�t�L��@��@�	�45�?�*��߂T.�h~q/~n�j�u��1���{k#��0����T�?������a%_��d��l����+�O��3�^��a��F6,��$d�kFT��9�w��?��pԗ�'�H��I��|lZ��Q���}����������4��wϣ�-�K<��6i'o$�5D����;��\p8H7�K��iw|���mk�q&�n��Hx�u��ϒ,b���ȟ��c���\����$����\A�{���,�7Pr�x�*I}�%�V���%��YN�٦"�C��<���]�����ԔF6m�����gK��4�� ������^q�P��,�Ī���T'x���g1a�8o��G/W'N"�rH���
�\���x*C!�h���u����|�2�&�[�j~do���1qr���Q8���gu���]���ri:nŪ�����{��Q���d��#�.�+�[� ��X��`� m�h[����Y_/���MUKh�v���{n��b����8�[�O9��Z}w��
����.Kf��(0�j�����_����L�
�3u���X��E5~��:�~���e}��'I+�ѻ���32:-���T���`aoUz�	A�v��v����L9XU�r&3�^���r�))RƝ��!�� !%�=\� ����H(:�/�Xt��}E8X}{x�����4�V�A|FudW��3�+$.z=/����&e�.)�B���8-솀�8_��x��	�d��I .������B��(^�A�=4� <��Z5�fR7$r(�*)Q8ES;��`��Ϩ����+�V��B��{��o��y�  |H+r7k�Ƚ�����y����Bx<����~�[��-���h�u[1f�D� �"cQ�^0�S�]A3����2t:S�ۏP�W<��i_�I�!�i���mɔ���/O����Uv�e��*�uNA��Ə]Ps���0���3���{V�xW��
8���0���%�i�[$S���b�1���2PQ��!�Nm>C�zzJ4�ײ�x0�f�K*C�VT��O/�	MF�6�Tqj���l���*oJm��؉7�~��V$cf�
{����,�>�0�� E�+���h��C���K��x;9N�"C���AOfj�A0� �?b��f9ps'��s ����j��&��-��a�M2����X]��\>����
��l��^K5����P�:fC�џ�Y%�R���$hj��o��-R�`*�a]�d�Z���<HW��^_t>�эP�-$�SNʸ������	<��(q�603���z�Hഛ]F�E3�;��!1p���j���v�+�w�p"�a����d��.�4_������H#�������F�Od"^��ڦ��%�a;+0|L��[�s׀ȹ��*�"�i�n��HF�&����{hE(1lgkN�խ���!Γ���P>VEsH<�F�>��U ;��4�Ζ8c�p7�q����J��(���V�.�Nf��

������g���cY�S^����D�m��5�f�QJa;��/^5D81ز�5h�%$x�.%��,lJR5������ �;�_Z]Z�BV2���d�U�z��?�9_�k�Ű����G���b;�?�*w3�޺�J�����ִ�C�`k�8I�j灡LZ���R�J�=�b�R��W�	�FL�v"|~�I5��vS*�s����0,SK�z��0P�1�}+OZN�=�`}#�X�}ؐ1 �k�������ǂ����
�#�3 }Q��Bk�k0��c��,��t�Mh=�ep�CT�F�:Z��������Ց�*m!t�I��F�}Z��@$�)+SUݘ�*(���p�?�s�A+��9(���ULF`�h�<DM;x�7U� ؉�@�v��0<6�1��l�Sݞ]̫3%2�O�8���d���A��x��5*[�S�_<�倭�>�~ޕx��"{��)�/&D<�Op4���:�Q)	4����ty�*y�HP��! ��^ۇ\�g��L����nG�� >S���;jO���峙�=�4�M��[I�"���eＫ@�~�}-��
�X����P=�����u�8�E��\5Yy#�V%��{��<��
F�9�^<�<�X$Ϊ���������MS���A�c�6O)6�I����~�ݬ��I@1��jIbr�(R�J\�e�:��B:���`"��"?c�G�x���bdsL_�I@8��8�i#g�āXY�v�Mb޿�Pci�߿{d�:���|ӡ��g�T�2]���	J�9���D��Ȗ����!`�d� 4j����÷�9c�N��I��AB��������s�Q��UCj�~c� 9eu&B��h�M6�j�-����b6��J�c�9��ƱU���.�+0 $e�8M B�}S�����W��rv��߉�c�Z�j�����O匏�g��AP�P@�Ҩ4�<K">�x�*��c�%��͗�-L��f�?���)����V9+�3fD~�_�	���h��Z �2##�5�E�@�1a�0�u,�V%��,���Y���-o�0�+>j����s�n�A,Z�&#|TQ!��f��
�Ci	��E: `�Y���k���v!��IW�'��v��hh�j}2l�{�4��q���KO���O?e��w�ʣ���\RZ���F��%�~���ˈ9�6N�~���/���'q��$�<aQЇ�h��O�-Nt�n\���Y��y\�ω�Q�[�YO�wW�q��J-:�`����M���q���Vl��j��\,�1�N��❔����j����V���o8iF��^?Mq+XÉ����7���{9���oQ��L�e���Q�048`��bg�ґ��aX�灸PF��+���Y�6x�7A�}�HB��v��Bp��i'��\nmN�Y�}O;�u��r��fZ-�	��q�+)����@���*���v�Ygs��7��o��yQ#{��]8�����k\`=B�܅=ڂ�����#d��6\���X���]�_6���R\�R�Y�ފ��J��=x�yޝ+1p}�=� �*�b^$(�>o ���oy�x���Å��!��P��h�� ЋF$�i�%����0d����ǆЭ��>�`���G�ˣ*�N3ef��Ƿ/��)�Y�pR;��[�q�:M���Yˈ����ݞ
91�E�Z*^�0���z��P����I��jI�LVюV�i��#��vLt��f�����C�;�&���چ�0��<�Y����)A�W��.��6i{D�Q�B��k��X�~��$�n��+p�?�r��9��Uj� 7��X�P�w��З���:y��C>`�4���s0'���Ė��W�̈=~¸�L��t�#BBp��u��ʪ@�"0g�H�غ���������w۹<���(���";��Na=��8�".|-\��[,��[tIT���e:���T�*N}*<�Cd�_2߹� ���ў����='����ծs�CڰkU�B��{��k�q��Љ�����weW>�0M�m�0��~�������*d�b���}U;3Lε�!dQ�_� ��=_7 `^�%�/��]�G|�;N�у�p����Af�[�,jP�ʖ�-=�Lg��1ίD�����ܧ���)U�y�hkeϙREM)G1��kKI�6rU��G�v���p@Kd%��]�A��������oD�=Y�5�6����}m��܏޹�͕�X�N��0 o ӎP9
S]�x8g��An+_Rb�s�utl�z�,�_�@�������S���Y��1t���\��T-��j�{B�F|��ks�n��Vi�/7�C����#=z���uk���O���,[��w��Q~����0�8���FL�t��S��gd4/ǘ������G����<��3�Wa[ƻmp?ɋzۏ�EIP��s'�ZX�8'��-�`f�]��è���ǒ�9���
�)Wߐ&��[#0'��RTeN:~��67�0?d�bU> ��dh�<��$���H_��6����r,���J�_ZG��0ʳ)��д�@��[����u۲FA	����ဂ@����#�.p'��e��s��&�wM�%Q�QII'q����X��3�0r���*ܝ��9�����;Ö"?6�qߑ=(��>�IF�ݕk����8Iv�%v��̒�9�2��4�b!�l�fY�t0 ��6[���,������@c����*M��:�KQK�D�N��ꅱ�7�`m9eŨ
^e�������v��<%�ٛ2��E��n�2���2(8Gr��-�d�k4K��k|�:bȞ� �=��5�/���m���
��٩���q7�ȯd���{�)���^ps(����5�2��v+,��(����	���n��Yn�6�SXA��ڹ#�`)��34lQ��.���&.[i��!��p����0�$$��(�ިۙ��g2�0��� �QI�Q�>��	|�C]+�w���Q� `-�H��> s�v���X�C�(p���W��j�#��f\`Y��zxPвK~M)�-&l�r,�M}�_Σ��A��*�Yt�P��� c*�x���m@\�3BúΤ%�Y?��>ѵ��D�h6��˘h�l���.�79��O3q:಼��j��#s��c�j|>h��N����Ym��9�f�5-���S��5�CDldY+/��=�x�/m���j��l�0$��M>�en��X#U<j��~�#w��#f��c��qO�	wT0�t�(:¤�ˣ[�2So��:���MM(uʇ���қY��ıRF^*ov2Zf�x�U��D�g�e��Y���uZ$[��pf��7�p���LGՇt��O��<�G+2�D�p�&�K�~}ɩ���?��BIOǖ��UC~Ɏj�+z�h�E��C,LQ��qw��� `���4��]�m�F�{�؝Q���L(���~�NO$^/��F�9�V=lT[E;PM?��J[D ,�?���{���q��M��#^&,�\�c(�vA���g*N�៞����+��o%�Ȝ'Ӳ��:t^��x������.e�Y#�ݳ�A!6%�֟af���2�6fo?P�-%YIWy߽�����ڙ �5 ��n� ��|Us��gQ��!�HK�E��.�Q�`��W�:��u�v�)*t�����8SC߁���v������Lz�J�rф+���'��G�n���U��%�tSo�����z��(7�P�	�	�e��HI+�(`�>��r��Lx�&���&�{��I�/����	�b��9Ë�y�sX!K=��ub��8�1�M}V���_Tw]}$����K3T�ߝ�Fֱm{2Ѫ�܆��Ewc^�q�v\1t�
r(W�j��ޖi�1����K�!�Z���'�ՑG����������T[K�V/6gPش>pJ�@�4�o�EٛŖ1=�<�"����RA�YȇK=�\r�q�!j�Y����7MQ�#�8�M$u��.��/���GZwKol*�Y�pϒ.���
#����m�!�Fs����J�M���p���l%�^�D8ZJ�T"�z�؉٣uT�����d\������N�����ޱ���C��|;��~��<د�k�%�/cFKU~2���a;�9��V�4����l߀���0?8���`6�a
��='�~X�8֨�����
=�=��7zk۸��8,�:i����L�h��^�L8�DlY��# <��х�ނ��8ذ�I<ϲgҍ��)��q�Y��BJ��Z��[I�[z.���ey����KLn�-1n���gy��z��^J=�mꝗ���Sl��,,�:4�q1\���%�j5��g�Y�E�������X��s�OpHE\�<��j�tи�7M����U�/��欰�x�ݩ�x���4W����MK&�vZB� �)p��K�0���w_��+ fiZiP��F�wT��G,�ߚ��L�������E��8�
�8i��]�(��0�/)�)y�'���c�ߞ�w���;'�e$^g(8�0���ژ >���e�F�πU�b�8z2jf#i��=y��y�3y<AY!r��'�a+�|�@׼C��4��S%�M�i�y����\��vIt,6���^�u1P����hP�P9\̫�8	�պ%�J�B ��G���e����ǂ�[�5)� ǍLD��̹!}��r�1~v��Ŗ�:H��Ɇ���-W�ۙ�!B�Yg�X�X��)�ƭ�T�8�Pf+������m1�Zĩ��O� ������2<�d&ɭۑ	!��.IX�m��O����ꭗh(B*�YG8�W�	����n�����M}�����[;�GY}w^��ߌ�ͮ����6.��hܥ��&�S����F���2`p$�Β�|��ۨ�.��P~�� ����h/6�'�Ë*�������O���iey����J������e��nu�̐6���3L#��M�()��=�p;z�N|]t���X��->gݥR�p�o�5L.[�>��O��=�FjI�]#Ⱥ���,��V&�����	������sT�q�����n+��v�&��
�X���4ȕfrlW^�S�n�;�nv���=�H�z�&���v�N<��O��&�PYX��KKW�'Q!0���%�����W�M򨝊�i����7p;ܯ���6麀�b9l�$c���l�#+?[�����5�̣���;-�\G�)��X���N�g�\��ř���q�劕�R'H�Z}^Y��7d�7tl�쐧sE
dDל+�tFw��1B�n��R\,"�yo�V�6��$ b�)e���˕H�	c��e=�am�Ydc�b�P�*��{6,��啦����Q�M����fv�>֖�
�X��.8 �0��d��?G������k�8Bqd'$̀��Тdq�g���f�U�c��T������zF����������1p<'}����[S��ELH���v{��x���R�-� �@��D����$+&Vֆz(WS�S%H�r;K���z$�ʥN�a�]:Бm�֫z=3L]���Pǰ�WŇvܰ��q�K����H�wσ�=_��T����P�)���G^r�s-�N��%J�]@U-��{櫳��K�I���[�(�$�D]����R`
�t�~W�y���?{�o
�\>u���S��1��v�C�ԣax�I�?�q]�����ݾC�oޖ�6��=�<���>�_�3[	P����sJ��p��֭��;��24�FK��f�T7�}Ʌ�~#gЩ؁}�Q�?�줴����@��C�Ԑ��k�#�z㥈��G��'�T%8����� 8�1��KG�Z��Zo@������x�I��"p�٢�B�儽��,�ǂ�l�X��[�3���_XG1!*�	-$�t�M@3ݬ������rZ�v$��t2]2�%GJ@t�<'���p��aml���K�E�p5��vW�[�;�]xZ#�+N �V+mRD�Kw%�3z��-��*�a�j�(���t ؑ��
��i�2����(oW�s�>E$�֭��
�G1��N�ȓF+ǽ�?K�}7��4Φ��-�4Y��R�'v�G^y�f:Q�6�6W.d7�P�R̰-���J�����>W�T������$��@`�+p.�+�
z����v�[�Q�2�����ѳCc�Ō%��3��ZF�.2�G��&�o�b�0$�DJ,Z�^�%4Txͱv�{���E̳{v��{��:)�������vGZ+�[wȑ��B��s��'�H��"*βѕ}����r*��?6�fc�<�S���N�������a/H�jey���r�ڛH7x�������4Ym���~ �ݬ�\��6�En�|����P��+� ��� !~@o�i�y_�+����r�N�&��z��ȱjcw�.6���,����ĉ'Z P،-�>1���8g��?��ٙஒ���=>�m�K��`8�g�D�k����XG��$���5��t#R�3�5�b�_p�w*^	P�	]�)�J��0KN��r�Fީ�ԧ��������'�Lz��fj��f�²�^$���6�@�e�{�B/8�<����\��Y�/rF� 2��SXi�JX/��=�I�oXu"L
�#�[�D[u@�,w��0��}ޯ�e�[�������Q��#Q��qx6x�Ш����h]���k��<&�
���H���|��+2��|
�%X�O>H�Ƈ���D���G��
��1�z�Wc<;a�C^�����pKn*�[�P�V��VW�G�b�+%4[�zQG��N���_��J�.�+9�{iÜ�����??S�A~����+�#���wdT�֏2��m�`
��� ^(�@�ɺ�Q��E�?�����X$+�`�A�%+9T/�K�3깪��1�=�Z"*��E��Q恇k��|�L����%�6V%���.��@)|�����3�}�k���! h톼�ޠu-����h�ל�lHd@,U���cS����"H�]���}d/�y�Q|2�>a֛J����}�� ����C$�Ўg��(8�z�7 �=UM[Lc�(Ŧ����v��I����+�|��Ƭ��N�7�Q�6lې��"�F'+�G �>��vRx���-A���T#���BA!����ܨ:�Z}������fX�Pv9-0%�l�zI��������f���3JLa	�M��+��G������P��ݛ��VMx�V�����d��~kk�zOJf ��s�Lh�	��!+��ex/�-�\�D'�h���f2G�$�>�9����B�h(��%S�P(`�	D���$���A�J�9�e��H�}J��E��3�a�|�,���d�'���R:uq�ɑ�H�oU{�f�I�A!-M|ض�+,�4���
�iHp��41����V�@�Z��������3���u�*���mBg��u���+ ���4J�g�H�{�����fs�f6Z��De�ߎZ��CNF~Vu�+�����9V�`�\W��n��'�'5����dkb�X���ğ�ڝ���g���U��o1Vy�oe�{;de6�~��J��-���&n�>�T��+��2dǷ
�_�Ʈ���x�#�Ʊ����P�fo�s}��(�H]����$r�߮�]��������B���Z�2��.��Ԥl�/_h�u7�xZ��S��3����zQk�^0/�#狋̳ǥ�|��8fsg$U�޹����%��f^���w�,&'E�����4p�R/�=�.�rE�x޺_��]��j$*�f�+)�BQ���3�́0��~l�Xb�q`���F=�d�]�D��G&>%���ȹL^Mo��~�H�s:\�����w;����������$�lR�kv�Ne���`~$�&�I��A��L_,���P��.������"�V6��҄��þ��L!�I$�8�*w\��e)��؊�z��2��tx����exhs�MC%N{�B�RM߅ʚ���)�cǨ_)��u)#;�(�+���D�\p�.��;7���P*�%���/-��Q�y�38�����2�s��� ^���xj��:&!��b�sO ��j�k�����"��2�h߾�����!�I��W���U�=ǌ�&y02�6�-0�`�V)�b��H��[fqb�y?e$�yFz�	��8�t�jGl-vE���ӂ� �5bV�az���n��At���Ϥ�`��Xh�ԵS�(��<�s���M|���K%F����xwS�y�����Û���0�����]�V��l�ys�^����/��=��5���uB��/ʹy�*�6�/#m(#�&*���*Y÷)w/I͇���n�#wc�]xHE���~�U�n����f��%�'����V�K�����@}�؂�/���[w?��b={�^�������NȄb}��$��}�xwԇ�n0 ��P����hNa�L1��V�iLm5�z��(sޒb�؏���NFj� ɐ��Q+�J�RL��CQ&������Uɶ+ԭn�����R�(*�k��N�c��rV^�T|ޥ�׫���j�G ���>��o�����9_m	O��u�0���f5$�
(_��i,>��㠪YY�������r�3�K�}m�C�j2����c�'T� ��ec�&{��Ճ��_�����Ӵ-���=2v�ۛ�_���J%:ÔB��ё[��u(�؀����8}2]N4_���6O+#�ǂX�N ��I��ϐ_q�����͖���a
�G�/�#�����=�S�����&�����y�/�kqA&��'��aL�d!3]t 4��eJl�#��6oo�v���6�0?ҲuDg�G�L~$nl�CtP��\qNd
Ww�l������-}V� B�Dx��/v���g�<�o�u��:���g\.��iGx�pw)2`�a\	����fs��'�Y<�t �%�
6��ӯ�A� ;�f�`_�+�H�!�� �X}������y� ;>�V�&_���ԑ�D�ދ
��X��?^�%cMs��w����g�`PS	��C�����z�΋��Y�k�8� �
�5~��=�����ly~]�~�F��ȃI�<�F�F��9��I�C�T�t��v������g� �+	HE1"Wɀ�8=OWD�0�^�,7���E�B����`~�v�+�x��Ӕ�ɛy??�GN�� _X�ܴ�s6��"|r�P����4��z�}n��3��$T��\��*1���1(�H^��͌� [�j���w�x~8Mg�b�G��Ix@�P�u��8��;[ѩN�O�o���^�C�_Y0"߬d��xf���`��f�%��<������t�د�)ՈzNoR$;;��"�I�)o^=%�C�*���I�R�����2�6镏�Md��:�k7�� ���ʙ|Q�����Ґ��\^լ�u�\�W�6y�C����`�8���-�#�8E���:����SJ�E(�rf��cGS.$�t#�ru��SŐ�����<��w��j,[�q�yh]����UĘA�I�S�P�$x�� Q�B��ͭqE�̰�c�ϳq �����q(S�����?P�� ��`�e_s�����hP�6�O�Q�6������]ݽ�xo����i����X�zE򸮯z?W�O�N�b�os�m�Ɵ/{�ro�tP[$!�%	ac��gݳ�)�Ly'B-U�^e�8w��P� ȁ�Uo�s����i;��&�R���<�8VLl���_>�����3[�+%���?Y���u�?�7s�A�����aL������Y=�zםV8r��c��Kx0v���(���5�%�M�c���L���]�	��h,���l�ԅ~!�h��3�pU}�<��	=v��\4��H��D:p�v�{܊��#���:�)�� 9�Z��@�Q���k�o��+��4	8��dY�$"jz�"i��19�r~/�1��,Sl��������.�S��Ѧ}z�1S ?q��ҾT��0b�-<���D�>�C>�����/��W�X����N�zαv+f�{�;�U|�}>��孎��2/q���_����WS���m�NN6��H�1߰*�,,�-�.��A�Wj�m����3`��r	x�j�N�7��A>S����)̮��!��'���!"�r�:��Nw�|�v���lmB�Y���<��T�/���.����|�5h�cޫ����`'�&��04q#dͯA!���j����&ըޮ ���$�N�|!�/���Y��E�R4����x����Djz:/Z9����)o4�9�p�(ΫCK�X+�G�H�#����������B0闎�z<�}S
n��D��KR�F� $௙M52'ץԿ��za9+U�#J�|a���[u�b�{���M�EV�EX�Z�h)q��++��w��dr�*��������˜���.z�Ֆ�I�.^�BE�CNw��5���`9` hJ���E�XO�����3����u�Mb�a)n�Uq򶕛����6I)������HȒ�g�Η��9�\1�����<֓{��e�ފ�}>l�~Hr�y��Bٳ��Kp|�����=nAt�!�L�3��9�rR�O�jxu�������Ԡ3�Aq�z�DJ��Dѥ~ĭ�{��ȭf�d�'���.�,,}+�����;��>滕��j�L��l�T��@�B����>5�t���g�it�U?�KZ< �d����L�5��+I%!��!H��̆~��5ԩ��_��©W�x
x���M��{��t�;(����1y�`�#6�D���{ $�!,_�������Auo���F�wQ(t�0��;H���:s��(�����"D)�2BqZNwЭ{Bg�*sX�}����)V�W�2%V��F�{�&�͈�ơ��.q)��o2[T��*β��ԋY�lm������4�H�?y�3��D�@%���arl����ܢ��mDX~H<�N��1��a##�����,� �r�2UZ8�UA�$���o.C�OBF�>&�ފ�V�Ql$а˷U���R2���(˧k04��'���"�e |��Q�f�x��!A���Q������9�=ϒ�K2'Km�prl�h��������*=��g�*����~�}a*؞�uƒ�F�! 6�2�o��A͝���[�+J�q�`,�r�%i���#zp�`XѰ� ���,��l��1��5^O��_�J�ߟ��?}���A���
���X?�3��ബ6�ɉ�l��v���hgt��[ ����O�e6��n7�h��q+B��Q��Sc�����шN��<
%*�Lڞ n���|�EK��>}(�#�7d��=DE�I��`��*���$��z���++��c��%�L^����sT,�[�A�V���B8/���ghG���V�,呶����y�~Z��9F,MF���Em08���ܾE�]�>����<xp�S�>?y�K]�4�Ja�H��5��b�
�S�t��tE&*�Z̘�K�S�z��j)	3@C��p�Y
mQPdɜ�<-5ж��a�`�K�ܬ���d�޽�v�(�2�V₀��HV��en��O(h�;��6Ct����2.����>�����(&7j靆��sl��1y��v�д�P�]��AW��1������\�U���:qBi��рhZ�XG0%�t]��/Zk���ɞ�0KW�Vh�������4�
t���;,�8��۞þ��~ږI|��Jy�|�v
|V��y�ʭQ]AĎߐ��O�-�i���ĵf���0}�ؕ.KD�y�z����>�d������@�B����C�}:��<����f-1_<�9�z����2@%�3D�1�r���e� M��X1���	����n�����ٶ��ҟ���	����d��3E���_f^S��Jz�u�V��{M��{�N;t�a>Ib����o�МV{�W����3�л̕Ϊ����+�e3B�|����s'~�n�B[�[�p��~c}�i��O ^�g�~?�P�NW�&�����Q$$��%sCLD���O��s�[A6)����`?�C����@��jY���|�d�`��<��b�
\���m��&k�X�7�:�Hi�u���୮]�R�R*U�}9@!�g4��c���Ϗ�}�&�GY� t�龫�Ɠ+N�)���E��ХtzX���_&҄�5=��UV �lBXʨ��n��ET&H�s��	�u��kJ������7C�>FW�c��}�����U`�1�kYOI��w{��!�}7�VQ����372�t�%I�������|}��c�{��|����9���m)*3���gg���ʩ�2�K���Z-�[L����C��?pj�R�E�I~������r"G�ك�}g���e���KsWi>8�<��t�s�XR9�e��R���[N,x"9�e�JB
��}:�Q����U���nt5�r$V���Ҹ��^�,<�S_/X�N����=���;}x721�8�;+��c�D���v�(H)1�;�UF���Z+-h�?���	"�*�H��w�/�-�W���\��"���7	�p�9FJlƻ'�S�����L��vB��ڠ�R�^S|cƊ��R��i,o�D�)&J��ؓ+y׫NB�l�ߧ���j�$�x�H��i���2��'�P��A�Lfv0-�l�[�v�����ܕK��5���]X3�#.���w�R���8W�%v�)h�_�A���q�-�d{S���IT�_���h��L�KB��#~��9�Wû�]@R^��-�'c�/�S#͘��˜�Èc{�s����;���M����w&��{k��7��K.m"v�y�aZػ�D���7��{��nb�f����Jl����z�͠�B�Dy:Q!�#@�a$`DK��+��8�B �Q}m�i��Q5���vy��t���	o&�?�h�Ym#�8M���\p EF��e�F��W.�v��z�q(�ňBq���ש���.�,��b��N\γ��h2d~����{�Q�XJv���Y�.��d�P	�\�@�������KbM�}�2��K�ꓝe��FU�F�N�s�g ͕�<
�֝���UW>3����ڝ�7��9�&�ÍUo���|����d��`Ɣ��x���O~���:�R���[R�����<{�;\�eQsO�ㆌ$�~�V�}�oǄ4`�>�d�|�B,�F��� ���kS���N�E	���n?�󅢋�)<d���������q���︹�$�J98�.��S��c()GI8W?��9��T�����H���Ϫ�GED���>kO�r����`�Z֤��M�������\����4$A[�c)�,�`M/
��,��N�Z�xS�bΠqrM�ا;�������2���(u�4��M�8�$�V�&^��a"=�e�4Y&Dp���'c���k(X8gH��v�`d/I�go��3Pc_LBH��l��.;"��T7���3� �	�I�S�2�\��v��E-i;���2 ��R�`�`u3�N��M3�;eO�F7�;�A�4��HDCA]ztw�+���S��!̡7G$�;"=F�cKB�:|"����`u@�n�pѧ�T�H������;�Z�ًM�9k�s�UX[;8��& /����lo9�N���ג} d��B���$�heAC[�{�I	��Ӳ; Ƴh+$�X�� >�^��S��f���C5���������A�� ������"#�ZYitܽYc���p=�٘�>�SU�}ڀi��N�b��s�(�1U>��l�*Gߋ/1=����}G��q	ɯ^T��LNڤ�����8��]���� BK�T��4>d:�&N٨&6�1���;��ux��t�}���IǴ������|1�@�� ��1�w2O~.��eT���3[F�8;�?�t���+�oX�����t��nK�]��X��k��b�A�_�r'j GP5!���q���%HP��J1I�̼�W]_�Q��>S�)W;�q;i��&�U�}=c���J¼���٤�aٽ��)�C��0֜��P�^(!� ��}�#�8o;�U�p�1��h{k/0Z0�Q����>sc|��n�㹹�`$g£�2�#71/�5UȒ5�^V4^ |6sOB���E�swW{o�k��O$��p
!>��Q��Vv�����ݯ;c_ �ȷ8�m��7�<(�c�������W��e'T1e��Ӟ�-�nXY=6��*�Y�����b��0;9�娜$��:{_a|�:�R6?-sU���Y�[�N�����lE��>�}�	�[�9o�#r��wZ`�ܱ_��)5�>%��P�x�=��	s����LV$`&~vO*��9�@��I�6W�`������s��J�%r�ɇ!=.Y�5�y'%�[�i�dF�#�f�i8�w� �y®p�����4ITRWOd=���\U��=^#���LG�Ym;R�k�))9�T����T6̂��\�I�j��ɜCA&��ʑ�g�!Uq�Akzw" d��|2�'y��R�~�����@����@�03w���Ђ<#�wb�Plcb�J����ar�$��AHK���< �P��A<#k���y7<z̯���h#k���q2�r>��R*�pX�����Bc2�{�h2��͇��#���^��ȈSF�����)�4C�<8�z����aCPî��a��3�П�����3�	QO�PH�aH5��V�o2Fq��H������gF��<�'\ �y+�9�T�v���)q�洎��)t *�c�w٤��6E�*;���MCwF!�6Vvs6CǄlq�m*ܚxʸ�;�4�^v��{���n��Z�CJz�x��+�T�.�š��%��������#�|;��� )<�5�h�QV��2�6�4�#��A/StU0�U9Ƒ}�|$鐓,	��L�P���g�xtf�۹�����]U}�89M�nk�h9�Py���&���6}]�;Y7�C���8�KL�g1/���]%�j��С{7���@U٪�gJ\�y��s��A�K�Q>�[(am�'��d��j$݀�F�Y홀���ܓ׉��L΅��0������̕�4Q<t�i��%�����;�^�K=+~E��'��W�Ԃ��L��l�-�ǿ��'�BQ��@�PF|�n�)�nh#]YB���p�[����B��G3�a�Z�2XM��O�߇��1����j�:EM���x�~u;)�<��=(�<��9B���5�3a
�W �Xz�9͎Sw�F��e��7�[�Q>�:yj��������c�ܚ���x�@��7^�p���{[-�+����j/�V�@���|�������!T?V�x
e��V�'Zg>�'�]Ѝ2�g�dлt�]���)��'�N״1�U��C���ڷS�ʜ���
e`U�v�����%��wl\X�2D�k�x��
�ˢ���$��F�#���i�R�:��D�׃i#t�`�"�å���~iei�H��ְ�f���`$BUS�)_,%.Py)� gE��E�7�ka���G-�N'����j) �ֵ �V��b���R�70Q����ש��^@ �3菆�H5��b��Bj��I\۹����l��1�J~b�4�9����ub�����q��s�/i�����M o�C~��ox���/�����Л&�?̵M_3 5 I4��)��m%��6iO�&�ha�B��w/?��΋��vX�����3C�F�.N�o�3 ��ێ1�����;ow�U��Φy���J���=�?W#sD�nV�q):K�A��"����t2����v��ծ��uU�;�㽸���d�0��!��P9f��1*�>�3"�"d�Ǟ��i��������3_=�+�?�+}�IT��@jj9(�Z��vD�/� j��P-_H�2�gvtL��s�	���)�~�X����e���j�#���oWtrpP��u�-����7�r������i����D
��SXh'�p�������r�S9�����?�zak� ���.&_�F������Vӣr#�46V��hΊ5����K/2���#��������~���8?���$�r�HG�	�s�Ӽ�3g��0O&��i?%|��t�
/AX����D��ϱ� �W?4G�η���3�-hk$��tBM�*���b<3/�)�vn��k�"тq�-)��C�&�/���gQ_�=��W9�+ZQ���<X5���a���"ij�G��}���mr�=��}����!�Ĩ26����&q�X�NM��-g�������5��}��ټ�Lp��j��T-ZZ�T9H��*1�s���WK�)�*��SY�Q@�?ef�]Dձ�m����2g���:��������1�Bc���?>�(�e�Oݓ̿T^F��>d$�.mR��C�A�ȹ�!��]˴������E�u,�˝��%��v��-��K�MOK��8a����٢��%���_%>�.��Y�§���31������g�~1�w	�:ܔc6�,��s�ia<����d��*4��-�@�X�Z���t1�9טlR �y}3�E�d���<Dr^ao$�_�^��(!Pg�?��q�/<k��w;)n<��a��_{�ZĚ>��:�V�$���|���H�;-����%��x1�l��}���������&~��r�8C�g-G�ua3ƝW�Fu}a�fh�A{źq9m�^�	��|r��S�G�6���͚� ��݉��m�%���-�g�:��2�v��X� �{N@I
��3�%�!4�8��ǃ�vL	|�
��	h8���x��-�vuݪIH�D}$25/=ݶ����,$cl�n��ɗ,g��N 0���b4�!&�0���{X-���z}���|�N�� }�޾%6�RCJ�5��r٢�Ƚ�WЎ�[>r\
��m� T ���2�c:�5��c����D���!窺��q7:�w�7\���w\he��F,��fvݍ�ޓ�:�����N��.����M�~	����|��h��������N���o�lA���Ý����S�n'd"S��v�C|?r�o�uW)Q�,���E��U�ÃC����N|��$��a|Ңb3��2[t�^��t�[��/"Y���6�.Hrʋ� ������~{��ܭ�1R���X�n�c�%�f�KuP8��U�m�C�2�U��|���q��yJ+N��% ��|h�B�i+�{`d}��p;�Ȕ�\7O�MQ�i�1S�\\b�T�^G�rC����6���w?�����_��xʃ�����Z���^uP7�8b"�lF�g��������`ę��K����Ly��݉�2*��ub�Ӹ��{�'q��Hii�c����eTl $~���IM�e �����ES?��p�u�������Q���a֐��h#8���8�]VuGa$xPlK�� ���H��{�I$�p�,b45�Cϭ5�9Cٲ{0�!�bJ��p$�CQ����V�6v�r�n���d O� *����{�����3��3�X6��%���L"�����+V�viҝ�g�Y`��T?��@��_Ld�d�Qg4���I���0`Z�#�i�x�1X����Y� a��ő�Pp���I�l���B�Cs���V޻��ըҫN*<Z�	��
���'�NM�+�ʲn!�CB^>y�O*6Ʌً�tJz�B<��\��\��o�H�l�oy`�&o�2呕\AQ;'�����PU��ي�$��k���v&�T���� ��(�B&9� �s� .fA+(�E@�H>��Be5�;�28g��-M)L�*�&q6�XFE�׵8��E�&���s�WUNˏ�T�Ϣ7���Z�����,F�OWg�r�VF��\5Қ���cX�yA1�;A�[���rj�P ۈ�q�m��Lz�� ��mT^�N��������ܣA�&<�C�5ťtן�#嚊υ*r#����[?�eS�Z�����HK��ݺ���{|N��-5�~��L���%�mb<����9\��|�(�����hǮ=]����e��m��,�؇nE��8���m��bM�5Gܽ�Yu��Q�NE�$7���o����̀�Zy]�虯|u�ȵ�fЖ�X��[�?��TS�� #Ė�Et�T�9�$'^?�l��\�a�w��GӼ�Y����$[��!�L����n�N�u5�X��80���Ý,,��I���zs�:�cM�B�#I��V1�,�A��ΰ�b�w�΃+I�z$#�6�.E;/�y���� �n$�h��r^��Z~�ƾ�y{��^x��F8;��~���<z%ip��Q�<�b��8ۂ�#��.��@�����s3�OA���tT���9&68>�h.����U�!'������7l	V9���.y|V�N��`=���zT��}m����Bn��I>m���������j4~�������Z7`ꔔ�����>�W˥��|L3H���� 9���_���v���9do[1��)P��/c���4uz�x�/�g!I>1�_��m�
Ӎbk�uĺ7qk���Ptʧ=�Aq�_L�A?�,�i�e$�c��ƙx�ܟn��Վ���\��ꫪ��w�oUy�"m��c�8�;�/��-c��.h�:?|tw�'a�����'R��ة@�NQc�X�vЉw{��|	��� q�����u�>۴U�B^��+0$8Cqܜ']�1���5��v�#+���3� .F0��]Բ���j �/�ឿ-3=V���э�q��� r�`ȶ�&��e�Ǻ��fdM��I)��p�Rߋ ���K�ky��b��)���Y��ƶ��\��:st�;�S�%�%8��Z���#wO��d��/�Pڽ^��G�D�X�0S�Uw�����2a�Ý(лM�0&C&sR��������u3 �������HF�ڱ��}eP�؜�1�t��&[�<�2�>���!���x�����LXR�`������՞��Z;��`�\�U�^�PM9L,�<"D0vk�,m0谁��I�#S�T�굳Ѩ��V�2���I5j�_���iHp�����U�o��NG]��O���}q����y�'�H=w��#-�
�o�j�D���p~g���&2��w�tw�bn��g-�`K�\Z�<]�������%��8.l�o���+�8-`�=��n!+O�!�4gMB;s��?9	+x0��+�klŔ���?}~�,U�+Sg�e8�/	X��f9��'� C� �S��l�.Xp7I�̄����ج%�"7�c�����nY�%7�c�%�� �W�ڏTp�y/��/�ht��$�G�=�8+��>S��8�dP��]�{� "��?~Y�V��'d��[���~�{������yͳ�0l�g�2�*&Q��7xӲy�؀�7w�$ K�[�ڋH)�V)�IVe��tvw�v�	����Q�-�T]u����
�Y��Y�U�2��?
���~�8-<�Jhx&��;�f G��""{�z�` ��հ��k���%����Q4݅�G����=����Q��~�483�Ęg�6%�ʆu1�;Q�[�@���(�=�p����+_�1ߢH�u('T�#s= �8ʳ&��;3H�\"h ��׳��]3_��1/��>K�(�����&Za�s��r��K�Ҹ8�\ѥ�i.��ZP甈����V�=.�y���~�����c>��1����	�P������M�N�C��	 �k�$�y��~�fF*�V��6Yi&�Y��}'���D�Ϭk`�K|d��6U���T�زh>Qۚ��ˎ���p���s��P@�]r-�t��4nx��^ډp��-�F��f�HL1iڛ�[U�Wʇ���{��&g���6=�k��[Rg��:�VG�P�Z�4H���ϋ�>\��z�|�R�p�;�ddd����$K~�Z~)����z��3�D�5#sX9)IlP�ư4ccJmRU'͋-�*bԉ�@�4u�"N��B��n�.Ѭ|�i@��:��jJ=4R��ߘ a�,�&�q�vY��jtc�,��&{��*R�Bg�j *-3��OT'�"L��?��c7���^D�`螐I>��������u{��8-��Q����F1��gqyK;o���\y�@քG0.~t�{e�,��,��: �o�S��ͥ����{ܿ�x����zz�N�3�TɄ����sWI}T5�}Y�����kh,cr��t����F��!���,���L���%㠤���m�0L�����M��|ʙAG(4�]����n/��������!���j�,�m�b��31�J]�vl/F��Sǃ�ɝ��B�7�#��O�NTj�cM"[�����z7��>cza�}�t}7�����{W�}Ź��_!hALX�fڽ����[E��.�uy�S��T̨��$"����a��y���ڱB�f�,��}�ظ2�FE������sp�_YނA����w����9e������� �0uo�x��KS�F��"P���܊x�b���X�cBT|:ZGh��$ ն�1�?Ih����ƒ�p	��� p�י�\�R�"��#��%}_��A��נ�
��M�b\��P�w��_ O��(yR�m�����EH��'�LL��a��^�0j�Y�2�6�&r�������6�hQT3��ߨ�1�7	�"�K��E5Ҿ)��sHd�oU���Qo�����ʡ�n�>�i��7$]���bR�F�H�����?�#�'���~��|��H��^BUo�h��5ٕ=�k�V�o����⩒������bV�7#��yN�0���6���чK���"奭)��ٚp��U��_�i5X1�����f�y�s�V�4��/2G��ޗ��>�Ck<��ZV�j��{Oޔ�k�@k;-���{���	\k"�-dDt�q�77r�#r
{M�l=-�~��ń�'�y�(��e�b���e6��J���gO�P<Q�ג��E���Vd�oQ�fÏ�%b�;��>ձTO?`�AN�ŕZ]�&6�E�������&R��KS��I��5���o0D��3�p�94����Z��NeӮ�_����[��Hi�v�2;��e�Aq�ǁ�0&��8����	/��tz�8�>5u6�r[�"0��"�c%�e��O�O�]7�����_�(��>��QIV6�~�.Ʈ��L4tIƄP������Rm9�����H�7�������0��K,e���-�ZaEpm�?%id���B5;�H2Y��'�&̏�n}�]C��qڐCz���D�q��;m�%=�<�&W�}�gwo+C�Kӓ���y��YB4_<z����;�����ߢӭ�Z��Ɵ�Y���z��p�\�m�$Ы��D62�N*�,z�T�Rj{I�˧9��Mti2�,-����td#HI�����t%P$�ذ�F.v�jD����Z��ڷ��j����$��eNkv�䀹��L���#
���mBQ��o�Z�]޴�Ѿ�n+�4¨�lu�D V�rzS�*�����h#vQ��i�xքxP�XQ$��4\�|N�p�e�:�4(�j`�>,��t�W�ʼ<�]�x��1����"��ͬ�ɄΒ4�s�a	؜&�vX��G����}.��|Ⱦ�*� o�(��3bƉM�,I&�ӧ:'��4$|%B�D�k�.xP�-͢��O&V�	g)ԟ�E�&P���l��!���9b_1�n�L��r�ndcL\�E�(p�����D�s����k���.X�%)�bae18M�vԙ�SZN�j�*�/�S�q��*%E��B@!ZO�r�K�L��Ut$��Ț ������P:��D(	ÿ�2y	C��|�*��݀M��y���9�Y}����C����ɛK���j}����f�SӨn�ņ*�֪�=�x:�	���{�;�Z,N��`�~N_�{��eDB�*Ê���S v�3��6s�5���8�(�Ѵ��I�3)�(f�Ћ��s���V�'���9�ĕ~$l��!@�(��X3܄-؁�#���QX?�f�&���ڒ�V�ݿ%�_I���Ӈ$��Xc[��\@Ǽfz�cLx���Z��P���������m1�U~|1x��v� F���1sBL/��0��X����}<*�P
���r��\�8`�v��Fj��֔o7]�D���d<�Xl`F�����GK�w��%��?�@����p�>�7K�a����:p��O`oU.u���ּ�ў�?�zR�8	���=:���f�Z�s쉄/����>�d���|4uk~a*�=���A���hH]���?I��� �����s��2t1�m�_yy�0��F��ώO8�a8N'�9�������)oeWxY�n��*��������o[�Th���E�r*BG��!�@����=�(c$��Sp`6T9�ؤ�=k2{j��I���/�v[�e+�&oMn�F��������*	�I݀����H f��NW�+��XcԡE�<[����>:��uVʓ�1���^�[��� ��j���
�߸>�_���K����<rr��Z���E�d�ʨ�y������a��L-h�e�������ׇPyW]�Y4��o&T䂭Ĉ�7�bY�Gu��:%q�NP�s�ۼz��n�US�[qL��D���R�]َ[ϙ���oa���π%�Q�
�N �e ���РU9���Zf��:����`��~�%�N��Emv-���wԢ%4�����������=B^���X]V�ɷ h#����rP	� &v.�k亙ؚ�@���v��!�^�"*�j�+��b�'�9�a��6���;h��
[Yik;E���1�w'�]����c@8''��I~����M�)��k�}�9k��	A�C��ɶ��i!-���-5&��u���!�po��$����Zs�x���2��׊�ͭ⩙���;�L>w���x@����r[#��ۀ���׋(�th��|԰՝IŤ#�c�,?����߿�諝i��Ѝ_�|�G��ʈ��� ������B�t.���i�I)\�d�*��F7Q�s�����L&��^\M�2� �<�L���t՘��Qc��}��-��J'��M�N���B�/�u#B�Jը��//5���Cri����m����j¥��6V�q!�SlAG.S:�z�V��M�����'�Q�%i���x�]"#*Jӽ�Qʽi��;�Jo��U���j�Gن���4Q�:���a����T`�n�}�΃XPc!��o�." (�"sXO�32��+*T�)r�0r��qF�E�~�H�t�*5�]
�u�b8M򔍕Ԣ������X��/���I�!����AUvX�ٺ�xљ�?�1J<!��P����,��#R~]��5�j�����O.\�&%
$/��O5^�.������3Q��t��Mw6�|e�۾(�6�taC�_��껾&�1�q�B�0A{�Ι�k���3s�ǜ��`)���qc�È\�&��M{rqS�Thj�'�������;�~��$|��
mC5��h���67��r�� P�}x��!uL�!�(�	��,*�;' �3w�}�?v>�ˀ��*D����n�[R;:"c+���Ѿ��3W,��$��hvq	�(�5��Ϣ�wf�y�t$T`���m��:z�1tuV��2=�z�v�#	�$�P	�-/����e(",ݯ1Kt�܏g�G�FRAZ���T���1��Q�o��C�p��Î3���{���?.Ϟ)�Ȓ�R��e�Z�DKj���\�xJ�
�HW��V�}7ږ��VH���A�A�ͻP�����m�d�����RU�D��i@~()*���������4@��s�sd��h�1T��a�Z�t��}c�����z����5~DI:
A7@���݃A�զ}�k���'ift������Ƅ��o%5�&���F)֓��'���x5���k���PR�r�/��TP�.��V���_ ?�[y	sk���"�Yh��>�aq�_r���0�B̬UK�"��.8J�Y�i�0Q%r��5�Pa�S��}�Abaɹ��!Ǐ���w�_�ZT��76�Ќ<5)U�q7�L륰I胇���U-�{��"E�1��B��(� ^�)@�(zN;d�����1�L�u`W(B����=������1*m�_.t8�}���v
�g�w=��^[ ���y����H�����Pmf0�+o" 4z1RN ��97P*x�;��u��t.�!���m��ԙ��5��@�5S��&uT��h���?piL��¸�ƽunF_M����1Q��G��O�St 4��Q�O*�L#�S��r;��{�h�	�pm3�k�x�$j�]B�o�҄m����^)�����7єh��zd�.�Rte}���_�fѺg��lםs�oN(0�Kq���B��8sz�v�\�-��!O��I2�����x���
���p;�>��P��P4o/����^���5~vL�"�oe��	�Ǭ%R�2�9�Hó���e����D��7��坯F�Q��\�R��}E�p��*���J�%���{��+#j����}���F�3��88�8��3��"p:k@,�ȓC'M��7�\F\��z<�!��)M�1����"E�Ũ���(�*��; >�A]�]��J�D�ᬇ��C��d�EQ�`X��߂�ڑ�?J�I��ma�>�:�H�g�Um�}5g]l�w��L-|������P,�$#���cL��;�⌄��|����0UNv��Ð����)�#+h$x�傿�FIhB����d2�4m�.��q�(01~�c|����o'�O<�
ml[Lc���&��ܭF���>�JM�?� Ζ�9��D�3<nH,S��z�-�Ս��Ey�(�?C�^�C�d1R�L���<z�T4���{�Ř����M�x�)�)8Z��8��	r!��)g��	���Vdа/��%�}/�(��&5��U��aNh<.����e�A_f��mq&-�ո�%�JY�N�'YNJ�� xw&�%Aw�p!5�@�&<�+�C7��꣹��vF�Õ�WD]���7S�7��il/TQr�9svC9=�E��&�kl4�r�!�I��*�HB��6�y~tY3�zЯ�G|�2ܤ"sV�Uq�nL��T@�Ъ���f�m�TJ�c�$��^�4���Q��[���5h}�K_8:�t����d$cO���kև�͚Z�^�4�D���Eb�;^�v�jW�Ҍ�� A}dTS^��׊U�`,v� I�/�0�c�9LD�\�����#���]��=%/����9�fw$�ӍY�V��|0Zg��#��9���6��3��τaʬ��dg�g_�jщ�[�&2�W��&�. _��aM�U`���ػ�+D.F�@ý��f��e���E;��՜��1u-.�x$��A]�<��<�����e ����T]I�9�n޲HӔ�$H��i8�-.H�{O�(g�z�_��YB�\��Cl�(c�������w�?J�z�e����\�+x�q���2�����c9L����r���K�ǭ�����nM����١}-R�c_06�X|��'K�_J��@t��zD��;���j�-���I!ؔ�1�A�t�����h���Cu���,���®^��nC���KI�ԅZ�!�#�����46~�3h����w��N>^3�s�r�*��q��+Jvz���H͛@�T�5;����P�$��!f�&ΤAL(�AGpH�0���m��("烶���`��_�NfS���b�DP�g�Q���2�v~� ��k`9�!⹠]DL�4)�i����E�l�����w��qӷ#����q ZU`_O�0K?�Ä�ިE��V;F
(Ųл��?�ĕ��T;A��Pm;�S!Ɩat�%�����\9����i��P��	�i�۞}��ɋ��b�8�[�N:�BcW�'�ܾ�S�[$"C����a-�s��;+&E�t���N~�]�;��L�}M�3��#���L���[OT��b0�e��d'�������`!������Ȁ�c��#��x�aX��D���a}�g�`z�ݟ����wKi�Rݥ�J�\
���-iϼ��XH�4-?���:��J�a��@�TI��mNy$�l<X�g�0(� V�#3�Q���8��y2���pu��ѯQ�t���f�O�G(Ί�;fG�>��v�T��c�\���@>��H�At�q��'9F]-ȇ��7?����zk�tP9��a�r�"���M)l8��	>(��":����k���O��uPQ�)�z�(�p�#� �Q�$��fXq�w-S��8w�����������(or��S���V)�;y���g<,gojV�nP4j��0-mҐ�����	����L��Q�q������*ct�
�����u��nq�������xY��ŐPU�U�(�Ch�*)�)Z�<N��d�t۟��"e�o��5՚5[pk��wF2f�ѓ�a}��[�h��U����QW�:D�"�e\UE�U��{#��b��o�R���e�K#�ӧ��g�^����@���Ӊ("��7L̢ݣ�/f?_kA-�< H��,BI�����hc��=Y�R���?���<�U+���d��K�N70%}ɪM��}�@49岍;V�Ys�4�������?!�.�7��xY�L2�qfOΪu����F�[��|��"��o�:q���ϱk崪x&k=3n�s�3NF~�8��v`kz��3Ta��,Ɣ_���'�e_�[g�
��t��t���Yuh�y�N+�4^&+��ꪖ����׭���K��+0��ui��A��㞫	h�!EO�ň���A�<���G�z"���+j�T㇓��=I�K
a����c�z�W�r����v5P����U�圤50�߬Ѭ��N��t�{�b%������?�6�(O�ɧON��l�v�؞k��g�ָ_�f���NN)�z��%xyD����pb�+�G�]g���(1*�=�������E����r���-ǘZT����ԝ�K���z���̃s�T��&=����>�Y >f��D�����]��6#��q���a���	�]�E�[����tF�.4�\��o@�_㈓��� �1�v�:��%�k �}�Z?Ta����th���U�-؄�U��z!�Uh��4���;-J�2��i57�Qz8�0�;m4�;�ί��4�W/B��0�|�@������Ȩ&��f'~���6���jG��ӄ��c�Y��H�������gՠ;���@v*�sK{�C��[���e�7�n�߄� g�L�67�wW�,�#�H�EoA.�	b��8*�0l���P�����JdAݦ�0�E��PG�=��b@BƸg.Q̦�q�qc�����=���ْE3QA�V�W���Z��ī�yw���	����ᛣ�4H0����N����r�a�V3�V����Yf~J�"P@ebotE�8�0mw�J�mG8 j�C\*��_��KB�q����Ȝ�j*�O��l���2�fx�6�˔|�g�8�-� 
3�N���?��I���������+������0֜F[ȅFO�w�Sѹ~ ���k��nLԑ�]�A����|���j�zg���ϧ&��J.�
��& ����R#N��
�kc8�;n=j��ZB���kqLf��<���,yo��Ⱥ�]2�Un8CvCn\��"^�	���-�g���k��3��y *'q'Dذ�)j��V2�{р�}��Sa֗=��'��=i�/��׉���� )�s}�F��!(X��0���6#����#FMF�e%|�.�d�D��s���&�A@ѹ�/��+�9���1ي���܌b�^!��|ϲ�V;�j�G��@�ߩ�oԶ�&oK�S�,<d�cg ����t ������U5����&�.Q���<GB7���>Q���<xŖ��=!�&��������S�0d%����z-hS��S�o���~�CRQ�#Fg� x�mO��_�ŅY���f��6Щf�m�w�KW�ùa�;Z��౔�����p��GoL����N��tH<j=w!E�+���ܝ
�^���.Yw�kdj�^� ��6*j6�"L3�d]RM��	 /�#,bn���u�ZCr$w�B�Q�<��X^�(E���dIz?�<��+��+5���2T���DF��х�;�Ȏ pքb�Vu;u���3�ʫ V�x p�#�~���d���t�CT�&be����|Br�-	) ��ͱnm��Hf�(����|�k�7�延�M�2X��p�E9=#�(>,
��m�E�%�_�%�~�lo�J�J/�Q�Ao��k�%�%,�������u�EY?O4�o~��-���D
�!m�e�^bƕ��$Ot�n�h�\�&����Ƈ�#%�yG�xWs���������.���h�6K����K)�eތ��V��Or�?9�N�P(�	�ٸ3bśd��=������2��\�Λ�,sX듓Uܳ7ρ��p�'7��{�k��������P�Mi��I[*�X!�7Em ;~��l�)��ĆNy]�?���z�o>i]�:�'e�]�:�%���\i^��R֟��Nv(�"Q����".�ͧV�]R><aoY��H�#f]ȓ�[\� ���U���=�p�^��<�͘�^�=>�-�IT:=c�ࢅ,jNP���u�A��q�C_��(J��?��a�J�D2����@@�`�{�ڍ%��-��rX�$�]�����]��̇@q�R�8)�D~���8��+ �>�H�?��|�;���Lk�l�ܻz}�֜A�C��H��S�٧?���ػy�-��VL#p�.�%�_!q�zp���i�f+a�]�r�={��jE8"�K�9q朲;���5�S�ps�oY�����J���"O�M�^�Ҽi�Sm��^���e'cJ���5o���EZa�v�g�ݸ�URu�y�+4�� �.m�,�`T�r��E�����(��t�3  %/����<�����q͗��
��D�}�U �	��H?���s����S�Z�"O�?|#��(�&!��J\m*DgU�S���Z �m:ܥ��V�m.�?�����7� '�.1
?��dKؗ̾U�F����"I���x��2��r��F�w�]ha���bϙ�lX� \�?>���@�Qmq��<�j�ċ^��bq�8�;��Kh-�Z��:�Ԅ��<�1���߾x=�V�O�OF�%��7u�aȂҢW��7�$��8��.�^�(z��ڸ{ތ3�̢��k�rE�����6x_��v�h���#D���=��Q`���#�W��Y�]�Y�mE�D�'��Eޒ�n��X�j����$���JJz�����Do�����.��-��1�o�}�}�B)o�>���y�q�K�5/�'d�$�N�����Y���8N6W�
���,Y5:P�����$�mR:P�U�W��p��Ƀ�Ue�K]{��f�t{w�߉�#E@�X[��Dn72�!�oG�Ǥ���3�8,��	���)�ÚtZyw{l��ڽ(��.&�bV�e2���
S�嗬=�����-|��D��lL��i���)�'O�����!��10�_"Y�W��s"~��jZn�v_��G���Wf��EK�6y�D�g���q\`l�n��� 6ӗ~iwi5�*�jb���,]��*�OSΔ!{��5��2���D���֓:�Y�����"rk	��9��9Ǭ7D;ّ�$�1hen[Z��R�@��j�}�.��s�Y�
�_�(���ҩ��92�ƨ�I�{7�o��]�s�~��3�ʘm�9���/}�&}y������)�=���N���=��%刿�Ckb�d��Վζ0�'`k�� �A���\��רY����_�Ub���	Gl�/�Ō8�C�=$��0"Ԉ����Ql������jN�3�Gi)�Ȑm�IZ���/w~]7�p��z��=��>t�$�mT�n�G?�����>d���'�]>�\'�k�D�8-�e�L�8Z���\F!�������޺`wD��7�"{��$�.yT�	'�l���ԡF�G�y�/�m<�g6�itO�o7��S�+%$g:������"2}��d�XmZ� >ݺ=Y^�
% &
�LU�J�� d�=���GB`0�x�+P�_��9n�mZ�kj�(RT�"ըK,d�߱��������'-/�&K��<�H��rOH�K����\����Bm��Iz��][&¾L_�'�&��a���:�'���.޻D����E�j#,u�(�9lUl �T�$�6N
�������-�6�<;{��ȯ��}���J:5Ŷł7ꝣ��"C��JK�����w�=��*���PY̑���4�<�x�#�ڜr��d�IA� ;8����d"��$��w�*�⑯РoD�9}ވK㖴އb�����|{��<4�btKk����3�4�jc��n��/�KX���v]��fn����C�VY$�����/h�ڽL���B�÷$�I�{>���r��U>��>xO���l�;��T������{�����-��������vV�G=SE�f?*	����l�k��k	P(�X�7%�lk�,�#�bS�5�Fa3��#�o�̸�s���q��P��l�h܄[���^��b�p��ټq,�&}V�/)=�����:j�TF�>��v����z+�fj /��Z����hW�	���ynL���X��@'|�>{瓼ݚ��'T�C����|s[�s�{�Ji�ڼ�9�Xb�۹lf,��q8l��eJ'��J��ӽ\�6P9A!`�!�b���PC�0E�,ЦZ!R[s��eњ�;#0А&�n%ƗK���j���,MKf�ޒ�b�H�8fr�뮳S��v3�n�A0�8��g?a{�.���`΢�%��`��9��� �N&MZ� .�mw��f>RWuxsG���?p�@I o���7����|n;L�	�:�9�<N���ѝ��;�b�Ѣ0	�H��᳨�U�	t�b5ߣ���k�{�$>����֚O��݂P�y]�?�/g�,�=^���Q�쀃�� �=g�xz�������x�B�O&7�㺈d)�a$6tm�:�ւ�V�����!��5}OjC+��Voc����d��FR�Z&U�s0�����Z�`�"�b�J�sV�.�>��=�2�h�8,��B��C��c�q��8.��f�B�����KR�xsm�f!�;&��nث븨�ZX��D �Y��g����7&CS�����7Y�"������݃���E���7����
0D�>���ɑ�bީ��_����
;f�*z+fu>���[��6�լ; �W
�ҳ"�o��G��c�B�J�_e�8��ɽ\̷6y�<��v���\�>g�ҳ���#'ԁf��к|����G"kb��,'N�d�����f9��n_:�X��[����뚆J��4����vC}9�?��Rqt��텅��7g�W�E̓q>�yg!7B%mm��e܋��g�3�O��4|p��?1ӻ�c�1Y�v��p���ϋx+D�9J�Foʥ�'~��:�)K� ���dE�r�e���Q�)J�x�:C��m4�%K)�8����`�(A��� � p�tLN���*Uf<:�Hq?�(rJ�ʇt��m/EJ���J����^�e�+���!g�����J�7�����I�:��=_�=2h$���X�� �W:Ti�")R������*�y
�]T9Kru���oA�b��,2��B�`�ns�����O7x�	�d��e�	`�$���9'���Cw�Y2�p&����]�G2Ԝf��<�VW99�0���p�>!�ݗ3�eq�q�����(~R0��60���>3�QeiS�v�[hE��;����}5(:�T^j"�R�ψ�ǽnyd��(T���H1G>�[�u�.�����3^��F���0Q5�m,5K���hd�τ����w�ldP��I�j5�<Q�:K^ �>�����0�I���n�xg�n=B�t���%;<֙�NC�B��Nz�`����:�j�#��ܑ���;Y�I�ZeJ��������B�s"�"?�I�*���+\�P�	�vPW� v7��X[%Y��t!��ڮ
;����R�{9����7�"����N�۳���T[�]^c����y/�LPrZF�0���$7���o���ae�Ś�W{칍�y��]k�,�7/��ݟۚ��7�H3(�S'(`��0fe|Bt䯂��\����w�'��^��D�@b���I�D��V�|�*0#~�m�m�vg�Y�����́�&v�=����՟��Y��m�.�a��780$����]x�VP�$B��M�v�̬���R�gg��^D��;�ۻ`t���������d`�"E�����qGMZ7+����B��$vS86܈�0�fU>0I����c{{q�L������[1�*�. @�;/өR]h-��E���4���o\'[KM@x�<QJ��r\j��y2���b�e��,�����-�S�@G��	�	9y�T�^[_S?f���t�Q8�J�r�-���L�6��%n��PQ�]	��a�����3�CF���Y�h������?mj�4˭�i��3n�׹p���vf_r��M@!�Px@*O+�*8�B�k�T��LI�-r$n͟�l������hT"Hwc۹I^�L�U���e�$KR�)�VO��VLFj̼�Z-����?U����S<geN��b����+<��4d�K)�����P#��L���R����ɢ�7l�z�j?��h%���2�-��s<r.�i��[w�����(mٮ6&,5��� 7�W�sn���J�m��J}͠=}�o���}��� �}�pW���]!�Vx��`�g�J�?�� ��^�=�������
嬢���6!;xn��7� �3{����9u�J���qj�K��>ᴭ�/n����Q������y�s�CS�3dU6�&�Q��6�?�/u�FS�#������g�|��6҇��;�]!J�p{y��2Qr5�r�yd�QZ[���S츈cS�m�����U3�"���R����}=0��<kS���I�����Ӂ��뢴����0%�����+�K��W{K�P��z������Ga3�n۪�0�(�8�c0��B���t/����s�K�fJ%-^�p~%H�\W��ݧe��o��8�O��W�F:��Z���˟���v0����Wf��I��-�N.*�[��|��A��C]f3rIHۛ]i��]��w�"�=�:'�ēhǰ)�b8� mj[xp�����-B^�f=�����Q'm]Cj�+��E��}�v����^�
��A
'�\
×��@ʐ�ea�M�w��,r�vV���56/S&3�<C��&�R�$�noŕb��P"}��r"���pO�	��9lqE.���>��g��`e�D����P�&�a�L�m�>������c^��yH�����li�=��&t����OE�GB9Q�7��g9�� �lr�=%��䁘���!&eoYz��i�k�ɹ뜆(�m3��Hz�f�����J����#�?����?bp�~��~�Hh�������P�d2���!���7*�:Ũ���r�k:Q
��/{tx�&
^L��}r��WC���bIP�aX��!a�HE��|��P�%9�V0d��� ��Y9��&�J�l$�5�'��I��uc,�z�+ǧ�=:��,�C�x�:9�����]j�_o.��R�#)'�3݃� �]E���G<\�$d?}�:��ɻ��ċ��,j{����U�ڋU]l�(m:�����4�i5�4P7ۜ�A�b�*`����T������C� ���I�gѐ\���K˭~C�ְ�7�<�
E��%H��4-������B��8���/����п8��\��jی��g�	�Ġ�ak$�M+O�k�EE�M�>T��fi��J!��4Hl�AHa	�XfXZݠ�|?)�]g̣��a��k����pN�67���;d�b	�|���⤯C�Z�A�T}2ϒ٘4)������B���?%������J����;���)�(���ތ��o�:6��2���5�2Q��mZ��%7hA����  ��(�V�E��7�/���ݖsP{�6`?�zvJ�Y������rS�NBJ�� w�%��c��'�ᜫQR�` �,e����3iAc�?�4�L�����Ì�(�-�	+���}�<��`��í��~	�m�����KJ
�8������^R,"a9x�=&���i:˛��6k1��ۓ���<��y��}�y>���g������
I&�f�ab�����t�
��&��U�biO��D�]tR2��X����f��r���V��w�֔z42�P9.
����� 
�U�	����3%�J��Ѝ�co�����K���M��r��H[R��ɜ\E'4x��>������\��a��cm��,���P����8�V�6N�:����$%��`�1��sn8 q�˯�v�V*��������{�2E��[��e�j������;�]Hl�]g?ߛ��X���r��;�e�%Y�q�Ф���tW����!�J��`�8������7���=)�$|�����ob����W@�.s�Xj�Ew/���_6܏r�ݧ�T��t�sXA6�m�0��)�L=_=��a��k�+1������ ����{f��#�6�o�
�s���Q�--R��(�X|W�U�G���MZ���k�GR�vo���b5:*��P���"���߁�YL�q�q�͗�It��n�'�6]��f�E��9'����0���w}F!�xj�3{��r&�e���4Y��UZ�⌞�p����P4�O*����{�O�"��:q�D��D�[��o��,�w���L ;��h:��+�9�2����˅\���s-HF�­��4!��}�/��v��G 
D�L�����!t~+6#n�|��SglZmpXv�B�\�-����q�S��f�#~{R���N��D�|q8�ꅕ'��c<.{���{��K�e���-g����$�:�\%l�<(6��Ҧߜ����C��%ݨ?��#�0�tRk�ҍ�)wp�RX���� o��C��>�)qe��*!d�* �ӯTq�s�uG�W��	���L��fY�2�������-�R��q��P��}�ߔ�0�`W&D _R�3�RУ�V��AF%F!2�Ē�y�:�e*�x����(>~f"�f%��@�����:������=�Mc��{��qb��g�2��
��mh�DM�`z #5�ĭ�h�sq�	hu`<1�_�ү�^h� jBhEg�� [�i�瘲i���5�H��d�c���XmNx��)�8��&=�^j��oq�uP�z'0!������8�Y2t� T%�s!O2�?��L��jӭ�|ׯ��RΒ�q���~]�М:��R�S-����'��#�EY��0��{K6��\�5�hܶI�\�U�K�8V/��U	% ��dA��#)QG�8/Ѥ� ! R�Gp���}`�$�\6�8�i�R�?�?E�s��4=t�>N��L9#���K!�x�F��@������wHT-l|�9��8�!�v�q�ϜZ�%'E&v:��gծ:�h �rZ����V�,|��S�;{,�ݎ)�I����bјt$��EÀ�]F_xuī��1gTy�YgI��
�����W<n�$���<��	�㩵��_.�� a���B}�:����,��lU��~�>��T:ŷ�ibES�cfv��|�J�q� Iu�Մ~/�8C�{f��flg�'�c���lb(�k�R�JM����
��s�}����Yx����̺Mm�ƞ1���9e�(���/�^���)(�MZ�>c�j��
s��e'/�Gq��V��E�qO������y��&WRѬ"z�����ku�!l0>�POkŪ�p�03c�Ml���7-���ol_�e���h�t�W�Z�+��j��\_�W��}|ouo1���.V`ُ>T��<+��$�I�1���=�FU�s������Bh#e��V1.����~���b�ފ�,�h�_�=������i���`I�}���?"A��7=p'k�ZX9D��b�ېn
�@KsuC�@��s�}J�;G�gm��qm��ZN���N����s� �Щ!�e��$z��HN牻�h/�Rߊ#2p
JfgB�c�"�;S��ƹ�M@�8UH��ݟ�H��@6�2=���R��`�)���1p*z��5�Fa�Z7���L#QZq���� eCw<&503p���mlE}�����D��_ΐ�B]K=x�?�˧�~T���@(=���G�M�>�#v��-
�uWRM��ҋ$]��>����\R��WQ��������1�s^��~�R�@֌������t��U�/�)�)�k�4��z.��T<����̊
U��]`K5����"�x��BQ�ں��i�Ż�����hw��Vz����J@Er�J���}Wbi�B�w�-1'����o`�k��64��.p>�ui�i��{������e��!�Ƽ�^	ˁ|sQ�L6�́Z{�@ݎ\�X� FNG����h~BGiU펤�wR/k��Cl����R��UP�
o˰�E��,i�ı����LG�:���k��P�9��^I�J��o�Na4q�U9(╅8y�E4�lv.����q^\8U��.}����ӷ�}�r1�T�;3�dL���Lf�gr���悭K�t�{�l�9ߑ*�vq�l#%Z�6ͧې$]�L�:�q�qv�}$��y\�%v!��QC�!R��7rI*�� ��ǵ����
'� h)��M�����
06o��θ�tE��O.�͞��sr�2J6�r�ĂKbV�sU!o��͛R&�E��>]�%��f`/�i
������^.�i���*B�$3� ]a�i|o�"l�;�j9���sIL�{�U��c�����S����^�8-��2�ݺ
z_.�������J+��C^E����#vH�H��"}W��S�'3�I��`���,�s_�Hw��.��#c�=���
����"�*���h
 ��B1�%T��ftEI�'���L�1k�b ';u��,n���ͭ��%�8�� P�	��$�e$QV�C$@Y�Ę����2��53q��:�ju�����k��&�[�	���_�^e����ZL�ؑ��Wt6*����-B!�@�
�('�a���0�׃v�8���n�!W}�X�_��o1&���'��!����}!`�c 	���<�9�����d_�?7�_R�xu�`�7�K~�C�sW�7���F8��Բ��㷨������A1^|b�ת�HCB��j��棳����ܚ�o	m7A��>���J�{u�% �!W�߱�hĲ^�ᶨ��tu�M�>�9�r�y�o���_Ĩ�i��Uy5�2n��S�?uv�z	"c|��z��>"5�<�]3�M���:�k�c�s'�Hr��p)���˶cg<�L�Kq�H�����@$�+j��F<n|o�Odoɀ�
,�t���$
+w��o�.5�S��-Y���"�eN�`lϯ�c}��%:�J�� �bu���Ñ���*��<SA���������8y`�zn>��v1�ئ��X!ž�H�4���w�Y�6-�xl��4}�|�` #
�o��9m(�����~���2�f3ylr�vo���'��H�ƉJ툥8�w�jiP��*�an\�����G�V�H&nC	��3��H���b���ki��/�lx����ݾD}��ہ����e�*�}6�T~4�!.�u�gǛf�봢����)�NQW�>���-r ��)�o�A{�"��Sggq�M�`���o�:,��2�a��¢!b�<G��Q�Z���GD���|]�C/��I���f�ˤ��W	��.�bag�1	!oJqLO,e�6t�	T72��x��x���@L8p�E�d�x ���z�@�^l�Qa�Ī���������_�W�O��ZƺZ��r�ȏ�3Q��3��9J(q|���m�����ЅJx�z�@b3 *q������|�Yӵ���������<"�ygX�(\��t����TD눍��Y��$��$]�ESm'O[Dp�2�!���juϨL)��Οg�������0ۄf���O�]N���JdNѪ��Lu��Z�-�7�B�qq��@5�Nd�<k�{�h��x�*�S���j��d.v��Jt6� 4�N��ώ�`˭Hv�2������k	�P�;����V����-��L���V�X���j@�t$�G;`�#�����H�k�K5�����5o��4�N�$��1eF��x�>�����:��e	�!�Aꦋ@�6܁Z5&P��r��Y]$��c�x|��xX�]Ջ6��@{}�W��&od���zI��nܓ�k<�E�����^��Tk��s��'Չz�3B�7F�p� D�O����T�K1��b7\:P��0%��@��a���y|��x��%�	[����I���,���ėg���z]�0���O�oW�����m�txV�q�õne�mV4?����_PAb���>����H�����r��*�ވ�b����y�Ba͠�I�u܍��y�D��cZ��`�^�&`�	�-B2fS�ZH�e$���� 
���|K��7�<�A�ވ�o��%�K��|e��{�H���7L�)E^�A$�2Oi�c�4�>��x�{c�7�U�%6R��_���2�����;�9�2���{�P��U�S�^�4���?PEV�X��6��1Ӯ�(�<;��
 �Y���*d�}��Rx�_��A��K�i��S����j���p���f���Bl��TIJl%0a���^Ϟ�3di1]|�Y+y�����o.P[}�l2�f~%���L
4�t�Q�~V���l�������r�e$f��tQ�\�&8���ֿE�r��PV���S���c�m7���bL�@�ȿQ�����R���nt�ٳ{f���,�+#`?7]������Ɉ<]��L��n 5UFd�rQ��cx&���:�q?�+��iz���J�C����,��4��7��nS���Y����5k>�`u^��w�H;�C%D��*��u�����l%�Ɂ��Q7���K�gb��8�f��瞶�Ƅ���Q8������A�`�;2Z�۳bs��\]�>Q�*��I���Z�ΎI��)N���F,�ʀ�BP���~V�!I�<��r4}�@�p
��4�16�X�86,�6R��Ƞ+�����.�TA�Y �3���U<>�Fl�����i=�.p9�B�z$��TU^oV7���N/�1��o*j6���Hu ��HI��7� Eg�J��Ә�.ftU�����q���Pd�@��)K�P��f���H"2��! r��9{��.��S��w< ��ǢCJ��(3�4E��C�&H�|-�5<��៳�OP�w�Բ,��|dfK�8�l�ĚtF��2���f�6�W�e-㛍]�Uj���(����U� �֌���Ē��G4����~��&	�ړю�U�Ԟ�#�؜�y
�n�S��Q��#@5d	�@m��@Ҥ�ׅ�@�^=b�?A{�>�W��AumZ���D�)M����\?�<��'Gl��㜾�nͪ�Æ�B[�O\n%'�@�����x��Og¾
��cV�E��J��M������ .G���AdA��aYQ_��ڭ���<�j䯣�#C������#R19�nl޶�����F?N"��쨢���Y��y����;oZ�
�wl������4v�xR�%�ɝ��u7�%�{ʐ!U]px.�XD_3�2�d��Xs`�d�wƓk��u���ԁ�A"Ի��C�=;��}�2�/�>��/���y}0SPe�Z��U�О���*g^�A"�C-�r�~?8OYz��p�����3:��2�>�������_y�~�żҩjB&}�_l1�����;�,�	 �d������`0����%���V��kx��b4d��>d'���Xԝ����/A+�L�֙ Xg�{E����@����QL[�=N�̙U�KP�ˮ��7��/H��k"���S,\-=s[�_*���^�\ʖ��\6�����V�deD`Rð�C-
2�{��\۹��ZaE �{����]/.*y�	�_9E�W~Ut2vfª�r^.�晀�L�TuC���3$X*RK��SPIO��2 ��Q�u�R�,�Q���������.1��S�c�sZ�w���p�@#l"ѹ��3�[��|�.cqI.�o�/������v:g���A�q0U�	�+�'.�w b<j�jt��Y��l�6�s��ĊJs�����1�?�t�6�"�#����o����wB�P�,U�eͰH����)��(�D���zY��}/y��A���Q:c\�������bѻ_�\��h73bbN�9�nI�B17�5{bq������-�p�R�][�n-�)5hEO��+:�=��PL��)���1�瘽�c�J>�s��h�ȤM�7��Ғ�W�X�&f��Ԍ~�|@�}�_��4L�]I���S*���C% �4��r���ix���0L��h�]���T�}0��a�N���nZwf"�eē�Q�C��-�e�]ү�!{�}f���_rQ4Y�V{uڤ�U;��7ٟF�������
�3���;��X�Lͨn,�*��Pd�eH�9����%�������l�����B�SlYX��J����~�tԤ�O-�ּ���8�w�P(r�=ߕx�Fc(1�s��v��tH!�K��|X��I���-��r�BA�ka�d�/��f�O
�A-�f`�qg4���1иu9)S����o,�*�Ӏ���-