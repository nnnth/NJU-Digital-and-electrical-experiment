��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��c����"3�p�7��,�j�gvì#Y�+b����W
�j��{�6B<��~�=7���c���qAG�V��l�^��k�}[+n轄k���2����%n )ie�Hc�k-���gpKU��g��-1�5l;�,��g�ʳ��}��d�P^^�ڕϳ�Gʞ�5�ќ�Z%��l��C����I�mI�A���N�	�?y^^׹Z=A��祐w0������#�Y��+�ϲXJ��PW���j�;��&�dp��1�{M�~���q��ż���O����l��6/1ĸ�V_B2Rs�y��^�37!!���� ޔ&}�-��r���T2��[(\y�_Ad��p���9L��AL�5�ڐ�l��u%�q�6U�iu|�J��U���iG����ԕPZ�:��Ԅu�;/\�dZ�vV�|s��+��G�r7ǿ��m%�_�4V$�Ɓpoab��f%�Zm=3�$�X��B���\h��� �Q��1x�!�d�3j"���r�qIu��HO@#/����ä�m���,��8j+c��F�6r�$��Ju��m*�W��
����{�tB���_�x1dgƅ�F����/�{2>�}f00w�s_#Q�����Jȹ7���?�����.ϐp�g�������B�5b�'��.���\������~-n��5� &l$�ds���Nk��\pOI�nbc:E�$��t�m3���V�Adj����d�!��Z1H��#}u��'h����hYJ��6�(pÕ@�����d�5X ��AdC8+� �SKj* ���z̍7�B��3��ķ�L# �Uܫ���z��KΖ�+WF�_�2�=
���q������6�4`[,��~oV���	QS��f-�t
���f(M	�W��E�7��m�L�P�6k;�MH�*Akۅ�H��U�o3YE<[km���[�~ņ���l��J"lر8}��>{4������¼��i�������'��3�y�] ���݂��Ds��g��b�'IK�����nK���[T�c��]mN3���v�ZPvo+��*�l@�Wc#�g4�KD���w%�3a�5bo�[����o�I�AK���}\	抣�U�=L�7���ɰ�'�%з	���!r�)�57��I�{��f@e����4a�4fן^��^_kU��gc�������(�8��ʤw�X(�r����X���HU�藸�J0\^a_,`�q�x s�̃�Enydt_��F���$d�㻪����͸偭`�p葈���g�К�w�F`$��J����;w�u��sk(�"g8Ya�xk�N�b+��\�+Џ y��u���I��;?I�=�ԥb粄O�>|��]Onީ�
�._B��!��N呲�.��S-C�5,=_�?E�	��R�0�з���_�����݌��LC�%辳(ح��*@�y-��W:�x��挽0�sZ���mR�����#�4[���Oi�E��ZO��M&W��g�_N����,���j���N�SRRF�^�K'�5�<�g����bA��m=9L��m~a�gR��H]��-r���P'�љ"��*� ]�V�&�0�3X�S%*	Z���x���.���W�o�e�y�>�)��4�4��S!�@2a�c��bn�w� K_u����c�e�U[Er�D�8�hY�G�|�W�gI������?��8���>�Te�P��v:���R�.S�����<~�� #�8���77��0�Э}5�:�,Q���j_n"��W��;1���s��iya��Sۓ�T�-����&���2k,&=|i|����v������z�(k�D�����h�1��푲2�Y)E��	�k)Ug��Ð�:�Krg�1ꖪ{,j2��`y��<t�~��%��S��7*
Z$t����O͔�#X⽏7�j�>Ɋg�C,��T��:�����%n��|�Rb��'{A�(�������#d{�7�{�8�k3��i��,�ϵ�f%w�Z��2	���S�3��6��O7�,�i;�:8 ^�$�ᜇ�/V�>�F�O�>�z�~�������,���)��[��-�-�)����;��U�v����C�2����.|q�Ph��h���Όn9{-���������_�Q%��Tw������'S���.��@ێ��I�V���򣽡�Q�=!�:/�<)���mw�$�B�_�Dd��"�}^L\M��2?ܷZ��x�����n�aU;��ܰ�N`ȳ1�\�����vԦ������NF���&����%�������Bg�t�$7����C��M���9�|�B~o�4x��:V[D|��7C���!�d���r&���o�͝����z`ϲ��⇦L~Hg�%�;��?����px4)���u��|�o�]A��-�vC��<dh�黐�C�Ӹ_@�V��}��:�~g��q�*T�&��G�O.�zA�>Vs?q�6�-�a�Ë�t�p��D{��ƴ���Ii����hB�^ꠂ|�ٯfZD��'�x�ct��?�^���X���a���]�M�{_̝R �P-G�6�bo�S�傴	i��5
�C�!oZ�M���
�0��\�|ߎWǫF��KɨF�u?7�㹊P�c�!����h�j�@�	�![����c��Lz������TwT� �2�[�34P����+F;�ލ>Z���_:h4'FP�MD��:��O�H�5�,�	�E�K���	W04\���L���jS�J����2��?�9�Ɲ�#N��f�|]�ܔ���`Y� ��mNd�v�y_�b\l�9�g��Ϥǒ���]<j�f��{Q�l�D[�k�*��
!��MN
����II�|�f ಷ��7�j�%�Al�[�r���*Я��q����|����<�����J4������+�'�8Pz9~��~si)��էI�����[afb�̻����
�ӄ���<��.��S�}��s���C)ǜ�3����C>�Jg8'�����(�.M �Uq
_f:��?�� ����x�h����uu�{�5���o��l|Fb�����*�r�]Tal�}��Y�����/��ٻ�������1�g,+?TUR���r��e��R@�k{�jq5��eԍ�*�@��8�}%n8h.Հ� ���=�?�/^�+�m���) Ԛmo���{sG��}��BU��1��R�D�߫�\��΁��w�Ycd2�2%u`ii*q���E/m��9���`��,�μ��ԛ��q+��?�$q<���=�MЙ���]S+��j�����Q��gE���SC&�
�v1#F|Ӥ�N�6��~z�~�I��\��)�+D�2��� �?&�@vj��՜Y*^�Ɩ��	y�e�@)� ���\B1�=L�Si�
�!�|e�N���
�pG{^�k�~�9k�Bd^���s@���5ɜ<b��(��踍��=!�!ͥ�n�{�S�n��}[�{q*M��ф%*�%�5�4�d�++ؗ+�Y���(�x1��0�Hf��0�]�©Վ�`Z��fsq/M��w���"T�� r�;ٖ$�}J$@Y�j�w5����oR�'x����Re�G�e���AdB9U��}\�b���"E�:�a1��A�B��6�X.S���8���W_��ƪ\�=H|c>K�����#Cb9��CΌ�͡�'�'�\��n��W���=8���H'�k�۟�Fl\�۸E�^o�H7�_Lh�@N@�w��L�v���.�u |��a�M)�\����RʎP�+�UD]���A�^a�W��.�9_����C4rI�r����@S��2��ވ%D����ݹQU�9���$t�N*,��fJ�[�>���@6Y���mM�!�%0&����V;e*pà��
e[D�qb��u�Zh+y�Z�GO�(���	����|��R,|R���E�[��	DL{Π��r� ���)BU:j���������Nܻ�Ƶ%@����tHl���,�K��\�?[��-�0��n�'Yr��f8�zr�˯�>�L�u1�iW���ߣ��ܭ����I^��ȼ��|_5��{��li��l��|�6������ɻ�cƗ�w�
Qy�(F�6]w�dxE&6iȐ�:�}�AL��7�|lː����%{�p.RIm�Y����z�_e��T���F(hN����G^x,!�����T���{�Mr���X"�nǝ�y�xӆ���eхcw��W$A��}͌�������i���·�!O4*)�/�z�������TP�m�N���_1�s$�0��'~����dQ�o���ާFrl}�}z݉�yN]L8U�J4��ҤmI�ô,���ig\��)��B�3�s��Q"(8���7� ���,�y����Հ>����dĝ)(mK�]�V��I���]���s�k�ZG�ͻ�.�T��!j�ogN<�����`��]Ǻ�ѣ��n)�E,��D�\'�1�t= `���~Y
\g�\����Yڗ����?dyU��z�[�B·�	��ɻ����5��%֍�m�
�
��i,�]xD�RV����c�dgC��rhf0�l��qIQ����1õ�c�~��_��^�MeX�5LP~�~�~��{�IWcf�/p��M�Ս�͟�6�H}�ܠ/k���_���&ǵ���b�����UJpX�so��u]���Q��B�A9�����GJ(��YN�d�6�;�J礪���<C���X-�a�ҭl�[�M�1\�Q:t��:�ȳFF���-ghD�p���j���{�{�4�%ZcY�jd��a����ْ���lj���[t2�.�-��������k��a)��k<6�|��QS�y����T�_����&P�!hcɾ�{���^����ڕ�-�V�	n�<f:7W#7-d����nb�� �`��b���r<؆�"�B�>��m�i�ᅚ���0�"|��YJ% ����@[ɈE0�$��"K�f�\��K������|����cE��s�I�U�Fb���hy:;��1�N��)5�_�����h¾��/����S�K>� �u6���⛺(���L ���U�宬�텉�`YR�WJ7�T��1y4<��b"Q��8���%C?��q��ϐa4��m�/�`�ɼ�����(�&y'D�w:�^��q�g�SW�˴���)O\�@�vN ���teHm7���I�r,)�ٛ���꺂&�(x�ܚ%�EKq�Ŷ�sc1x��\�P�����NkD9{��
��ٸQ�3a1�]7��\M��z��u�B�Z�ƅ�`��}��34cV�E����;��K�Z�'��J<{�R����O�&�'���N|�p�m������(�E��к>�
ǁ�;5��,{�J�B]�"��>Bhc�2�f��� ���N���� scNZ$�׳�#��Uy�"HP���Y@�+�@���ڄ!a�f�F(�X4���3EBq0x��;7���T_���e������-�j�h����m~ˊIC��������i�~z޹f��2�Rz�Wt�ħBL��HZĬ���3N����Բn��I��#גc]y��o
}"�{[@InW<VR|@v�j�LIz�_���y��7P��;�3cq�Dk*J �N�i��X+�$f�НE�lZ�l��}i��^pV���.��tĨ
��ژ�Ɨɤ���,T0@N*}�<�S�J��~1�_��p�B�/�r&�W�1
��/i|��\�e��a4X���K�TZ���o�ȳp�>�r<}���E�4U��� 6��~�$�@c"�X9��ݽ׏�N-�8`��v�'%/�P�%H'���:��G�1�98��Omދ_�떹���.o��-�<��GAsO�2n'R�����1�,��W�����A1�w:�O�w�p,e�Y����g'|��ޚ��7ݨ��Cr���q���k(��*���L��?J]�����ڿE�a��i��S��+��-'nt��p�4~�͇}2[�@ݕ���.+p�:Ա�	~}�D�tU�1�d��8�n����=���3��b2��Q+�إiz8��AR��K�bPZ��L�u�F!�7�Ipqp���U5� �Ւ7�j'�:wVU������W�=@��ݲ�]�:V�`���G�L���?�d��
�n�ZG}�,>qh������Ԍ�@�S�ui����!�ES������埅Uy���c�ձ7ɴ��Bwi�ҵǜ�;��1��0�pH��r��h\aM��[Y�+m�@���eN`h�c�U��o�bXbbަ	��W9��k����k����i��zs���)=��XPI)[�� to�����}x���"{w�u�ʅ6�C���3Q�YN
��~�x����K��
� W�ދcI�q' )���O�cc��z�"|~
�P�}�?�X+#8���1~-�٠Z�1�}�� �*��7úJ�|�/�O��.�{����=�ԃ�:d���a��S����<�JW�cBLru���Uk��:��&�������*|6s���=o.���[>�'Z�c�����3�}�zFQ���!T�'�����%����%t�S-�T& J���(��Nn���������j�)�O�i�����>�ӏ���R|�D<�s�ʬ�$�l�:ax7%6����'�<�C�\��Ǌ�H�TD^K����������䩋��w�Hh��q�������M��pF�]�(�L]me<��`\����dp|����?��Dۦ��̏8�@N��9k�t�3]���Y1^@���`�,��)ɷc����O�x��FN�q|�+��v�n�}��K
�
��p�aca�D_��Z%~3YN*�M���ѥ|�p��q"�L���!����%�]r ��@{/���j`�x�˽�n�lj��.%��-��7z	����5+e��=�ŵ�Yl�v����slgj�z$ʑ"���&WC-���ӌ���nF�g}~0DC2�2��)��w�9��H&T�u��=��5^���m�\��s�Orf�6nϛk1��fmm�9�_���dG�ëYG��؛b�ٹmX�dh51��D��D�5��	ɫ0Y������˶��"��;0|�.Z� \��b�����GX�B34�SH��y�>u�{ �{Z��ё��[:v]���-��R�8�oB�z �a�R����!�[mեO�sO���jgzk{y�h�Yx+ F$=5�Oy%��w�s�֖�a�p'��0�����D�2`T������5���l�0E`���*�ȺӰ��ح�w��e��%|�LN~"0�\V�?�<����u�bb���L* 6���]�e�"���Bw�x�E1A�)�8(�q��
L��V��]��5�
���1�2�p_W�-o$��[�CFy%-�c��:<��NG"O�S�P49��Ys���*O����cea@�0[y���'�px83��2�C.`���Q�kI�	��6��A� ¡0f�쳼n*ȇl�	0��LȂe�j�u�r�81۵�q	�5q�OѡD�Ha���:���*VO»j�-�@��GbUɋ�=��{���nh��/0�o�F�ض*bX,+,�Kf�������Kɋ�WuG^�XWFL�����L����O[~�)�0-M=`.���P�2��{�7���XLF`���`��Q�N�,'�I�抴
��b�,;��Y��s�����vՄ"��S�|����
���㵙��C*�A��9�3�xW���6��=�*�L�
��([����ͪ�+�0�^�����?
u���n�;�zJ.� <�Q��������ӽ�S6�/馅��ڈ&|W�i���I�S}h��Q���r��܎����ڥ�e�s+9��~�,��*J:����������Ԃ��V���5rm�pϿt@���4���)�d�$1�a�{Ge����eW];����y56�L���]<��RF��ۿ��,��Q�sŖd��
�Z�����V̍m6��͇�ܦ�^�yС,�|�J���N��d�M�E�tda��AF������S��S��#�։K.��I�r�{)�[���T�[?�i��.�"_����Za_��<NJ��bk�e�c��Ǣ~*�-.z:��+h����kKc%�9�_cs�F	�ה�fç�F�}G��-�LHt�fGː��Py��bOzI�W0_��t�p��,�]bq�c2L��|���)����{�Ϋ�k�cA!Ɏy��?4�����e9�|�[+��TM-��F�W���xLgڞ*����x�L[�o͑W�=�]�ش���²	l��`�� ��*�ˬ�����>�@+/��RQ/x�]�����A����U���ۢ���@w�H���d�Uⷸ�
�WD-�w�U^��WD��C�0�-��S)���}�C!$�O�W����"(9yN�<&_�<	Mx��5W��m���m^Z��Oй^ܔ%1������Üq�.c2_�@p�Qג��4�w�~jr�ّ��96�܎�lKtzR6��J9���@�Uq���q_��
@MIB�EŰ���:6M&`Pt�JC������<�9@�` 6kaZ�%C����F���{��/S}��aB��n��DUT��r�x��K��p.��-�1�f�j������=m~�ط��`�2\����'��gQ	���]�~Z��VH�Z?�+m�տ
�Wmt2qf����Vic9L�,;���^q��7F
a�
E���m���=b���' 8L[�	�E�=(� ��8{�
�zҎL��9�S���.i�j�ɷ�c�nE��6f2��.�q��Aj
�,g���Ȧ���w�x�#s(#��}������j��.j�rNK�	�X��t)�[�"4��Y��]쟅�'����Aِ1��j�������7�3�2c�����8H*X5�,޽��c�a�=n�?�A�]���i�TT��{�n�8w�F�("N!�x�k�L �ԐMϲ�RYoF��W�`�o�ʼ�����,��%���?���ڹY��Db����ѫ\0�s<���������vȽw�Ҧ�)|�Y
E��,J_��")f�կ�����"��*��KR~��'5��/�{�*�e��I� 
�{���s~������k���Y>E2g&��9̥\`�*�f�~H2h��n>���C�<���b��<'����,�ۄiPA�)�^<9����iQg�h�H���9��}�/�"�x@K�8"�����࠰�B|�~ V,�R�8����ݕL��h �ݔR��a�2sL���rЙ�����5<h��C�0�^��Y*��I��0�k�XuR� ��,��D.�ﰱ<����#9� w�G5��M��ޥ��L�>I<"Ĺ�t���C��GO���$٘R=Ȁ���㍍O=��ɬև�������&&�5p�VO�驟)KR���qS�eC��A�.z_i��%p��7_����/J$e��FO�`1�fF���u�@���+0+{$i$�6�b����%l���1��!y��R!B��"uX�s���q���p�Jܔ>��ڣ�%�!�R?���ʸ�
����$��^�����|�ǼYl��,�
Jt(?��Ri����0V`��f���,�=�j��1�85�k��K�@�T&Z�%4�K�r�*�(��d�q� z�e*�h����
�A(O�y#Z�?���ⱊII�o���!��F��z��ZC�E��Q������{ckɡ��\��eB>����!�R(��#����#���[y�f?S����7X]��1�))�r ��'�&��v�LR�"E��ʃ��s	\��sh�]&��$)L�Y��l�ϻ9-��h���՟��m�'F߱|o�s:u���_M���'�c���M��:��Yx�!Lkh��e~����:��4��}4)�����afqw{����A��o����Uu*e����V<�VW�W�Ii�Õ��E����ii�>�#
����#]��S$L��W���9�fM=ϛV����7�L�p��i�(ڙ����5�i�:y�ֹB���xNX��~�⺾^dju��K
U$ū�V^�IȚW��T���ŉ�E�7�#��>�Smo�3Rf&Lة\u�α@���mjdX�cgg�����e�z
d�O\4�D� Xhf:A���	�s����`�K��%�m^b�� �r�?�Ge�y�6��&F*#*)%q��휮}ZYP �ᾂ�U��t�L���a�5 �h2N������V�'����
<��1�m#�]��M�̀���q��J�i1޽4
˓R��<p�q���n�v\�9N�<�S�/�]՘��o�¦�߉kX��K�'RQ�`[��Z8?���+*PƜ��D��ձi�'�F �錾�(98r#�r)�+�>(9��?j|4����n-���'�ˍ�P��pdK�?Qg�}D.}	C���i{����L�n/�{:��od�i�LV��k��@���>�-#���x9��zv}%���b{����xQ�v׈��F��H#��9�Q9b9��C'�%����rMزl���Q�k������HAt�GS�z����xC˞C�5+�N��\N��&2ۙ���%�_��4仳��G�1D|%��n;w�f10����F@��?�W�P����]�6
�@סp7Z@��d$z�*h�8���:
?ʆ&�6�g��7�E�q���c*M/��%�~-Y���ʣ3".���)�2/��1r߁ҫ�V�n#K&�ѿ',�xYBE�`�2"����M��m����&�ہ�>��c&��I�����T�뱇��v�-��B��r͗��(��(�0�tǲ�H�ʂ4�Esӫu�C���2T�Kr��}���:�'l�Y쯫��BC�l�6�D'�kb��[[մ�[=>�<�r��q��/Fv[�gaڼO�\��	�ti�Q)��o��y���`��Qz���`Ӌ��T怛V���I��U�1�EK�!���Uk�}��qlm�m�6}JkSyl�О���)�ۡ+f�ŕ<я�<����Tߜɷ���+�
j2YjmC�%��Gr5��B���L���»X�-X�i�]~ڔ6y���F`�L\�vi��}����UF���b���'3�L���
noI;���[���6�]@��mCZջ���Gⱔ�p56Ɖ}jI�)�c4�1�=�s�Q[8b���0�G@�S���6qaA^#�V��m��Y"dL���JW~?.,c��cnϔ,I��x�^�EL�΀-�`{��`�V�F��ޫ3u�o�F�F�sŞZ��y�.7ۑ�*�C�^v�)��p$�6Z&/1P6t@>ګHM�҃D"*b����m6��s��G 5��`PU��`��I�qkM�3�W==(F�?⪘�Ds��� M'�%D�S�[��O;P�z��dW�$�u�E̖�}l�T��On�MۆD�9<�O�!�� z�aǓX���b!j�y����������Mg�����U�:�e\��[�'��j���2ߋ�f��� �5/1���`��e7�R�]��'[��(�����&��$r?�q��'#Y�������
����L�l���7+ȢK^?B#��4zc��
2���z���o�_�6/��朩H�7��%̋�F~0�)(�A�Ў?Ώ�̈́�Ԃ}�ujP�S>�.Uq�!$�-��#�oe�_�
�gK��]�}o��b�Y�\��ND#�p�_�
�-�����8��G���&)Om%x�R�_	����9�'��?v9����`8�9x�g�Y�N�����J��7}�&��P���t�(�H��X�O1�`	�QGˈ��Q�v��0��T��h\�,>C�r�z���8G���};�Ӱ��n z���H���-����6���M
�}3��/c>9D1H?JPx���q2$�b?�'��I���w@W�ZJ�d��N�B2v�k��Pb���~q��)�5l��,Lň��BjĐ.�������GGQ=�s�	��0؊�J��ݲ�ռ��RY��q��o�,����h�$:
C 
@���a�b�Ѷ~�Us{��@ٸ�i�9�/|�§e�*� �)�o�Zm�x�_O�)^n#�C��V���v� �zj��WC�+:�}����i~����Wc��2?���Z����Ӟe�3��詰Z��+�}����6�OyV{M�� �	�-���2eJ�4œ�����-y~�[G`�c�{��������P۞����&9��8Vԗ�n\?�yKf����5�E}������De�Vv�.	@h&�[֔U< �N�Q��eK�w�PGņ~�i�&;~�A9|��_u�aC׵\���]��	������z�|��~���7�w�T4N�#p%��Ur����rMKP��^w��V���x����7���#G�(M��e�Y�fI�1����2郞;�ަ�2�$����P�ˌ1��s��t|���@��~'Yڠ��V�����`��k M��j�~�c��}�q���%��|�@����x�x�Z�	�X-Ajٺ_m=x�CX9A��
�j:uA$�t�?޿�,�� �N�����9Yy ���J9n��Z6�uQ�S ��wZ�h+�a�E�\��*�����"�����:����K��m���ńJ��{W�]�!���Y��2uf�=��m �]|��`��`���-%�S�k���c��ʌ�(�y �֪̇b��$*�f�5M��V�E�"j�5�����@ձ[DZ��yrVj�y�T�\�>Z�+�jx[D��-�(��t��ǂןĈU�;�W���xid6�3���"���Ok4oY%ܱ�]Nb�= ��%<�	���kk�kHBV��~���Y,+b ʹ<w:����ڸ+�p����8���K��^/yr�!�4DuU�$z��Ai�e�GC
L��A�����( G������f��^�����L��0�,����S�@1�9y����[7oD�U��	�JR�<��m�`9���Cߣ�M��>�fe>�@�jRb�(D����vօ�v�ó���(��w�Z��eK�����w��f���}��Tn��U���e]�r��'AD~��z����2�ak$����1�s��ά ��Q�&�n|6�8�9�QC��R{=�艸Q�wc)I��N�����M�V�3���y�Pe�8/3��Q�#p�Ho�XI���E)0�̰�s�6�&{i�(�~��G׵�n<��7h(�u-���॥<Th��瞍���+
%�!O�﷚6���H�T.ItU�e(�)��W��v��̍:���[>L���a�x���X�{^hVp���uC�7E���+��Xn�c�.���Z-09< ��a�k*�D樺K^nD=�O�,����ÝS���4 �y'ii����s�o�!I��Ҵ��N7!�ٖ`f��[����I���U:V�I�_�8�r�2�v(��.2�w�hJ �}�M���Z�ە	]F��yAR�a�}�n_�0�2��uZS1ۢR�q�	Y�5D����� �0�Ýi#e
�>� D�ׁ^w��/n���߫�z'w�
Z`��)al=�z��|m(�לEZ�1�'����l散��Y1�`4Y`�����st���h&|�6tA�-�b�^Ɓ#f����i���d�܏���<�9��16$�1���.4�{�X_���X�z�!7)��.aM�S�CxW�@!�U����(�Y��o�ɛg)J�T��#��w���}��Z�X�����&�G��:�v4�=L8$<:'��Ӑ�� ��
{�����@YҪ8ѧ/���hs�j���P�/��.a��I9!-��&t�����4V�)X���L" } �{~ ]� {�����J�d.���c�L�5�~U^�3�"���x�__7�'qXJ�՝{(~�oA؎����Ç�ώ
?��Uea!|*d=�z�d�-�R(o<���ɫ�v�.�TMYb-��Xj/y����L���>�`o�� �媇x'�)C98b_�{o��5�O��G=5��.������AoeJf���)�:�ڙQ�,�S���hUN���w�|`��_ӛ�����܃o$��柔���ݫj��Ay%�G��t^�Cjb�u��`\�>wn.l^h���Ǫ3(�x�S�Eߑj��Y	�7���P���<|Ԟ�Pm� ]S��ߎX��+%����N?�Z��Q��Ϝ���:Ȳ8�6�s:��͝I,魚>�"�����y�=��	  n�����L+f2]33�Q�A(�*㐣1v[m�6[Ҙ`
i��(O��)�e�Qzy�8�3�g��~��gi�;ןr� �'T� ���S��S��+t�G$���'m�Z�GH����q}r�&��@1����;l<��"a�"�f�����ժ/�3?� f������W �]<�`;�o�X_�%l��G�Z���pGA$��zh�������a�X��n�P��KJ��!*_�1��+���*��TN_�9��G)!��
"ÿO�O8	H#��/3�٤7c�ʃ9��}�*9}�4C�*��Lw�2O2�W�����'b=;�C�Ob���?{�%rgS��k Ԓ�9��5b�ȃ��"L?�豬��&ڵ5]ۦ�W(Їu|v���G�\ERϤ�֯�̼1v�2����H�6��{ ٱ^�b���cD�f�@D}�X��Tԭ��<�&%HJ����T���Z�fP�J�&�RY������ɍ�S�[S��:��M+�U#[�lZ�hZ�ܻ��w7����^��_b�#��Ɲ�A���Da��,�\�r�KʯY^�����!N�O_�/�����:T�V�%�"bTW��Lk��y8s�9�WI�`	\�0�ɘ^��e(!-�b��H��0K����::�WO>�25%�� �w��T_U�է���IS��E�ZR)�L�!BU�q�M3^��"RW�˞;���#<�{(��$^$�,P���&�!,�/��o�Cx�vI�����$��~��z�	�Q0��R�����PJl�����7G���ㄌ��f�t(�~��n����E��D�E4�Qqk*���r�T}Vf} �VA�1�����9��`�������t���Z�΂/��@��	�� :*�uE�jJ;�wv�Xi�ܝB�O�2�C>��	�MA%K��eZBm($G$�B��0J�v�V�̟9������+�r;��{RT�"��F_���{<�@�&
 �yD0K��?5l��{m�Gi�9�HQ��-��Qߩ$xYδ��K�Y;���AZq�5w�K7���+�G1�Ltpʸ�g��rP-��.�kf�����/���BR]�[������?/�{�7��g^�QET�V��J��p�Ж߀�=���>���w�
�ӟ�|��%�N�@�iM�<Gp��)K*t�\|��T�N�V*+X��f�:9e0���̮��>}�V�/&���nEc�,���Z����.&�/�z�`��\���^mW�aGxT���WFc�\����|��8�fG�g����Z��Q��{�sv�K�F*~�=�q���B�/��k}�7�S�K���r�tIi�^X��v�����I`lYP�Tt.|���w�tJ��C�[ɖ����[��_[�@�Ma׬;
pThG$�) �B���Z��?����}�8@�9��C�������f�P�EUO�j�}��غ'�����K���W*�5ϝ`sR �=�:�q�'l��"�؟C�^ȹ��3Fj����;��@x)������ ��َa	6	�Q�b:J<-��h�����
L`r��^ӂ��.Ė��M1���.w�~�i��#�8!���M�x*o��a���`�����9Wu&���^=�j����N�@.ݽ�ˑ���@�ģ6^a ����`���ܑ��#;OJBmwC>�@`|6�?�5[l��,cQ������`[F�%b'I��M�~8m�e��W,
}�(>�n���=)r�ޏ�X������ ��QO�L{܄%�{[�ƠAm����s�O4n9�zuv+h�Yk>̅�x�rl���}H/��r��o)-��"&�z~�0�rz�`�n� ɷOVob���ƶ;���q����BigI����(����k�IphO���k�9��	�}&��6�����.-m�/�Y=l�<���� �	sU�MN�dd��P��6����eȡ"����Y 0���$���{��3Jb��������0/�x-1׫D%��yގfyd	���a9R�M�ѯ2�V�_�!��w4pܼ�|X(*�i�s)7i>w`4"�`�0����0TV�CGpEj�'���Qk1��EQ�$�)�8�4�ێ�jKA�-T���2N�*�m������2��<8��9�H4׆�J-qO�z�J^vz��T8�WO�,~������$v��55�)�\�{�k�t�Kʞ�z�^GFU��G]�u�c�k���_��]��d���`m�)�y� ��SK ����ä\ՠ�/�5�>i�s�/�C���Z����dl6�~�a��]O�6���2�m�M���XY�x�H�K((O9�ᯗ2"�������؞Iv�-��K��]2<�0��H_#�#��ۇ2�@mm�*�@R��(q��;����.~$��qU`����r�#��U�4BePƬsh��41�-�p����.�hul*n�#�C���{*B�&L9�Ɵ���z>��
g�r�bu���p�=q �z�Y#	�O���Č^"�KQ)e-/
Nn6�r�c4d��~�``� ��57D2�9�ܔFQ��\q����n
��JE$�?�B�LP0��,��P�tŐ�u�j��6��P�-5z#F��n,��>���V��PJ���z�e�*4�t��j\��+�ZA�<XJ���|+�.���bhz�m�cV `�N�T����>�a���Bt��Q�h}Z�z��p8Ok;�Q/�G��8���~��d)i�����$̋�)^]��So"��T	/օ�GU�;�"�u��)��e��n�E绑Eo��t�|*�?�G���8�
���e\߫�\�$���
U��t�gA3�h"nl���zJԪZ|F�ysфע��9skX����t����M����,w����+�������g��p`��Y�1P!��1�h�����#�D��/��_v7���(5U�q-`?�%��}�<QY{�GjR�Q� ev���ϝw��`�Ҏ'G���)A��:wr!ߗKj� �[�k�a>}åZ����"�|�Zk?6f�)��V.	���·;U\��R�Xћ�xɇ��n����Y*es7"�q���]�cK���#Q���4Ü��[����L� ���ձ�W|�D޸h��x���ѷ�
l>����b��S��Cލ�esB��i��S=F,�ޙ~�eu]�=��y��f�o]���@(�sf�޲��c�4�(F�g꾻%>t�.��^���F�Z7��w7!Y��/��{�O_kO�ǜ�m�\M�6�i��Z�UO�j�==����^�
��@]1wB(m-�Yȋ�f���$���=�ywQn�/6��o�����đaS\>�Q
�$с:R*D��yqZ@�r��V
Ц�M��$�?����ɳ��E��ܡ�*����
�ץ��@~���S�/ �N��X��VO��>�:��p��zv��U�A~[���D�\Үbk;�^���y��>���s�AZ�K��S��C*�G��ܘC�H���`W���뒙g&L�4��8\ˉ�Y]�>��Ǚ�\����?U{�Q����=��nv��f��~���%�2k�3r>o����e:N��S�_J1�d��R4����S�܃��JФ(U�S"���mk���I�)}���&�c�q�g�����J�ܣ	5�!M�:��U��8@XR,�J��Cr���R�q<����@�:��t?&B�"���	T�h�e�� �J'�Vwi����i�Q#R���٤L�[&��)����|2�I��K�a�\4�@�6�x�}����U>��A�Z[m�,�gb"Pfk�|����h���0j��[u��� �tQ��搕V�2��9�X//��ҲdJx��O��ER�W���>~��3��2��-��[:Q�~�F� *>��dNN�����x���>
g��z�p��Y�J.�b���95R!�1��o9J�i���2�|�����P7�����q���X�� ��>�H&N��ny~��Z<��I]�_�5):��r���:)��О�� ��H�eA��y��i�G3�m4+�,��ޡ���r(:��IkƼK���Ӟ�t=)�iSb�2�pa��3%�<��ъqD"С��n�?�c���#<;?������<�)�sjr�#Z�������>f�r&���$�A�S�_C�C�y����	�:��Augu�-ò�����A�����J��������>W��kT�e��;}�3�����u+�;�H�O!-�j�pz(��݉KYl\Z��T� �+�ۓOp���
/]��ƍ��j���zc�&���O��0ݍ���N��5�V�z�D
�Z̄ ���?�$T������6��5�c�c����&�>M q�Zn��X��`���B������ru�f]��n4U-W�����G�Q�I�>���LbvCK/��;��'��Ň��dK�af8^poNc|���=gP($	?�M���lޗ��r���R�7g��|E�25l���j���o��� ��k����M$A�=H,�|����t1Xw�vAb�0a��*J���(0
M��"s����8�X�rA~հ�BI�YlU�ĝ�>s��\�[ ܷiN���R��y��\��έp���?���A�5gJ�8�
�3�)9r���F	���2������ %�sݟ���_�3�76D��e�#dE3y�
��^wG��q��i$��W=]׭Q��ǁ3D1h�@՝r_"�+52kO����S��P
ނ�%{��I%W��VT���'d��w�Ԝ�ǟn�t}�����lT�@~D����� &E�^�N��ت�d�@012��l��D�/^]�Ҵ��{�D>[��t�����7�e��0���ו�w:�"�wX���̆��T�n��1~Y(8mz�,``o�C��^�>&ֿG=ffǫ�h���Ep���c	�&D@&�����ˮ0#Ի_�맃���Y��qxX'_
�����.D����,i�^���+�>�?Cs�����2��cZ׳iX1�1����=��X�9�#�(�T�#��+���T`�ב~1�p��'��x�h�l�b��;�Zי��.	O�K/7N��o�Au�$�w�' �Ւ"��#5�Kgg3UN(����)��0����.��k���|�b�N�<�N��B��>�ZBG{��sz�bjTIdʁ�mO�(-r=7\S�	R�9�w�9ڂjѐEFdG�U��+�R�-�jL��vrz�H���8	0ҍ������;���C����s	
8�;�%˽d�/i�AB|�E���ToH�{�B�H>��!tO�yֲU4X.GȊ�	����1<W�<|^g�:�Vr!Ȉ	u���a�����=�>q��HV��뼼��т��c �p�����G��4�\/���1G��n�	hK]�/�ˑi��_8��t��� �t�M5k� �G��Va�7Ơf�7��9�%L���S�%��f�^yeS�;Iw�@���UJ���^���=⣞�o��DPJ�p%���(Xh�ܕ)�׫��R��'�*�}������l �+s���S���� f�6$�CU�R�Q��gAu��k!S=s�V��Y~��[��`��W4��>��v�����iک��b��h�կ?,���;���N��k�G�ps	�,�1҃d�� iΒ����9,*t��r���~w��9�������.�qu���n2���e���CI�g�����]�,�u��$3��>��sH*�nR2��ųl(���
�qo
d���7b��k�:Q���H��G��9�r���8O�F� �����z+�R�ImK�8��aN���N��̢�!)���a�gtJ����z%B<ʪS\w&IcK��}����z�ɹ�@M�_+F�R��EX�Q���Ti[%y	�mx`ųT����x.2��G����K�j_h�l[�v�G��$ʼ��4A���fC��[���G�#�C����m�JԼ�*,�)�B6k*z�.n0�#f��%]�`�5CA��s[��1-���[*�qY� �W���AWK�#�}C_���2�0q!1LTɼ�h]�"/:[T�Gu��^��a7��UJ<g}��Ț6hHM�ݣD����3BR� �]亐��8~c[Bnk��3�U|i7,ɜO�8�]��}m4� ���.Dło�	���>��A��p/6|�K,�!3���3K.��"�F�}�.p�n���A[5]���/(2���m!9�!c�5��"w��韴��2a=����\���	k%Q���7H:�B��n3�O�R�~ɸ*�0;[�^�J���������f���@�'οR����e�gtڍf+1Um��pPq�6��+�[N�ٍ�y,�0�Q]�(pX�j��n�2I�������IB�v �C��B��9���IUMKs�[�g�y{���Դ����C{�a�/`�G��$��4b����b�ԞZ���M(Iѝ<���(��]�ѓ���?�b��%$��^�In�>2� ��}\��O��2���̖E�җ4y�������f�����@b1���|$v��X� Ӎ����� /~��$X����8}s���;�����>�aOҾ�Ʒ�Y�wD��&�f�#�G�1*Hڢ��E=58��Kz7uq�	,A�yR��dv��3��[�<�$~�~ܣ1�U4KM~ɏ3����
SF�*j&×���RH->��6�b�$������ iz�1�U�>��T*�?�:�Ӱ�<$��)���A�����C���C$�`$��w��T�Y
� iV����d#a:m�����zXhsVE� ��Y1zY�R��B����k��E@yO$�O����mKG��ʴJ�~u(~�mI2j���$,�\j����+�����4�ȴQ���O�-}Ώ8o�t�$:��B�ҍ��[���Q��N=��{��6�΃䉳�8A�����:<��n%Gc�D��.v�	o��7{+����n���i���+��-��n�\�k0ݝn��uA����	�`AKzq�n�����.��á�ax�<���Ku�!�I��w6��M�&s�^aq}ґ	D��R��a
�x���l �s|��@N�e�F(W(b`��YS�0jo�c"Ԙ�����9���Ծ�yb�*��cG��Y,�����a�qH&>�ֽ$���~�Ԭa}r�Vˤe/����oc�Q��	�t~<��N,�R
�'��i�ۆ|%�:7K��,a^��[�"�0n�|82�y��p�:��0�v ��j�V��G�c���pU���렯�*ǿ�n�	}�!r~j�:��Q[�C�j�n��G˂I�58�I34�\�� �H�|�ު&����-�$8P� :�<T���=˃[�o8��5�=�PiF��>�[d���'���yg���]�d������U9uL3,5�ȸ� ������c�1q�*�o�D��u�q�d�퇍�`��o���1P��� �YZ��7/ňYQa��Es���iH<���ݏ�S�qLng�����2� �]/�p?�LǄ�U��tw<V�(f�VʹMrL�<Wu��5�����S�t p,uWf3�����)���	wz�����ye!��LM1���+.�����L���{O�R8�w�H�)��T����;�Dy�&7g��L�7�V\�u�]n1�1[�ύNg�3r��L�	���|����u�_��^u��V�eH>\	���W�(H������Oj)��|A��	f��(<������&O��-㱒�9��&�XK�BN��q�@�t�'6�cHz�"�px����� ����C�`�D�Ë��w7�8V���Hk�j�²�{�5c���n����1$����ݧ���	ge����+��-r4������\h����o*���������8�\��9�C��ߔD�p�B���Y2p3��um$
uPpH��U'	��hɴg�SJ��j��<���0�e7� ,��\���Q;�
40��f����h���I�`��2��^�~{��'����(�u�w@.��e����5�'q�U�2+��at��TK�9�|��9�+l����kp�	��
Q��kJ�6�3�Q��K��g�2�C�>ǺS�y��f�Ti��К%9}����j�0ZZHV��\����ރoi��%@ڐ�ѺNC~��R 'pg��fJM��yCﰷ�t��p��W*��L��;jt���QWd����JQ~��U�!���j��U�}��x
��&��Z�$2��uwܰ��%ڴ���7���P��)��&�Xjzy������n���FZ4����Z搨|F%"�Z4s&j5O��"�7�?)(q+l�羉R�xGN���$f�{�/�,�wrL��P�㏡��m���FH��%��ن͔�p�A�A�cۮ��,��L���W����8��BH"=�(Z@Ԡ�Vho^�}l��MBZ)���h%��{>�b=��΍�h���+U�(�g,������{��㼷K�Άl
xg&��K�Ŗၳ �e{��8�ԝSp85AO�$H[e���ڀ���o4o�5X%��4c�
fѱN���I��&jm��Y�
�eO��8_������؏�/ph�a,���r�5�c&�88�X��1��V��r��ŉ��׺�G�2'7P��'�r��u�_��썌��,���3	;�
>�!h�����>&�/���j.w,k$Wކ�=�D��#�Za�j#�1��?&Pb�����>�X�p���tQ)}n��P���0�����[A>���s�h�v+�I~=|¢��iʊ㇓��V���}u���X��To�����/�y}�:Zl||K-�	��4~����D�W�<-L
�;2o��Y��&��F_���0��̗eu��_v�U�X�\��sl"���2wu��;��,�40�:
(,����(E���='�A=_K�DC���;�^��+���ǗK�1�OĐ���Æ`��������Dab�$i/rEVE�I&u�aC~�t��L�*�I���-!q	d^}�1�����6[�"��)SFo��x�
+#�q�J���|+�9>�<NO,����� \��:��fN�"%�u�٠gW=��Z+�l:�d�j�M�g�6���T��wױ��)Ȱ[	MO���hX1S8i�U�� ���م��N��SN�k|h�Tl����A6�]�:��W�:��i