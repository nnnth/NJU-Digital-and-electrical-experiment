��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�_���v��	����}���g�GH����U�K��*Ѓ�!N�=�Bb��w�����9���\�9d�I�S�D\��i�6����-�S�9�5x��
�hx�A���&m�F��K�]��lX��%��3�}����r]j��N߯*㾡'��|����tiN����H��7խ9k��-�l�m��DYk��B`QI���,��BJ�1э1z�:��sf�ch�	c�;�_s�5���U�?�t��6��&-G ��s�NHt�_�M�ܶ� �c_2\��1�s;D��&��9��'{w�g�s��ab؞������h�Xg8���2j� �!C'ǟ�A�)�ę9��pA������M�Ȩ����Q��	�U{Y�z�%���cY�X��ᅔZ���;�qo>y��%Ti��Qz��M4�JL��<ц:��?���Rjs�]:H��P�R�A4��6`����|f�x�K��f��K�����G�4"C���F����d��S�x���{je���{��ȽU��������S��J��1 v�7��.ް�?d����JN�c�}�D���g���Y ���u��=��Gtq�&3y �d���z6ؼ���{qz���*��u���f{�eEN�}3���7���O��S�8���F	��(GغW�D��Sh���_��'��V*�nK߉m�#�jOc6�e��N�6�(�)�Up85(fN�����Fފ��F�]�/(�C�e@�(Es�=�z?[��İ)|�i��˂��{L�|�ύ�Ți����5��86Q;�rb�.�r<��F}`�����Z�H�ji-���s�c�0��:��B#t�r���`+[?	�ߜ�e7fDݥ��e-U�	y�E~+�7a�㚥9=�Ѻ_l�4��j9� ��;���	nJ?���r~z('ᒞhn�,G 5��F�A׳����2�/����2�t;����Ln)��+xX��٭� q�^��^Tɉ�*�nbNN
�8�@���)��_*�����Vqw�<�㗺�kFL|b4��B��w�����˭���#�CGr�W�?�]}]"3��>���&_�=�=P�;�<�66a�Y��3:#������ ����n5���J���25��G��e2���B��k>�f*-��!n�UP�[�uY���ǑC�'GL��:hl�;�Q��=�(н��T̓��WJ�O.�
OvM}wB����T��"u��*������7� ��8@7m�S��Ĳ�e�ć��U3���Xc�*r+whS�����柖�ކD�L7�VT�TSDyUa����Fk�p�,�P�D�H$R �^R����*��7�����N�n�֯G����|<�'��/d@nzm�щ�(x�D���S	9#�.���O�$��h��n�\XM��0 ���n��:�Q���5G�֌���-:�C�jV#-4#�h�)I�S����Kb�Z�u�m�;�)V|y%�c�u�P;��B�s����}���b��ѽ�����y���5թ=A�O��_^�y/��ƚ����{�
��{��}�."�����<*�gwkYI��I�oH7��k���R6䰂h�9�F��ʴ��U	���ɨ�O.C�-eG�RB_�
d�wIŔ,=��m�]d·\��q+�!��ք:�h�5��&�>��.+�0�����DlS�'D�HF�A%<��Mf@��2*�FkG�S��}��#՜�z ԑ�I�֠�V!7��)?��<��Mpw��	b��Y|����N�^��k'
�>���f��?'!�]�93�X����L�N7��ͪ�wk�o�rt����t/GT��;1��o���H%&�x��ȉ������m�Ξ������x���u��F�6�t���W�%��k ]N9,1?�{E�ϔ�A0�����\6M��4/�h���[� ��-#�"�)����I84�аq��l�y�҂@̲;[M3�X-o��]2���.B���%���I��U�f��y�qH=�0��mR��"��2��
�4.T�ؑ�����:_�Qm���y�Į6J��9�'O�a�)sxA<�0���A�w�0<����s�5;���G�(Ѝ�c�o�}B�P�5��-$*mŌ94��x�ur`�R�k[4��<+mi@!����eD0�F�\ťvK`�y��^� �6˾�'s��1|�����򶣍ɼ��
CÂoUKMZℾ� �k���_�e�1�'��GQ���]e5��t�B:_x�����.yNfӵ^v:3y%$�����·/0��8P+���_�y/�C��+�mf�D�ҫUK��`D�@�SL��l����9j�,mԺ�UY���������]���/&�$�ei�y� �V�J�3PJ]���'��Z9{}�|�L�5������^��#��	��=,��^T�<�Oj�-*Q+�����h��D�H(XLVk#�=J�����<+�/��	�9l���I|��F~:�����@	q%b��KU���Ad1���F�A�w�nJ�?�J\����b�3��%�gwa[���7�sb ^�tu�݋!/v�Z���e�� ���F4r[zpO�U)Ǹ�h�d$���*���O7�.��w�w�Z�؄�E4��搃-���]�r�8���{��9�t�|op�rv>x�-�k�+w������I�aSظ����yy<0����9��<xOV>$�({����9ְq�)�tE���牑@]�Z���)���N�<���1 5�/~� �mr��[S\��s�FU�9#�ZZpe��5� ��?��!���2��d��*�*��Β��z�F�y/�$����D��!��?���)�*��2X@��������v���e��G�K�d9����%bIh	�E�~�a� :�0����
=}��,�7^	v��3�������xC��-�]��ʃ�-��`������Ǉ��I)�T[E,M�!�ǫ�2Ą=�ɰ4o@P��ݾ�
(׸�!���4����cM쏻�u�;�P�(���y=�Q���.Al���ی �`��?�b�L� �jq�������������R��j.=�"P*Q<.�#�Q�gQ�W�Y�JO�C�Ë_)��yi���,55\���4�|��yފ.�6�X����	��9��B�BG *����R�rqU�Fr���t͘�%G�W��H���ʯ�E^�]sd�m��f��ա'�doU!oik�}2U*~���2���	������,K&X�\�(��@u��>	>8�Z�\NI��e_�t�hr.�G膛�Fp�9��B��h�ƋΤT;����L��c���[��'�,�8x4
5͸ �� ��?5�X�����{�Br�Tv����7.�\��ԍ~��U�qc��p������08!�w9��}6�F"��^���6(�l'�P�5��e�x�K
_�?gM�ՠ�ݼA�e7��؃�=A(�)D�qkLm��wtC�Z�8��(��CUE0:�v�g���{I ��HjK/f1Ⱥ�A��8�')���0H��:�[��<MNh���.,=2	��b-�0>���9���١�}<��c*ޑ.E�=,+>�␕�.-:�^m���Y|IYկ|�E�Vxy�6;ye�z�}a��a ��"�7�e��	�A�L�z������槶�}z�0��)���~�CM&�˄������Rf�Fs�-�jV�����_QGmb��<Q�'���o�]�W�ȃ�X������\fH�>��F�&����4笹���q;�	d�߰�AO�Fl,;R���%��J�d�OC�l;��	�Q�7�c�������Pbt9��>���`^�Ą�zA�Q�4x�ո�`uWģ:����R����̣�m�1�Jtd�b?z�-�@�ĭL�+��Q3Qq@'�}��kB����9򸧇�7<vk��~/.��F�V	?o��%��k�2�,Ã���&���N� ?����<�]�5��䆘_@e B��sf<������m���f�5��wl�I�]J�t�`Ͻ��r�r!�o^�q��~�G�g��N���ᥟ�oD��-�$`�ԈSSel� z+ 
#��PS"���Ӯ\���5��w����@A=~�g�pխs{'�����LEgY���p���2X~��3�9�F�1����5�Yr3ԧ��?�_�GB�>W�|���>��N���δ�с����ؓ�O�:w�q�7�C�`�����+���.�$ٺ��/�`���yI�Z��O���6�$���
���zT���31~q�����m~��ϊr�gK�َDS����0�0\�vޡ���s%xOJrq�?yji*̲�G��p,����hIQV }HƑ�p���w7M��"�G�a�W�y�0{OcPw��?�b������6����Y_��O�<�;�cW���p�k�ڜo��P���\@����:��S�a����P%��������j��ʞ�;�8ɑh$����,Krݙ�JL�j�	�+M.c�f0ۥ�4��WÒ��DR2�'�k�����A�..K|\��s	�)K�8˷�5�a�m��*�=�T�P��mZ��.٠鉺~	V��2V�a�#��I �\LŶwi��5~�^T�� �9�B�g��ݤQ�����^�VV Fٳ�(�Í���o���TJQ��F5�P�vr�/�T��Gb�G�����6�GM���H&eJ l�.*��|+EDKc��/Yy%s��rV�hs�bᦟ-~mໜ@�N���o�93rk�4kD+�G��hI���H�<1�t|+�����Fn�=`Є�6�f3����=��4q1��1ن��s�(��
���=kU�|ȗ�û7y�$?���ʃ����m����k��m����|^�	���l�����Y+��C�.w�P(�7�:L��8��X�U��dWv�)�N\�.0�N�a|¦���i�;i��]�,O�� �����������j�S��g�>��>q��p�^OF��iq���[@$���F^E���S#�Ww�kV�`���V��p�$P�膶{�7�(���Թ�˰> Wc�ʱ�����h�>!�=���Y�D��K1�_[�������ES�����$��p.F���^i~�yxR��1k�SRx;Y�����ݣ���ק�\������	��a���4����Ï�P� 8�n�<�-�:{%AJ�y���h�� Sz��S�lVG�A�g��(.O����F��C]dq�G�����i�A�l8�-���!4���zגm쬄W�m�‵�ep������z��3F��f�\�ƨ���w��9!M�ӑp���"x�j�K�Ȋ]L,�/��H��l��ڼ�/��������F%�g�YWU\�[���-o@#l\�S��JN?kq�׼��HW�'S��%H4ی����jkZ�WM��G��lq;#wI�17@h�8��=�
�z���fpЮ��C���+W�}�5H�X�5��F�D����V�u��>��U�5��j�g����+:���wg����nw���1J,�4�I2Y2֭K���U�C|N�����ܸ�3�tZ0g�T+m����c@k�X��ӃT\��	��rhttT�3D�Es�?/e�HG�AATU�:7<I�r��k(��8̍�PK��ЅZ���F���Q�@|�Qk:C]�&��o�}�r��S���H�S���!�O=Q\\턨�{5 �j�V�Ն`a�D�l�z"����GJCS��sPf�ly�ۨM�8�qHV�^v�H�'|X��3�QwZJ��G�"��@���J(s�#i�m��V�q�b����4�9�R�f��}�#�^d�U���Ӏ�&����,�a/�s����&M�o���r8��8�;�!����_;�æ�-��1�3��yl.KX�z>A��uA�Fr�E	'
��d��O�>�2L��j�ij��/��������-��~M���W{����:(�*�[kw�
*/m��:��nŶ�y��	�gI ��3��K��|�1�/��Mh�)���5���:�ä��?Λ`q�o��\�U���[ ���rF��^Ls�{�Z�i�����W�fx��@fD�v��AypFW���7���	0]V6�kib��h��%�|%k59�=���PR���B,���^A�<Fy�����֬�w��߲����3?=CA��Q�%C`��%�(�j�D(�����1hT��1��ਂX�vی&�|�W(��K����w�F�.�X~����ǄF���En��pn�b����mҙ�2�qȸ�a%(��ac��܌j�.c��"���!g:�k����o���M�.�E�隧�E��Ϝ�����e��B5<˷M0�v�C�i���D�R��+(�^孒�R7�I�$�~t;m=6؁+S@�cB}!��X��dQb`����dV���b�����RQӲ�����X�b�J��c:Ze��Oh���?Ay6�=�COW��T�v���6����e�d��@��:_�'��ۅ^�Ьb!@�����2��;��ݚ�.��-��Kh+�Ax���f�;��a��C�G���8g���$���$'w� БC���dݸ���b��K(�bz3j`��E"� 龷:c���D	[���� J�-��z�Dn�/(��r�?�`&��d���Z�!�j�Ǌ��r�f�3���K�7���׃����r(�%.3̠�v���~�D	�J�z���U��Kz�O/�r�Z%F�=��D/���=� �2��kĂ�~C܇w�������.���)@�qN$Y .6���ZsT�+���bE�Ѥ���_�l.G
N�������u/�.HUD��}^1ʏ3�q����L�,(����p:���=]����u�����+��D�7���İ���ٶ�F=3xtׯ�(��r��y��v@>&ފ
W<F��ٰ>u�%�{�H���qR�}\9��<o`Ϸ�J���ڏ*�J���+�e֙%�L�;5Z't���w���$��n�	�mRy���G����0o�U�qT����é�^���K�< ��hѱ�ߛh/-R��<8��xxL��P9qD0�)��P[���&*ZͩU+��k�76eޔs�#�'�����nM޳Agd�V�xr:�H]�7V*���%җ�F���OE��9�Apʕ�f�hO�����g��8/˛mR��3V�Q�6E���E���ZU|����j��-�>y�(~M�ǀ��L"�O������?�g������3X�$;%���RG�G��΋���K�@J�������Y�a4�˜
nh�};I���K�l���Q�����e�kK9$�?6!5��׋ꖒ�!a�}��j��#��ϋ���"���l�jȹ��W�8�8�
�-�a)@28u�sOީL?�
E�����o�Ew�u	rHn�b	��P�QXI�&w�[8��ly���f��@+Zi4\�j�Y~c-S�p�mH���TL%�;*J�Xp^�N�^�
SVXZ♔@�F}�K'���uu��#������5��=�)ԃb�t�x���Rry�)��_���H�80
�������yY�x����
)��Q�v����OV_�N~|E�|N�C؃�V
��O�]e�-�9Y�k�(cuj�#c8`����;^܄�_(�j�la�7K2��!<�ޥ��BD^�/����('����w���x_��+(���	��uTf��L�����m��Cؠ8,
��k}ys "�r �W(}'@�ȒѤ���l�k��1�cXg��)4{Fa_Zo��j�-ű�>�*����O�%i��R��u��}�?2ªm	D���Fd�¨��� C�˙�G���t�I�r��/�A.��В�9;��]�����,uS�7l~gF�9��S�<]=E���:�8��}�W�(W���R-Q�!�w˼J�⬘�r�a��0���P/���w������e�;������g�ۑ��h/�n������jx^F(E���/^����\E Z�*���u�X�$�3�ow���|;QӍ�2�C'G�(&�96��s2Of��O�yC����۪�+R`�?P�l�GEh
� ��%���!KdO�Ꙥk�U�ꕊ���|6n$�ͩ�Z��F��W�HQ9]6���,t�^��(�)�ui۴q�ǬCa��P����<}�;�5�&���������$2�*��!�%�h�?�P���=�7dQ�����߾���4�̆*N���,����65&�g':�G:Kh��:y��� i�R������j4���zp�
'K�&��X��Q��ǲҬ��q��.�3�{����U>J�o�"�cЁ�ث:9�'����F���+��s���,�6I|HF�.<|"�bi�t�.3�J��P�����0(�#|�LK6���1k������v�c�W�� Nr���(���Z�,? {XR�2��A���w{g�`�!Ė�3A���5�%�H!���(�@�h�ۥ��m���bF�=n�`������X��5�$�~Rn\���;A���%X�jT�j(��?�@ף��(Э�e{B,�:"q�,&,D��Ew��yK�f�[�4`:���`�oĪz�#�*S�TFݚA�-�O��n�KSz1��P�VKU��L�-�֐mD=n����n��!e�q��kcK�ޗ���+�s28�xiڪ��)�($G��r��׍2�C���a[���p���3h)r�M��e���S���7�g������C�j%��P�ͽ78���>�-�I[�0�؎=�/���<9 WAc[��m�J�.:�9�E�����L2~r
���!��	N����*���>wV��4<��L�7��n溫H����.2�]�Xy��L;��S����Z(¼uӫq&?[�ֿ[���T��߶�J����Q)�.	��h�l��]��BY<K�bR͵':��5�K�2ELx��C��ؽ��S�ThaP�S��~�ʵ�g�1�r�W�`b�Mr�2,��1-i��F��g����1#�4��8c;����Ӯ ������^�������g}����UG�����?Y�Dr���N�����Iq���Ė��*
~
G��1}�-�4�9���
����l�	���AK�U�#�E٪��6��Ō�2;И�Yܬ���pcs�s�>2�nZme��������q�va-X���G�zS�"��D��.*���|�J�0��c�.���C?{N�ƃ ��<;k*��^�fMcL���b��!�Z���W[��wǽu_��Ęv����j+�P�n����:�	mL�
<�@���X[�x�Z�23 8�q\���89�{��?���"��TWhV'���*h��X\��=.��7������?��G�\z6��y$^������T���A�b�Fn�o����@r2�Sl�Z��}M����X�����m��d�g���@P�ǂ;g0	��fN9'�h#`A>�F����9���$��B�a !�G��H�ɬ��b�9_"䮱��L0����@%=�7�F�wFR3���[UvDNQ0K$3��6�dNNSi���g���+��<�v� >�r�3�'08Ђmn�z��+g��L�iъ��-3���ai�Kp0;V~b1����j�Nm�\����t�{��\�����y� 7T0�$�碽ǥW_e��KA�W6��=���-"�"�G۞��뎝�xs鴫���7���'%����ۓ�@x'�ȟ3���1���;�����O��r/��15W(�P���j�'��u��+j[}i�yl�{ʫ�al<�g�� L*[1mE���g��S��"һ|��ś���p2L�V�??�}����C��Lh�)��)��AJ�)Z�g{W΂�@�<�a3�vU�|<�����N���/L�����h��}���=KI����t<�v�*Qm��"|�O�9z�C}OF!~�I*��[�Ǆ�%S)����Iȝ�	�{sw���i�L���X�DJ}�x�+q����~�z�_o�bA,�u%����:��z�7ʿŮu�������J݌X����֬<.����-;�1 *�C���X��c�W
��פI�R1^�b�Z`�V�]mP^r�ñ �[T�������۲�,txR�r�t2T�.֑��j��Y��?��JsDKcdx{j��T�i2�18�~I9��	dX�/�3��[���\H%����ɕ'��Z���Y��3�j��#@�qCPs�f$���<s���0X��M���!>BS��ѣ�X�Ǯ��^��X�8#P����Ũg
�;�]���s�<7>���YG�6zƘ��ol(�b���.�*�.�:}���YD��ݻ@��C�H�3�Z��x��t�b��0V.�t~�Fs��/�"s�I���ַ�/}.�֔z��װ���ά�_'�;��#J�4<{o�n����4`�#x���F6�*\
��� '���w&����©)RΉ>�'<�V��k�R~��d�
=�D@���a����+���3�d�@T��,z,.�_��r[vޕC�!O<I�rY�y bk���r�Q+�/�MU�0`��w���M�^��l���d�0��F.C�9=�A\{��$m���LL�m���
%H>�P���h�����2��f7��v���ox����V�z�|T�y�yr��wNH�q�;�͓l(��0$c�c/W.�P�
mH�e<��2��
m�:�v柴������E���˶@"ƣ'H��|4��ͅ�&��C�u�䒷8̙��i���8.�a#�ziD�`����N(}�s���͏U��j�����Q��L\��t����yt�TO�|�6��M��}��ˍ���y}�L��r"�lkr������x$�Ӂ�B&��1u�H�'���ra�%|�~��]�^��Hi햝���ٵNĳ)��c>Eu����is��a-�:ᰰ5F<��)�aJރK膔��F���PIϺ4E���7P�duj�50�S��L�����"���KU>�i/O|�S;0�+%��ZA3��Q���:��9�Ev�P��CiB��|�4�%�|hl�	�=N~Bx��l.?���'�tI\����M�1%��ߑ<F�sݳ�?���ܨb3[J��W�{t�N���E�K�d�{@疃]�EΑ��ܴD��h��÷o{R~\� �k]}�C�˻k �e��mZb�q�Jwf��}����]��p�c�C�bg��Mod�E���Ld�ᱳP�d#��v�$��(t�P:W��xZ4Up^�Ҽ���;����	�E�X��km��6�N�KI]68ր1٥�w�nՀ��H�>�e2]�� ��<��x-bEVn�������I��Y���l����64_Qל1[3I��b��6jJN�U0g1/]�u�I;g�I/�&�$1��p}�ZQ!cs�I���R�]V��z3]5�Z�FI0C��.c�C]eM'���O~�(೓*w�?���v�\�dN�p�Z�w��6��M��l��ܗ���Ԕ�L�6�k�m��)���Σ�� �,��J�SEi{�:tb4*�3�Ի4�~Z�����~:��˕uy�f��K�:�����>(�bM�2pFͭ�
]��ȧ�Ky�As1���_#��ȓ�n�2��w�]0����E �b�j�k�p�i8�� S�<�҄L=$1܏d�}m2�GUDZ������&��D�^e��-�['���ܨZ�����(�E���9�:\�D�.�FJ��J�7�Š!�~���OܥA�L9������D� So���ǵ�d�r��O������nئ��>�66�Et���*6Pdt�K�I6��qA�o��1�e��w���k�k��	����'G>\�?x�x[�|$J
K��:n A�Z�|�])܄Äʼ.�M)�.ц3k�_"ߟ�; �O��{z����[qZ_�F�r��������.H�,��/����>Ɛ*���Qg	��x�ވ�P�%�o7Ӏ�w=ghfF�l�Bp��j=H�c3-�	Qp˽��7�
�����Pa�@�^C��s9���t�/zar�5��+
��TcZ�R��.�1���m���!`<�"(P{�' 6�wI�)�2ؐ2�G�A`���Ɵ>���x*\�|�)mY<�=3z���f0��N�DtoI���r����Dv�DyW�FDWtH$�x6"���L{Jl���N�o~h-��`��`�0��&�!u4l� ?'(��"���H�7����&Yod	�: '��<���HB�3~re������'Mu���6�C�~]9��!���Mz��U�4�f!g[�Y(	�����y��ͱ�#Q�\eE������3�8`�s���E{��
^ȵØl�	SC�i?��\�R6���I��g+������λ�g��vh�V���ߥ˟U6��M�f4�X���AS&�l�!t��X*i������j�&��2���f���^���>󠯄Mkc��L�V�[��x#>��ȡ	��ĳT�b����-Ѱ�X�,�ΞO�G�<1��q�wHIba�얍��/TGX��� �7.�	�1�cSv`l.�(�'���DuǽP�d�;]�(x$?�ݸ��1%!�����8��se8 �r���ԘۥӴt�F��W^L�-�`6�O{��s_IN:�����"V�\j���TED��*�A� ҶV�g ����^�w{���Fx�G�0'�.���c��iZP�����U��I�-������J�&6{�1f�s[J��������U���Q�Q�o����#��a����K\��;ua��]����mL���6`?VS�ؑ��->|Ě�"�qp��A�2�#�n`q=m/^Fg���g!��\:x���8�e�n�y��Ơ�4�_��HӺ��� �@}�G����Q�#����I._Ln��{'
�����-��nH���+����_�J��L#�Ծ��A��]�'Q�/J�Ĥ�n�E�� ���	��J���d�����U&�o_���[�]Y�h�b�W�2���S+�����-�S�J�(���2�&�����C킺_�X,���{k��,�ɹτ�fb[�,�1���bB,�ǳ���0%!�z>��O����08���i4%z*���8v�vK7�|�0{�ӆ�{�I�T��띾��Dd,��˅EC@����tC�TTGe�^)�ҽ��ݒW�et�a��u=�W�W���1M�����%����Ġ��x���}S+[��ε�Me�L�I2��0�-�HH��K@`V�K$�ӷ���?��)���
����|=;4�} \���=(�#|m17Y���5u��`!!�e��	vs���~~�eK�1d���D�]%b�|3�,��Y�)Cp�N�0���zJӸ_��/�7�2�)sB����W�w�)hJ�PY̧l�ER�'6L/�˹�_����׋i.��h}���w��v&Τ�C)r�G��A�~G!ϱa:�Y,S��-[;��R܇����)��,Yl�@�f~6詐�r��'W�'�4�/�'�-�����7��A�>~f^̅�ݩ��BG~���-Z�ގ�χj��n�`�H���ѝ�1�a�&�N��C��]m�p#k%-,�ߤ`u�)k
����Y��a�=����Z>�&�e��A�f�"�C���o�T�po@%]HߏIe�d��>��ґJ�`c'DZ����J�s�j�����W'�Ba=Ϳ7X�|
3n��n��KB��	5�"��7�YLh���7b�f.:3y�O5�fS�4�$`9��4��i\��=x�6�$��Q�!|Ű*yļ����"�Γ�9H�������j�gB�N�at�8]/`�����y�-��.��DB%T� V�7͖����8�a�%���� �f[y�>�%q��A�1"5B���gAf���p�S�W�D��������G�+~�w�� ;a..RxU��>2�q�s��5˩�駤�v���1%ę3����)���&Y��b	F�pA��W��+P^�A�k&8Q!LY�C�Z�~:h��r3	���w�})7���f��چ�O?3�{7�,�~ʱGJ�G|tn�)�ׄcJC�wƄ�	�Ƴ4r�撐M:%TQ�({�P����/TM������^["��\�wA��}�}!�(�95\��8XO��f�o��q����͍�F�=)H�PcN,U�mfizP*���f*�TY(�+l{�5�g����Ʈ�"��|30�L�1Q �J^Ew���8�{S�=&�*!�s`?�|�9r�g6$�2��]l�S�z�]t_�MYB"�jZ���:v�Ãb�ﭢ�Zm8YQ���I
�|�l���~L�J�'��ߧ&��[\�����&�?°|.��W%��Ȟ� QG<�A�#�!�f/���4�T��,[����/䧝��s� ��|��.SUq��ef�Dd2�'s�m�@c2V�ب�{�d[�3J5M)ay���a0���(�?�G��]�U�}03�"���HjNe�����ۨ�@���1D�'�a�T�͞��ke7�֍v� 󂳮���^1t>(�À��@����-w|j+�e�4'5d�?
���~�6D�6���gp�g�%X;C��/�R�8o*��� 4�f�8�׮f����Syd_�Yx��a���+���X'�oW`�Hm܍�Z�#Dk`�f1�emM��������z�nI��������MH�C�rkL$���/zw�)7BŒx��B�=� ��:�-������vI�Y�.�'�s����+�\�>��h�#O���S���S��71�YtO�a�J��s�&�3�}������Z'M/}&��	�?�rpPs��,N}{�R�ߕ��1����:+�h�@� ��)�{Hߚ}Us� @�-þ��{ts /�4�2[Y=Ժ�	ed�	� �}��:�d~�߄A�a�*?<C����6�ؽA�2�@X�#@�(�g:�#\�@��l�-�XK��g ���B��r�c�˓?eԾ �G�������fI����[��	�� ���0�.5ڬ9-̗qb�w@��1#�G�����H��b��-k�D�Gk c�[Uw�T����ZU;|�V4��ۺ�us�0h�}ū��.m���I�* �(GE���]�lW�����;���	���*�ue�5"�}�����5�+mi�/J�%�A�r��{dH+$�]YY��ԔR���)+R>��8@Ϸ����ƺNQ�v��F��g&�=ޤ�i�t��y,G=1��� �Q7�tĆ����(�2�߸a�|�
D�a,&Z��]"�0j53J�V.�''�n�U�.Q^�߃ z���{.�w���t���q;�VhV�=A ��I*7�?<$�?��")�"=���|X2K�����EW��a�{pgs뱮Hc�]�X皷�U�>a3�3�S)@6�J�_�Gf�9�r]�kɅٱq�ֹ��H�itt���8`;�!�uz�m�W��t�td\��2#�zaFg���ї�n�kQ��Z:@J �������#_ �kXJ�����p찫�C�ϕ4��P�
�}�dQ��mJfO�+ rɱo���|�t��H���WF �s��i��o����s޽���p�Ă3}e�������k���3�">�6���ԥ���Xo��<?����-m�[���u�O�x�N7�!�|�KR��;�ӔMz
���[�!�Ղ�}��P