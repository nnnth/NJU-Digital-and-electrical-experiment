��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��t�x�}�Eg6�3)��I_T���@���B��A�u~1�c�(lW�7ó�I��o(���ت�n�2���ñ���o�!N�Z"���ƛjz��IƟC%?�X��IN]�C9�cYf�o�K�{���V5�h��߽fY_��~HvB|��R���XLl�U�U�Ɠ�iN�[6��&wY�ZΡ�{�!<Ȓ�����}���R~h�c�|.��
�o����u�|��
�pL5�6Nb2�
԰V�l�t�p��^_�Y�Pϲy=�A������P}H�6
��"`�k�������,�Yb7 ٦��jm���Q�DC{�ʍ��m{��='E�@]����'(L}�b�4`;�V�79t@(���3m�N������ܝK%�w0L�a#�O�=��n{���5&ƾL�U���u�f��w�4F�/u$<�劒��V�ۚl���.����Yli<���Q�d�C��[�DE'�2Ob܉[-��9<b��8��\�1
n�&� �P�7�	���ym{�AcU8_J6�:��"9�Ĳ��q[�3�~ߔ�,d�CJm'�P�����1�����?� 6CA�3��HL�şe��b��jƄ��'�4Y=SO���e��{�>�i�q:=���G&B��Q�L��gLߗ��SF��������Z��S����cM)\k�:z~=����&����������8�a����:�E�|�\.�L4`���ݹ�^U:�Ϫ���<��oʿ��N�j_�f'�y��/k�jk
�;��_����������B��n{�Uo5 ��֬W*�FPc�/*�
�_T���!�|��^��D��z�n��d�V9�	G=B��0�B����޻2�Jpt��%_�|�x�i��PƄ��������	}�f�A6,��ⱝ���B�e!�%�j��Ge�]���#y�@�MKP/��c�F�N��?�+~m��&>2�?&|�	�Ϛ�_�V���;�Q��5m�Z���X}����Qrk��9�d|�.!ç`������m,����A�O�Kd���w�*ⷅdH(�~����9��$�MW�w����3�� �O^��V�ń�4r����e����!�_=� 7�#�[��K�h��C��| ���K�=�u�5�o�4�q�u?BU��@�)�(a������Ю?��b^�)�fe��;|�j8	�Ҩ�٨�������v�&B,���p�95���c�3�]Ȟ�:�[G�Y���p�_O����qH,u�V��vhn?���Y��~�ww5�v�=[�A�.��~��o�d�dWmv�\����!^�š�h�I( E�d~M�Q���!Lp����砘�����{���y�Y�[�/����^�T\�|��rIōa(ܑ�S��@0��P�%u���+K.EY��:Tc��8��a%6��3g���?nq������!25����-�b5G)Oh\�ϸ��|�U�*�u�D�|���(?���t�Z�:�d��R��1��������x9d��E	�m�(��AFJ��Nl�Y��M�N��Ş��x(�r��3S�)��o�ǆ��_u*0�r��S�b�[w!��z�����)7娙I�Sێ�,����� ��!i�F�͆!�A����V���4�g�c�-E�}���˙�fv��	}�-�ݙ5�U��P���Pg\K٢/�і��_�$J�%����8��6-Ѥ���.�	Xyt���K�����.?L��qB��W�r��T��_UG;7'
�X0����K�2Y?���KC�nTO��Ձ���Z�t͹�Qɏ�VɊ�j�F/�/�Y0��}M%'��	�Pf�*��~����&؏D�\`�����y�|ߘM�}#��-�+*���$R��t��Ƈ�n[�ؑ�$ٌx�C����0��E��އǽ�7�{�B_6� J&�5��VSs^Ϋ0�7s����G
o'�u���@j(������@��M<GS�u1m`ʕn/@v��i@8+cu��h\=�Q�[Wz:p�����׻fVj�d0�KC�DL�������$s�^�`U7�s?{�R���)�',���@� ڹL�1��&s�'$���V������H����꞉��{�_s[:�6��|����`yAR��UW���mk>�]]@ɖ���$n9fyf�r��ria���)�v!�V+*, %�{-�=��C׊���^jK��E��4K^�n�>��@?�����������m�q�~���#��P��f�!�?h��Z)�]�Zk�'�h\}$��)�̃+���8DP.o	j���*�bI*Ó��]Iυ����-��<�W������y�[�^-��1o�y>T}(A�E�h�/�J�dd�^#��G,���� S�(�"7R=���!�J��0婼�c �k�����FAf{Tu�v6�0���| D~�M&��V�Y�xzT�Ä�r:n^2���������%#�e����^!ڛ�r��˞QRQvX���5?��_-��R<�	�b_�NO�>�H殂2O�Ш��^%�1<�P�T����N�AG�|[]ZE�]ѶbR�<Di�O�$�;D�T�9˘����s���ls~3���Z/ͱj�eN��v���P;%�8Zd1˙s-R�\���C���*�au�ع� ��A�7L�KL�ǎo5�Ji�)v] b�8�翇n��>L�J܆&cOމ�W*;�iO����X��Խԭ���4�2��Qi���m�F*�
0�%�?y�ٍg�ûH�غb����z�hI(?-��E)�:}��"��7�Pe=��zc*L�]6�oZ��4�\������N��ˬ,�Me� ��F����D� �o�6�xs�	�Y��x�;��~�|^UQ$�A�ɋ�L܅�,��˪1�h�<�6����S{��O��F��]�n��[(-���ݵ�����C�^o��hG��8uLނx2�w�z�[0A�G������kN[���Y̈h{s7WZ���>Νe�����]��z�Ԥ�&�8��fI�$�`���:���W99;�k}��v�Kl[K!#���ѳf���L�Rt�����3/�W��
R�����+ ������#���[�l�vm�}.�{3B��'?Ґ�ˇKC"�Zɍ����Y�>gN5�
0��&������`Y���r��ߩ��WZ�.��B�xP*H	��"v}6��P,/1��8w�$#aWB�|@ � �[X�c����x��D��RS�yE����g�X��р�q@���jdk3k+���5YҜ&rג�MK��ޛ�2�u!��whw��}	=&�Z�\vY�jX�	p6f����%�]�/�L����lN�i�g YU���2p���>�c�n�.��-��&�I���x���F������zȪ7IS��wթ���#��NTN���B�P6�&9v��\�/��|UCH-�FF�_G��,⹶F�,kM؇$R���9�I��'��C��򷞍���\�0d����x~}�z�C�pE�|e���M���z5tA�����eo�%v���J�ۍ��y�K@���m:�����=-��> &��^nҸ�T�!BԴ�����!���� R# �=���<��0/v��5�g�c o����uT��h��R�Tx%���T0����Y�"�ӭ����� U����,a���,�ɔ��nA��E�)$p�ι�C��Ty��|F~�O�JX!�y	��n=�Q�7+
����_1�a�|������
�i9��3���e�f@�!-&d��|G����V���ݟ�is�P������p쓖�}o^!^k銒����^�uB@s�)�̙����OE�	4���u�h�d����m�e��,h���T��¼$mYLQ�p�ƶ�(�����S�$�?��a�pd �Z��w6��rS?cj�c!�@��L���|��z�m���Q嶈����a0�ms*�Р��ߡ�b�CVC����a����P�?R���x�7"`�xnap�2��^�=��ʗQL0B?�#��}W���h���6�a�^�Z��}S�ow�V �ܻ��G���8�2999�?{>t�}7��[�K�%o���G>��5Q��Ç�F�W�Xy�|.5搗(
0c�N*��ܺ��m�_�T�ʱ�ݎ������
�7k��{ͱ 57g��IsV����o�.3�?P���T�}I���wu����koI	�цW�n���զ@��
�Z�����D�'v*�g�����
�J����7�Qc�T������2�<�pw�]���q��H�Z��&��O��ٳ1��y�w�;��H��l�D�q�׉�oޚ�i�G�`o���U��PU��š�o����<�(�>ʱ�*�r�4��yP�A�� ���;�E���bܶ{���ud8�b}'���#��=2o�~��D.v�	N=Sԁ)�����$ "�p���Ui/Mϙ�=��R�~�+��&i�K����� [-��q�`&-���5m�0W='o��Ax�]����
.!�����l����Cve��7���(����IgO��Y+��T�9���k��'0w�7^EO��w?3l�w�Q@z������/Nʪ�T�2�Rܟ�V�D�OS�P�Ryuf|%��V���S�Q��5RElQH�_�AIZ�"���K�G b��Y�Gc-%vΟWc*0���N�?�R6�z�u�yԧS���������Nz�����.��a�-,J�*���ߢ�����-�P5c��xU�G��cg��։�[�
�b-�	�Qs&�6цU���?y��+�@�[tl�_
��1�����KX��rPjrRS7��d��4��实��Sw� ��op�UvYN��r���'�I-�k�a9��c3�Kv����g��6�z��J�]u>:!��)8e]�;��W6�'��x�E�}`<�B!�|��#��t�-
���7���i�DЪ�!��f}�k
�@��Ont�Gux;o�M�`�Ur�]FZ������ʮ~	2XD�P�'��O� -��U�`�2�Bɍ����V�Y+���`�����g���x�sV�]˗�l��(d{�(��[�K.��M�3[E*�裍}�z۸Ɋ%���(�d2||�<�������V.Y���v���['����,�%�Sd^�g��f�s�şDt�N�d��pC#��=@��@ �6G'�(t����C
���Ji�^��0ii�d�p/�b�B#�ۺ��-��yB+}��	ߧk_�d�"5˶�v��;�W��U�oȗWހI.�F����8J*�;�# C4&W�ak`�d}�YB�ߺ���Z�B�T`��\��I��.��h�9����ǹ~�k�)TԎ�w��#�Z�_��.�����u�7B���Q>���Q�˦�I�l�HE�E8rp���<g�ь��{�'�9�n�?�a�3A�P���z��Hbм2�JP8��	{٘䜥B�晞�{��Gn�$ދ�%['��{EMy+&�U�SN�'+�|9�u�2��![Ǜ���;R��f�+�@V����ZV�h7"2G���]6y���;r@� �V�$�0G��7F�N�T�G�9��ϗ�!��q�C�*}�����t��哸���@`E���	9a�j�xcbR��ƶGM��d�k��'�9���]���6�k���GU���i��C������������=^Ε�"�tr�n�ppϗ�O9��e�:㜆n�2�nJ{�:��QF�W�L�ѯǽ{%�5�7	(w޵ H������`X������������b�ڝJ�Z<�p�=���)v��5��u]Z��g�� �p��/mB� �ܪ/Bqƾsp2w-*%M�M�<�z�\i�_�mV�j��,ܛ�CI����х�H����A�Df��AO��S���7�]W���L���� Y�f=�h�(��k���5������	�;R�RΡف��n׃۠�R�S���)���岢��revw�CEH��;�ݬ�^骸�!7Ằ?��ݼ�J�����ZP���t[���!���}Xt>Q�z�cʻm�`a�t*	gY�D�_^!��S�R`�,�N~�9�އ�XLau����
��Y��K9���x�Ը��Ɔ�S��fNo�Y���4��s��r��]^Y͟�Ӯ�]��E�Orb�ߡF�,�%���� LX"�i�O�t7D����{#�k9nӢ4+�'���������e�.3a��j�̲�j0�b&6���x�CY�^7�e��`��QpE͏��_Z��mްR*����ja���k�3��?���G�����,���6� �{w�qSZ����&�n|�	��	E��ь&)&4�+@'�v�4B�7o��L1��ɪ�_v��o�y{�����jO�5L��`y��F�=�;=;A9Tm�oW֙h���ۂ���a ��(J]I;{�0��Q�,�ַ�����(�+ ���xc������S�P���d�7.�P:�Fѝھ��t�>Vr=X>C�1��g!�W���!����}�� T=Xs IrS��:df�b�G9ܽY���h���<���ݔ��]ki��+}�n�v#H�)Z#Z�� ��cv1TP�2ʺ�� %)�O�vv�����͛t�\�$���I*Up<�����0^��-&�4����d/r�q,RM��ONc���ؓBC1�">�/����ֿ�y<K~=�׋P�WQ9��c��Ԛ�a�	Vc$�xp���<�ޟ�a}O�d�	��ۉz�����&�D���Ԇˀ�B]�H
�;5X-Q�����r��et��V�d�.�+҉SjG&�c'o��̱��T��w�m+�&�:���v��i]�I~��=�]�_���� PNM�� +j�hG
;�k%q�t��� >b_4����BB0�����*�Թ��̼�d���7Jψ���2�G��ŤL��V�c�MKPJΉ�ׄ=C`�$Q1����^�Z.ߎNO�8*�[{]l2mɀ�&�����z7�I5�yxީ*Er��+��k@n�M��|Gj"2.�� QM$�T�;@Ӣ�:�C?�z�Չ̟���Iq��Uo�����k�Йe�"�~ D��*����E��BR}��(��\����ǝp�i��<�A��|=�-�ض������P�@�9�/[KJ u�PU��jc��oR������Akw�V����S{��ti4�Bߤ�6+V�	�~W�O�k��A�\6,F~_⨘�t���9Q�Y�Ĝ�z!&�~��`Nk��]ұ��`�.�]�oX�>5 ۆ�����R�����>�WɆR������d�� ~d��X�^EG�e��Q��r��Uݦ�	��\2?�Q��I�)���u+������t��z�9������9�H�;r�	�-�}����R�y"B������]�i\�_�^D$Yb�w$j�a��!�>iN�Y��#ϩ��$���zl�/�m�:p���pD�O7�� �S<g"�[�!�U��P�����h7%iӐ�P��:��S+�爤5'6]f�M.QiC��qA���g!,�pm=��c̮O-N�s�I�^o�N[0'��'Rfy��O ��ϧ��g'&p�����v�n��y���5Z{���'ic:�pT�#��Ge�<�2jqoÅGY=�)p��@Py\S)E��Ea3'����.'�[i��J���qHC���&C�Ք�B
��7����.��Z����U�3���Q��K(^.zh�q�r��������8<	b��$$����MCկ��	������ef����e�qNhU)�Mr �qʡ��Q�`�|��O�J�y�9Br$��g�<6N�<pˑ���;��9��3����;IH�9�N�:���)l�)�K�"s���
qO��-��Ij�]G�W�k�'��6;�P��VhY���o�";6��壛� )ʤ�lEl⤓�&�j\t� �h��`�Y�6U2>��mvi�2�"D��19Gx����N�Q�:J�p
	L�/�#��_hM��w[Y$�u<c{W9-J�=��5f�R����N��k����n3���U�x��6����p�����>���r^���X�����Q_�o���?���1&����-�L&�'8cP���/���;*B8�����厏�G�7Â5gMtY�_ �)aߵ�1�B�~��4���+6U^&5�:>��mι+b#�8�Ź���T^t���7y�f@tu�t3f(�eu��OU<ޝ�j#l	������쟏�^G�ё��7�T�n$�dS1��2���MdUs����\��he�N��"ߠwx7��c:�����[�zٜ�R���� ��H+��W �]��k���c��Bv5b���	]#,H��7s.�	r�B�1\P�3�~q,ֺg����J>�	�&N��
*{1�䳲0�w�������d���W��D����>�仌��T�|?���`sѱ�4/<,i����<3nN5��w����'#$�c�
l|ϙ{:���i�M4�Cnuhŋ����#���@�E���9�_F��5#�d� ���b��Cb��W2� �'����ǲ��^2T���dD�+��T�&c3H�JZ$�|iV`���R\oJ�N� �K]B�P��@z�v$���aJx%�DKU����N����˵���k���\�顺'|��l���j�QJ�-T�ׅ�1��V�V����՜F�`�Ӽ�i��Z�<^��2��]h��W֟O����8��I���&�ڇ�w`��VȏCm�S1�C�/�m3�_1;���}�=�[�H^�.� ;����zPrn!����m��a׵[E�1+۹+�Y�_��&��hy|loFڰ��+h9�Z	�N?�s̙�XL��'���q���Kb$dX��t�+�ġ��=^�9h~R��b?0;aLBBY� ��2W��6��.%����k�׹�\5ڣ �1�7�U��f�#��ٟ�yo�l����X'�E��*M�pP!S<o�C���r�[�Zj��!Ug����@SJMt�rْu���s�X��Yw��䗮SYvu���<�V��@�w�"@�^2/ݻ[S#+j�\�W�"��ޑ����uI�ۤ��N[�,�)Q/��5��o4N�����bQ��0���.G:�V�wN���~�4`O5�����Pu�֗:�NH94}BSYOvh�� ���]"s!�h̫m{�p#O��MZ?�l������x�k�7���vR4���&��,�Bߍ�#�
n�ݜ���u;%z��i4w��Z����A��ѭuq&H:��h�/_@� !3 �)������˝�j�۷c�hv̟t}�f��ڌ�G�⠷)��)��/�1�\-a NiNs��.v��`�L!⦞+&#�B���-�l� 
����w��C���B:h����C`8�1�JY���AX�[��k�Nt����+uR���b'�׏5��{ēQ���9��K�?�ޣO�5%�GQ!FӘ��#�s�HT#�$�$ c�Ǧ�O�N?��ü��K@|���}B�9��M���n�P����W��[Y�l8�^�H�#���]7�L8R�<I�c�x���� �l�1�Q5��L����.J������ГѰ^�sI���v���+���ֳ�;^]I���A2E�\R�D���z��E�MA�Z1�0ѪY�7]*L�a:ýJ2r_�}�r�
�ݢh@�:ta����p��:�d-RCE(dx�<Ӵ":���J���J4����~�շ��vxx��|R��ӄ�T�~f$��LЏ�G���>��(&7��`̱mU ��!�ݒ󨫎R���e�!�Շ�g�x����P���ɠ�g��I��v���<�4���*��J׫�-\z~-#�T�S��G��꡴����1�c�G쮥4�C�������2&�ݵ�L��&�K#e�j��4ӹ��/*�MX��
�n�Q��є�{3�\���P�+�1�CJ��L�}�̇m32��)��X���¢�L�I,lͪ���77&X�w���Y�0h�t���Yn��{��w>
�*)i؂��;(\��+�Ē�}����ԅWR��0���d��_x�jpDF�������n�mR��9J�	<��aiXD���C�{[�����׍�'ny�#��
M�,2B��zp9��4���G!�qz��7�_��DYo�G��JF �!�{�����J!)�]exb�Oke�wQ���Zc �u,i�G<ب�AE>� ��;1ZL���'2�l�4ӻ�"��y���jF I����0����*���T{.��7���F�8G�5��!gb���<F BܮI�����Ѐ�Κ�gc��`�r�Z��Xˋ��T��]��^�"�b�4�c�a��z��5��0������߻���L�E1�3�p�5	���J��X\*��XU��6��4[�z��װ��i��= PM�'ҭߎά��oК����̖�1O0���6i46-Kf� (y�RxR�쩏����6~	��yeL������
�����;=�O�p��lӍ轅}=2������{(r.ihU���
��<�^���8�����:�v�G�)*�~}S�����Q�2Q�Y�1ӕ]?���_�KB��]N�x�*��D%��pu� ��@�,:(f�W�]�����XIG�A���ٯ�VG�g���a�U�H�)�2�y+�k�)�T�w�e�w��#I*��]����*k��F9��N6��{�.A�/$5"`�W;�h���~Z�l��<��t��Y �N���[ EjG1��.���;�i��S&٫�C��Am�x'I��)+�' ��[�܍�q�L������@���m�+!�X�+�8pe�Vț�H6����!�,p���B���1.A=F�hSL��b;�vq��%�2�x�|ۦzFe�Z%Z��?�I�$����x����k�1���sf��������k���e�]��P (c^�C�b�v"�h��]��(o�8��^��$��Tc��ٱIj��Y�􆢓�.���ϩ�5�a-.��9BW_"�,�ϚPn�lC�a�t�̭�
"��h 70c����^��b��w��
I���`�9��&͊B��(���:�e=I����ZC���#%����q۫ u"�:�:���"�$=�4����ޗQ��M����i��e���=-�Z�^�*k�&�i��Ǡ��4���@P�.���qۤ����2�Egֹ`���C�����8�#���}��]$��s3�8mg�ñr�Y���hw����QWz��a��|��@h�િ��v�I�A�d�����T
P�����M�����2�_�~�)��N�?H�V	ڜ���/u�p�˿@�˫��o����`�o� ([Y9�
Y.����Õc��YH�,��)���6gQPr���%��礈��WR�.�-O�1��,�C8i"~��g��%{�Ӟ����Qu"l`�e�������M<�Ҷ,]��?`�=!v�#X�{�����o����8� �ǽ~���F���?@�_e�l�(8�dj|�8������9���χ{���pQ�*gǂʳ��\��!�+K~Y~/2�R����-�+�*/�h��3�!��r�He�S���%X��4��ůp�fg\�k�/\9.t.@װ��ȭ�I"I���P�}a*ygTu =$�����Qi�l� �r��s1��V�5ڀEX���VgidU�9�.��8� ��k�����wnlG^�΢I��&��ǹs0a�	���$k����6	�T��P����q�b�}
�Ͱ �k8I7����&��%o`��#������GdK3V�'��nu#�Yؙ�J�%�Sa�sr���b(+Ll3
YU�t�h+T��e�Bj����~����QQ��X\ƥ?����� ��1��H�'��}G;Q�z�)�������a�u���)wJ�uĳ��=��
�f�'��)��G�LO9�U�'�ǲ��̽ #.^m����˥-�#Vm�
�o�U�����S��	iՏ�l^���D��9��iJj���p{.k�Kp�q(���L�9
�Lg�}����	����0<�O�H�^���o����l�᲌�j]�+KQ�Q66�C�.8�Lx�!��vx�/�H5,�7%�hO�ﾲ�%#��;�)��SL�S[M�^@!�M��^�̰&$]	��$�{�WxjaahO�gE�k��✀���
�\η����Tu��}���CN��Ld5G��q���$���G��r�Y�WcUd��l�9��4���������ʯp�,���"
cB�E]t���WI��BV^�9�Τ�!� ����ݞ>X !���&-
��Z��cT�9�%�{�Tlv|�z{�.�O�^�N�?���#�7�b�.����ΠL���e��o��k������0O����<��������5I�	~��h�� �u�ꫩC��n$�=���� Sܲ��m�j��W`!w�����bK&{J2��+�����Ƙ������?ǜ�_���*���AT�F���>���9�y�d��tZ�)��'��h��y�kͿ�bL!v2���3֙�߈�w�B�T��%�y�'|�M1`NW����:�����s����'$�W���w	�ewm�/�Υ��������f�/�܎N��g6(/��k1�׹�w����'^H+;Z�z�seިH�,��;�Q8G4J���nBx�(�wH��-Qu�_���q�vv4BE��|����C� ���}_�Bhխ��)���=���\��i S|�����C�5�Dwz�?x��H��0N�ԏ�uH3����R53�o���$�����P��(��:K���hn]�2)��A���ZPVV��{/z"��3qV얕W��X���=�i�yZ�O9�����d��P������������+�sN�4"C7K؝���0���rI�m�)/r.�C%�D�>M-/�(ؕ�u�`~鼽�p�o ��ӠbѨ3zS��*(~�:j�G���=�1��鯻�M��������T8��A�k+;ձ�0+���m[�}��	�O>\���Y 
&.�c����폞�(چ�X�t���6Qj܃���|���&D�l� ���<[7�X��5�-#�*�~P�S'Z��&�0�r�NܢsX���Tv��%��Ĥ�.a������)+�:���4uq����J�m�sS!C{2ӯ��Ş��!J+��^`��r()C=��;-�
qv*�zF����
J��i���}�H@s灠[;-z{|/���Sw�mp���@���P<�k8�B�A�7u�-|�M�N{K��W��|�;��0��|���"l���r�>�WE�,��C��ڶM���J0nE����;��� Vf ���;���%�Vy�錄�>fu�\��y��7(]�js��	�i�n���t)�@	�31�]'������<�L��ܙ����: ��'�c��{�
���t^;G����9��_b�7kG׏�7�:�><���(W���~k�?��:�O�haI�|O%6K[ƺ�`)�oL��Y�I�r*"�
�^�L~�O��|k�I�]��>\��tW\�Z&6�q�`�>1]��c0��
<���v�ó)D>U#Afw�=�����B�(�[�dh��x�D��6��Tr�D'�D�p6� ����FyU������C$R#������G�vj.�H���_19���L�~�A�-ؙ�	�r�����3�n�J=�B��2��+�4�������(�ב7k%�Ϝ�&�la6���+KX]������r��]���}�Q&P�Q���>�h
o@�h�rP�h���\@ۂ��vf�!<ۢ��Ӭ`�%+�ׁW2_&5�q�&��é��B�gd���� �<�@]y�^36B�����Ӻu��6r�w���F�UnԱ���6��g��'��-4!�۶7���;���+�[o(V����7����gQ�������:��=e�0�ߑ6�l��Jt媺 ��d:�#i/�^��M�r��%��A����Q*�6��ei��&����P���)����,x����W1�Tå��풇j~
^O"���T��x��4�^��8Qiy��/7�t�_Vk��H��C�٘�?�:��Y-o
�j��LLpM��s�꽌������m�S:k���
L��GOu�87���>W�"/��?4���&�Ћ�.P![M28�&?�$�+�#�
]�`�5l�H�^Ҳ{WH�?�ml*n|�C'6��\��٦
����T�H�� :��w���+�˞A���	!>5f�)�5���cc��ץJT���
�t��g���u�=��-L8.X�E��i!��P���Be��"�=�F���'�����b�������"����$�NK�����5�9(B+��|Q�rj3����꧒�d~Ј^�mAD�>�
�c�k��<t���O���1�9�4��Lh}�T�@���m��!��p��՘�����#/�O~H��i��KU�� ����թϼ��d���9�/w[2���Fެ���d�'��h���)�ެ��4+v�`�������0}3��0�N���U���5�l�
�e ;4�����'�5%{(zM�!��=�-����Due%�~<n�����9,�,[ʾG���!��M4����\��1I�|�B0E�&��Z+�F���ޱ���ܳ�b,Ύ�_d�>��ǰS��~"}�N�ak��*\�p>*5Ȧ�X���TnK-yZ����|BJCG��&�!P��_��׌E� ��1Ro���+�yf�Ε~���#�M��&���떦ϒ�g�H��G��=�D�e�_do�����4�]����>�2Ct쒚�A�M[#36q��K��"��r��S��h��ұ/�qu[X�]4~������FF�$ +�� ��m��ky�u�ZWj�3G����.#���1�"z�M�[T8f��7��"zU~Fɤ��Դ�R��¶C�C�^�HN4�^�d*g��FIaQ�	��)�P�s� �vz|T�O0	I��1ŝ|&��h�J������z��朣��|��摛n��x��tn����W�(�Lm��9���� Ȱ��[��V�uJ6���όر+S�;3�+�u2H����\#O�tnK��9)%���$ϑ(z�Q��U΃��'�������"�Y��P[��*�{"����B��uP�f�v��J ��eH�� ��Fw|�>\h���Ŵa��� ��Z|
�B1\�9���>�ۑ�_���%�>j�C	\p"y+7*�5��YZ�����
����!���#�AzR�2�w7)����P�e5a��4���y4��[l	/��Ë���X���vAg'��� �4��
uo�i���ף��l�@���u�}�x |�sycp��*+8mB��
�O�	�����;Fz��G�":�� ��}0�:����<(l�V��y�Ul�� ~�N��-�v��R�bj_]2�޿ (Ӻh��[�e&&1mB9�YN\�S����;L����i�Y�Ǝ_D�v�L{F�<QU��%g���e9wf�^W��Z�����]���GD����U��m5�_G��&]���+o=`���nЙe�R ��HwrK��<���A	��e+���F�����F�?Ng����������/�ǃ�(�;��f��m2|#��0f�j�sˁ����"��܌|T'�US����)��V�K0�_/5�)�N�f+;�L9�~�Ȭo��C
#�p�sB]3��g~֭�dԨR'�'�wK�9|S�LX':�PŮ���wXN��{%��J��%�"��;�8�c��<QM�!�7'�F��s��o��ݙ��`>Y�!<���Yr}/0�I:��]<&=��T���%�DC7�%���-a0c�h*b 8D[�Vp�]?�{��g�ޭ���\���9���a���Ew^��j��Ú;�|���h��;�=�R3>fq�pmdb�έ�b�\�V-�Wp��J�@��"�W��a�!L��n�"!���?�s� �S*ȄoQ�M�����g�L�8��kq@���֞�}>�.r�oH�Q��F����^O�g�OE���o=q�'�����Q���-C�z=~��];F��ϳ�$A�`�_8(�{/�9��1��;g�eƢ`%�?;�C:��I�}2zֿ%���3�]NV���.��j�rU��W�ne�F��#�!�G��2��)ἒ4QG�Q�9->�#5#��yˏE��p�zr�"�Vk�����3"1�1@��� ��]���Vq����E@&�"�)i�`
�W��z��Z�B��d(2w�ٛ@�:.��b���Q���;�Ϗ���G:=��|R��W�bn�ܮ~����/�]�f���)fd��ȵ��5�����Ec�R��m;p-$`��7T_4]��ĘvW�Ҽ����g�,�!��
��Q�%h�L�����~�$��@Rd��$��c�����T)w�,"�Y�4G�q�}'�\�a���If"k���F�Ɋ-q�s�c�7JI�6�����A�Pf�!�_ƿ:�|�c���D�Z�D��XC��uP���*�&EA�6~�.H�f�6��*I%h!��؎#T@_rIǬI�=bi0c��o����������{w��!)2U|�v`tr�5)Цu�2|ٟ�(d������AзUGc/!��{ ��PN�=��s�_�!r����4U���z.V��#3�6io�����؎���04�3�I�:��bM�&>G���/��n����}51���h��a'��k�=,��nڊM�I��� ���@��6�������[���|��$\���իbj�T^�`~�l���y���Wz����Q^ȽOjx���;�!tS1�dU��b�wz���g���ˬ���k��]~d)��I8�כ�������Q�7+K��� гk�|}Ŧ�E��=˨"0 qRI�*z��ZO�aP RG��o�F�6A8���֥Z�i@�O������#�"�?�QѮ��h�J��B��	��B�D����(�5���#u#X���(3]�C�-09����Y��*
�9h�*��L��s� ��G�US6T��Oh��N�Pֈ
9k�E��w7&��bw �9�h[#"�첬�ُHU��]��z��5MA��U������%(�V���V+8o���a��6��Fd�EsԤ�Q�`�>�?e�t��&aA}��c�h|$�����6�3��