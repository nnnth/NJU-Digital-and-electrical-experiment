��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t�CZ�-�b/��.�X_4u���%T��+]Ǚ=���a��0~/��4/č��#˺Pk�� w��s�9�,����	�DP͂�+V�4�T�hz�%��ɳƪ�~��~��ÞߴVj�3Va�u���5�g�,��$�>7;���['��c��$����`''"qb�X��"*KN���7=v]՜֓$;�������!���t�T�~k���h�,�n����P��i�y�T�� ���-xj�*�5�� 􋋹�\�/*�M쫷��7�WG2���q�e%^�saZZ|c�G��_�:An�O������� ���N��l�o�}f���;q~��������e�Y��PM�z9�oL���b�I��D�[u��3�؊z�{�"
ń��V�*�K]��jA)��+��|�t�,jIj��R�ӈ�=���ۋ����5�Nj��°,Y�v^T�����]��f2�gY��� ��L�n�y�[D֞L ЁfT��(]�a��_ܑu�4�vq/\�V���ۈ��>��!=>���y9z�n��B��tP�e��܎����M2��~Л43�)ڤ
���!����ٽ�
�Vt*W��ʻ2���X�R�EoH^Ɣ�����,�C�n�}A��?�%wϞ֙��(�USPY[Y��RhS�w��Q��918f�uZr�5��&�?�c��s9��ǔ N
��:q�����.�Ŗ(��-z+�8� �E�HI�D�����ZM�Q�4�<W2o�ۑ�q3�2hwӕ�8n����_b	����M�� �����}�l,�к�&��V ��;30b�}���<Ĉ]iCD�;��r_���=�7�Ƴ�~�"K�1��Az"7����ӳ �"SZf>B�=�RČ�Ę�]�h}S�^��^�`6��F���~����G_��Q���[t������U|��;1�&�_~VY>�f�<_�el���-7��ڊ�z��X�!$�*`��W���~��Y���l��ͤ��Y}-GX��Q�}#�gS�D�}墊	����d0b�A�Re���*4�/h�� }IHI�h�!0Ch���)"��̻JV�v���1�.�Ԋ&�-S/J���{�y��=���e���-�nZS���������d�>bj�)���@��J`��c���Q	 �1W<g�V8#�ZboYX�c|�M��iw���{e3ض��:���o� 8�ŵ��̒�p�a1��f�u�7�!�Q�2QދM����͐�9 }�݌>}�۪Q�VDkFg�>c�e#���e����K�ݛN�2;Zg�*�`��2#лzzφ�5K�?@�)}ʺ�/��qE�CU�\:�?�v�]��!p֫��������(N���ܱ�OY���ȃ3�:ZS$E�Z�mH���9�g��^���צ�_N>l簙�a�ȁ(��W/�*��?����0�X�<G�- �i	���L��M��%�k�'�׆W�,����4%�h�i���&%�K4|,�s(��0�R�6���U�mE���b�ۧ�"�C�ҍ��2���H"�gl��(���"C1xO�î��X�j�q���?'n}����2�۴ԊC���yV7�Eɯ+��^J��I1������5�Y(�V���5B��2ԫ��(��`6_$��4�O�����4D�7��Ih���I��Q�����]�X���3�C�!@��� �i]�T�८��	�D�u�S�t��<�C�ܸ�~ǤbX�Et"� L��Uֲ? #�^@��h&�FG�@���C�0�0��g������Z�.}��JO�tI�FD�����a䗾�*�,���F��=r:�waX*�08�!�� yD�BϤ֗o��,�<�h5F�-�G.����D�ȑ�rK����?o?�u�y4h���X�
���UKV�悮��+:D�����NY�B�۟�@o
r5�\�:4�P��4$a�=����,(Kh����� 4�(A��L��}��-=�;y2���V��{b��&=x���K��Z�_��!�kP�����7�cj�PH�����pI8!��4��ǭl����e��TM�ɾ_""��*�%r�c���\�E]�P�����2�-���F^>s\<q���������Z����G�-C��G��?��Z1S0�'({X���`���"v9��H����a�i��G���BE�=|�k[��I�������?��e��<L�PIz� _s����I
&
��$���la��\��M�u�{ɍ���ֻ�vg�"z�;?��^Z�<J�<v#�{.���i9'z@�,f��+v݆�m� +�B�=#\G��M/v�Fn�|pchAe�}�O�ł2��ÆFQ	=<��j�B.�Xf�P��f�3$fa�P/N��Qu�#6k�:��p��\5c7�kaF�-D���EE5ZdF��߰Q\��M�
���"��p��<���o�Z/>�jd2i���Z!YQ�W/!��t��M�%B�3a�o\�ZK��*�/S�\��*��,��+�]��?<�uG \� �� ����K�=�/�Z�� @I���2�Q 'é�v��PK�����P�dϯ
��	$�azf6_MԟN�蜾���@(���N`?Ǭ���֚��b>�,F*��jNوU��<r���֋z���-��f���?�|w���{��7��(Մ��D��b�n�W1g�|��4��aJ�֦�Q�'ɱ����X1.n�]	�����W� �m�\�_":ƪ.�ܾ4s]�j�߼�|x���!���I�y	R����xݫ���\��籜�/9j�|����*h�)���Rþ�nE),��ђ6��I�G��q"��R&H��e�<�!�C3X	8Ц�g�Uv�3����)������֞��BU�C��ZC��q�l�޻ALȽo?oN8(|��i���N642�6�{��J��K��W�������n;�54�^D
,$qvz���n�&�~2(��w�8�SPؠ��[��?���[�k#1m���|��nb�ֹPXW�+�'����=�#h�M@��c/����L���*�wv�"��%ܖn���}�̷7M�7�@8�	�<��4I���i��(��/Ss����7��u�ʄ�W4��Ի��.N<���V��Cd�y��5�2�
�½<m,���{㹌�!��ֆ��_+�N!�:�/M��'�Q���r+e�2#%�Pb�U�t�>�@+fqvj'���;^�^e8�o�⨗	!�ұ	�;�x���+�X'pP�aH����E��a���"zF���R?�@�Nο^��E#
Ա�,��D��O�bJ���+o��GKހ\�\�x�����4��>�Y��sUA��/˩'Viwq��=����Z��
i�~�����[ @RV��5e}|~�㇚X����� Z�O�mR �:���ɧ�D�����>�Q�D��p��]�:��D�b"�_�R��ڮg�~-̗�R�"D��{���uo�h�M�J�r	d_,,��רA�:y�]���@@��N̞uh�[X��ń&G�G��ށ��B������d��K��p ���=!*-8�"I�����dE���9C�"O�B!6؏���h�
v$6�Nn�5e�^ ���q�COm��G��7�VT�@&ZI�S���t�Sl�e����w���m���Х�S_ı�͖d��8Bp��:�!����^��	�&�y�1l
�19����LY�*�dQ�ÌtS��sv��%��;�j@���^,���-q��Tk7�!M���sr��FI��(��*�r^�;�d��Wޤ�1�@_���s	��:��0��CG��#j�����An����%ye�r_�j�6R&�.Yѓ��,9&B��u�KKP��F�u�ӟ`���;��(DU+����4�D�M�/Ϫ��<f�y�c
O�����qDH��DD�=W���a��5*��?�<��F'*��Y&�ep�8��z�X���AI��J�h��ƣ&��o�'Q�Q`8m��$�z�(`���!������`��\�#�Ё���/#�}���`�ԙ0�9T� 5��Ԟ��X_���]�[8S�s�'�k����qf~g�a�k�K���RD�+@i�'����Y��j��`�d�Ueo��Ǌ�Kż&7!�9�� �qǁI��=Ѽ�Af\�5�:�Kz>k�����?�lfl��*�a�Ɖ�{�vLa?k��<���@O��"�?�C|U�Lh���)UW5��7S�^�q��\"�6�����qq[s�i�'��1��?�k�~�>�o���]v�}���@e��#(M���?�@F݃|�JnUy�9�^�J�pI��1S9���B�S�Sԗ�wL}G��C���7o:.&��3m��D�t��H��ǻ�9�sו��8h����~�I��T�0�*�Cs����\���r�,(�=�dx��u�8��z#����>e����(c_7y,�t���Ww�Z�)�G�Ć�M�M�oMl�0{��r�z��LIGC���g��V���F��fn<v��W�6U�����;�0*٠u�J�Ml��B_��h��Zg���m�8���^uH�/��,P���w����@��&C�$m�~郥`�N�P4`�� ��ӯ��X�o���#f�k�Ʒ��G"�TJx�yf]���*F6�h"\���-�,���~����c1��3�����R���]�R����5P��p��qbsg��O�1�XB�H<k�W��C�'�� �Jjm9����ob(tu?�����!���QK��l��ֶ�>ү@�\!di�h�.#|��SpX~R�����6u݉E���Y�qOaV�-������Ee����$��b}�4�m�h6�Y�s�wkx��ϒ�v� ����S���%k�V�+cR^��v�m�VSJ�T�������i|�̿ɟ%�x:R����S��\�]�H0�_c�&G/�,޲ϕӃ�ѵk�M�L2<�k܋q���`���@c��~�f(c~�E/�F>uP���`r��[���`�Rp�BP�b虵���'��ə���r(�����X�rc��2p�]&r���)�)>0�e�(.g�lw*M��v�Z���,I�M;4N����W��C6��Ajv��D�p����ћ�O`
�m�M�]�2��U�p��4������e�=h���w��b@1F��#F����mM�du��Co�?�ۣr�p�d#B������8��nh��ҦD�[�{��L�&nw�/H'':�j�kE���_G�ʷ��}E}�kv��1ś ��￈�V���Lua�%P`eEQ�߶�0~x�ۣ�eF�AnW5���'s&`ܦ�89�Y�/.�r�4�lT|�������]G��
n�Q��><2�B�*X��` ��[ʟ�H��4qKV�
h��GK_��VS۽�]3��qj������G�`�Sޘ�����v�k���}����_�k���[X�,n)�>�K��aH�
�� �M�����h�>���/�h�Tr�l��聾x�燌�A�bd��G�{��VƷ�����4��fC��O��G�(�E��*��
��8���B�(�����C�3j�ޜ(�k7�C��(�%�=į�D�q�X*���D����"���S~O]}|��"~����e�=_����P����hX��%2$$Q��c�s�J�:���Y�߹�#��֏���-�{6��� �:C��f˞�Cj?αxJ�+֒~K�DO��9Q�u��WY�Olغu���(�1?�9F�ɇ��LOXH��y�����v�5����>���GzQ��/��|�w�gw��g���:�� rcm���Pf
<�~��J��R���z�/�s�G����p����Ȕ�;s�c���w�mÛ�B� _wît����q�yj����s�n�x���a�-fL�4P�������,� �P
K�P����w?�IR����/t[�x��
E.�غ��9���IT\0�rR�& �Nħp*�/T�W����Ĉ~u�u4���D�����V�'���"t`]!<v7���f_�3�L�kd��/���Z_;�����s��ڡG���Վ�_�A��VLɍ�6O��w��@�Bf������B�I��  =�����_b�3��|t���i�
2
��3��±.��D�x�كO�h_��֭�`�`1I���	)\{/�rp�Q۱�NqaS�w:#Wt�	чY������s��� �p��1�D:�?��}\Ff�AVû�M�M��;�j�{�^5^8��` >���TC���o3�5���x�6�3�>���P� �B����x�� �,S�R��Ւl��O�6��.r!��w �{�:��[�Z�i�UizT�i�v���Z*m7���	�}��?�F��6]�mrl]��/�ВÀ��x��~xFO�ĥ x��$���J<�j���(Ëm�8���,|A��͠H�C���I$S"X�)(���%�ŧ7�*�ٞ�*��V	�ե�k�j�O��""$�M��wr_s��v`v���n/c��$
�UC�?�+�E��'���kD@Җ#l|��t=e�`:�I"�`:}��1_��!��˙SL.R�� ���T>��п����֗:��kQ`�)Ndt[�y�@��zT�8f�N�{�ď��&	x)4��x(�Κ����n�	���˯U�7��j��h~��������� �!!���i)������m�Wu3���$+$
�U~$z?,���EUz��Y+{��Ĕ'�^S���1Eނ��:�t�E>�W���D����̫��fsH�ru��<�B?�~&���&��K��2.�8��H�:Ѝ������'٨ �o�K��O1;g���1���8����X�x�s%�]���Uw�u"����똺@N���_��QS�u�3��~��+�����U �Hd�o��>` ���_��.>*O](��{��Jg�2�:~/�\��bt��<i��	�	󳙁bd��_O��|}�OaE3#+ߌ��K,��!v4�N�2��
U	D��ej�d������;����u���y���~��a�)H�NWE�7#J�0�2�"�ciR
a&Q��++>Uq�,E5O��t���(�a�o6ʭ��d�[`:F%>���9[�h���P��!`(���j��/'��q��G���۹$�pL<Q�}�������I|6EE��.9W+�ads���!#�vs���z�Ⴚ��BMխ�&�@\hLFUe	�������3�l�蒑D�����˽�\���)�$�?شuY���Ġa��O(P]�-`����Lx]�{���5=��I]@��E��Dm���F���i,�P6D|���	�%q.ྒ9�D�h{:�'GY	�ad�%-�CcN��~z@>��i�R�%��C����G��K�+b�#��$�B�U��<�~��_���%cw2/��!�:PG$�'���`��f��t ]ڗ���y�l{I"� .�a1��G��\Cy��I�2�s+���3���s��4�³��� =�8r�Ęlrq��T'�r3|t���@�fx��'�[a�)��D!��+o�Aa��#���C�}�F�	�e���B"�L�{�d5��	��ࠃߙ�$�%弉���6O�K��C���m��<�`���FG��&� V����tw��c�mȭ���'�ta�QC��`��&"U�}�	�K����(�}/Vip�o����B}5?��~����* ���ݘ���K�*Ns���ػ�y���U�V1�6����{�;86t.캻#3��[���/�6yW�<��V��k0�Z�cxm�,;�o�@%��&���3>����7=ã���� u6s+ʴ�������[F�@�tǛ�q�.Ek�䎡��I�|x&���pY��Dk���a6����ַ�g�`Ik����L��S�(ou���u/I��,��n���������K��R���A5�}g��H_�=2`΁�x�2�"��p����`H��.a[C�����j�i�/}��i�$��❻N�j�u����"��i�Y7�wVԨ�������ք��O�f�?�s�|�o��\���|3�
���L���2ѳv$�@&"e���}�H	��>䍏�{��R�Z.��EQ<�C h�:9��sͧ�����u��X%��d�T�^ɽ�x��e��w�ߌ��tL2�,>߮*:#� ��Bv�����St�O�dtfz��;vw���̸���.�z���&����b+��u���[ti�� f�zjώV���@:u���b��q���F�}Tv7Խ�爂	�Y��ݜj�|��?�*L�OVE�'p�KpR��&�C���A;q��1���?RGU��rR*k�=��<4V�b5�x��C	�-��bI��&�֥u������UJ.�a�~<��3�9�e2�aFmW��2��Ivf�ld9Y�V:�~�����>��6���?�ִ�󻰨�	�"�>k9�	�-&'M'��y�3�����w֋�g���-yCk���Jy3RD�P��ս�#��d9��`\mB5\��g�&��ߜ���?�`uf��O6�������� �̽�j�_4��ru��tD����q��p6fu��/Œ�CVZo1fm|���[l'!�x�>���(k����P1�u:�G�X�
��y �u"�����!Z��s��,���P5�~�5؄�<\R���y�n���!_�����(e��4G�l�I�C�Kt����
��NA��'�n�����H&�K�*���#E[���:4�CU,�ӟR��,}�O��ߔ�w��Dw�td��9���W����X�-��7h�j�|�m��we�u�3����0+U���l����K-ZQ��f9!aO��M3CV����ͥTPxc�YI�ƛgt��U>���^�S�K�-��N�8v9�-v����d�$��'�~=�=���2� �O�	X㋯�l��މm�k�V*�?�6T���P���6f��`g�닠����0H����U��R�dKx"~�5�����Bl�4?�mc�;m{��2���F#�IT���W8��y|\�L8leʋ""w�nϥ�j[K��k��[��cfߵ5C�h�Ɇ�։�ſ����]b����Ǟ��?�����.5±AcM�S�m⊺ۺ��~{ �CL[�����_� 8�H��ج,�×1e�дBU/L���]�16r�86��������͔!�ە�k�2c�N�����UVp�[��fr&~ܙ����^��܂_��4�N�YI����������F�