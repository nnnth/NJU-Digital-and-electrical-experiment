��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t؍�^��FY`�&�o���9h�rR���~/� �s�s�7�j:OY26JC��;�Q���3���t��&d�Hj�AsO>i!�$ �Ϊ�tq�k̏��S�I�2M���Qp�6l&�!;9$25���{Յ�=�Ңr���ٌ�dV�*	��~�U����Z�{�*��Y[V^�G�au�+�
�,�&��"|iV[�|�z��<î�]�;�)s��'�Z+|E$�5�e��Mt�۟���*�݅Kx���T�О����x��iyE}�#�]� ɶ��D�l
�'��;�2$��z����Jw�<�p��lx���b���K/�'��ӇS�5;�	T,��rb�u�/��fqOw�.%�$h+R��.!�m��_Me�ٍp��Ը����=����{xj g�"��y<O�M]A�Kh!f�yyWj5�%��"�0&I�F��xVt3��Z��x�!���x{�|��QQ��i*˘[%�v:%􉅇�[E������' �5����/�G��}���5�����U쁶.NIc����������6�wY���%</�%G�S+@Έ�zx�cn��z[I!�bה���30CR�l6�B�l|�-�fN���at�D~D�`��ʽUE�QM�җ���02�@��^ZK����,�7��ŸӰc��!cE�(J[Q���&G��s����5
�.2��=��Ek�Ta0hD����ӱ���^*������	d�������](s��@�j&a'_�?���-Ui��]�RK|jt_�B$ne'���&O�?0�q$�/��q8TL*�h5	��3E���Lk��qm�i������q�P���Z�cc²����t�+�t�Im�e5ŵe��X)	\��bi��aɉ
f��@m����)VC�/5�Z��9���ݩ�����F{OL�{4�Kx�}��d�L^�CO;����3�ܯ�,Ak�v��s&�Ma��]����]~q�I 	v���遽�y�j�������0o�N[�rxg�Q)b���'$9�{�+[��J����$�Sα�j�K��TM�~�Gr�{��<�&��"j���i3�tL$ #>��i�S�E��+��1�s�ą�o��̽eU�CkQ���ta��nLҵߢv�%G7#��,_"ͯ&Sm�ǂ+�óp�Y��c���bv=�h��n@ P1t!�����+��I�E/�]���P��v|�VW0��C�E՚tc�.�Eh@{�g6�YT��d��%<	�D>j�H��j��*֮��y+���},^�m�����tF�Da�n���Ish<v��w�&�$��0
�զ�3�����F�ίw�?E�d����h��D�n�0?*�AE3Ӵ�[�rЌ�R�k�7��ů��H��g�gU����m��+p��-� ���=�g�K2��s���)�_� u��tВ���$�A1<��.p�h8��M�c$LEn;����IA)�]lF���N$�DN-y^w�C@���s1��8e0����[�U�Lz@��Ԍ��=\!)�6�-㧤�Ώ禽�¹��J"��Sh�ܶ+tma!ُ7�x��f~�Z�n.�L~(�`�^�s��Q����&� ��6��C,�+\�8Q�B��;l�@ y�P�E�o�D�*��z��[���4H�n���W���"���Q&�:;�@�O"y����x��׸�0a��6EW��k��\ �oy�ӌ�`=�T=ƻ,