��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������Z��B��Z����eS��D���Kg��
A�N�(�a��Q�n��U��N!8ߎ`ۼ<-:[�t1 �m��PN��߭J�]�V3E@m���nf��,rﲴ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��90 �+F"��R��ޒ��9�#-R���xL�c�F�p��k}]�U�!�W|m70����aˬ$�ɒo4NU��y���Y�&#��/v��cPƇmjW���9|S�7�XX[L����vN}��*0J &���7&`]�<��| y����F�r��P��F5[��x<^��=g�.:D$kg�V|����2�bٌ�G�=���L��e�]ȣ����[��n���r��m�O7�B�#�`\yO�1ld�5����iV�W��ŝw�u�}R����6��h��e�"{�+�ū�*����@rJ��<�g��~�A�	ya'�#c�G��!dk�]�p��Gr�0�)�;�k�/O�p�\i⸬|6�8a0N�y��p��c,�V��S�c/q'��D��)�3�U�!�q���N+* W+5���^�e�
}���t��i*�R�?���nB�f@#�T�����TN?�~�ڏ�՚�@�.,�G3�_
��F6%�4�O ��oG.��d�Mt�h�j�(�0����y�`�Iq�Ī�\���O�z��0z��C�L�3.WEe�vO��7+Z��߱�:�g�8n.�HS?i�xBT'I����[.��	���d�m,�8��f��k�?������:��U߃�������ck��aq[<��/,6;����@�7��c��e�,��>+2fI�P�\� b��y�!�c�Y��G��p�S���cё4������Ɖd�;,�pYB2��E7���N�D�IH��*��/H�ʰɘ���Y_������3L��#'�X���T!��{�fSC�z��@��w��q�S.;� ��[��\�=�:%b$E�ۭha��JSq�����V�#m��:hgq�pD�%P��Eί�_q���%S�j�s���b�Su����Nu�(�ÝQ1vifp����T�h�YO�<���=��#�iLg����U�a����$���ߜUՃm �'���.|g����$�55��x��u�����$�i��F�F�D�R�իݿ:{�))�T�s՚e$�ȽyߗM��R_uݹ�hB}�8}�L
�~X�B�;n�S��ɭ��v�$�#wa62�ƫl)��OTb�L�{K�	r����)��ZrF��?z$�)��^XK���)��:,�I+���b���3�R+E-N����tЋ�Gn���آRi���Ko`�zf|��K(x�tS�þ�QS�X%�O�~���ϓՈO�Xi.�;Z�U��W���;�@����@�����s|�0�Ü�H�'9s�,Y�5J%-yD�p+=Bz�' ��4�G҈�"�D(Z8�TcN��D�Y� �UJI�8��$
�Ѿ�X4T`7���Q�2%���a��qc�0P+i����?,�l�k�����B͕�saϵ��"[�u�����N�*�:�H�ߵ����T$U����bt�����Y݄'�᪇v~=N �Q�؆n�\�r�Xaw��>d�L��=��ih��VM�֤��p��EA�7r�%��!8�Y�M�9s<��|�d�/�v�K�c~�7s*�sQ6��uk��ix���v�]7;k��ꊌ��k��pe�$6�\���dE�	�"���RYS���С|4l��B�[$�c�o@Ք>���BH<R �Zchx�Q�+�Mя��]\ �l�Z/�j6òڛW�<�Kw)��u�k鄉֫������8���
ȉ�E��U�*h�CU��ik��7l,�T_�{) ������	��:�zZn�"'έ�Y��(uZh�P?�\y�p���-�k���r2�k9CFcl̠]��Gi�1����ӂU2����U A\G�������O�%���m����{���!,s�qı�)�:_��*��W�����L�PJ�I��=�Φ4Uc�����.����#���w<?����F�W�9E����=�Li�s=m�/�X����b�ZH5lL��������HŎK؇.9`UÔmE?��� �{��HUwT�����#�4O� �$'�~f�����A���݁E��!�8�g��ߵ� '+�~�,�F��U6v2c��j'B����Kf*�T?��1&%�o O�u!��M,k�}�Ιe�stY�P7~+��i���s
��jE����A�����0�E*5�R��YR��ƨ�x�ƍ�~�p]Ԉbš�9O������j`��g=N�K f�����\#&�V	~�������ײ�|@�8e�YNYԥ[?;NJT�[-��anC?��nL"��Y��8뫳���f�5}�(I������z[�����e�Z^`����5�
p}7�����#8�V�0��_5��9E�.��%�X@uҐ��jvyZ�G�9�/��_�#��&�N�0FI�K���+:h�.���?K�tU�֞����-2�!Y�_��9��C� Kv�����qQ�`��N�����q&���&�I�����^p�4IuxTV�j�޾����
���=y'��;N\��K���m��g%���Oyv#�u�H����
��q8o�S�ނ3�n�d���)��5G�lxY���u�I��>F&��_�2�D]����"^��D��>�@��G�7hЫN�x_�:{z���K������5�#?|I]� ��#����`�D�K%(�'�����e6�V�g���6�D�+�H���p0)�L╫���\�\tF<����Ȧ,������HdEV��D��$�o
�m$N�� �*-!w���k@�r��Q�,{�>SP?��R�	8�1+�
͆k��kJg�}�֑��v/�뵏�%{C
 ޻V(��M�ag�4+p���->�  �$����кĪ������	��R�>$�X�u��[��\e�(Q*���Yq���7Ԡ�4�N/���嗊L��R��4v��i��t���	0!ŗ'&}2����}��f�+�w�+c�������e.�V��C��F���qkѷ�Uۧ�,��L+
D��+3���̄_{��	����a����)�mQqx~�%R��?a~�ii���S�4�ΐ�!4+Uv(�Y��/�U`Zs� �!x�f!8�y�+t��p���Ԍ�tσ���?U����(0zݖ������%�����cLHH)��Z�D�訂�����d!�=�S�(�Idn��I��i�� 4��^�l��AG:z����3%�4�.<:]m�_j�a���]'AW��lVȈ;㓰��.m_$�@���#.A�c1_����/]B�j<S�p��+���W��І��$~��?���
\v&
�@*����#h�Uo�mtU:�R�;^㧆G�<a+ H��� q%���kƜ �JSdO{�b*��+0�� $.r0�8���/�`��wol��U|�R=�L_8W�ލh ,�;l�nCM�Fk�(���l�E]��f�Qr�:���xd�!�H��o��q��E��
N(M��q]k�Ddɲo�$�Q���C�+���J��z-���<F���%��;��7����7
�ȏb�&���q��[
V�� ��u��ZB;����3"����tG�˲�b�\���8��WW$1X�nHݭp��0���@�rIm��5KDD���v�/x�_!,=0](~�ǘ3�s�b���bH��>�ls�y���ڲ�����5���=��<Mh ��N@�[����}|�peQs(���g/R����1�~j�m�����N��Q@n�Z$/2��%�sQݘ�%�"By̑��_�M�$�3���Sw?�kP���e|=�֧��8���b8Ko��qZ��?���և���)�v�D�O}Sx2U��� P���߽sf�z:��u(�Ӂ��7���d�/�,�b�#X�}��6�]Z6e~�;H!��5X ��[��&�"N�PGX㉥�z�P��h��Y��)3��
�'�"
�`��'��Sy|9d,�Ӥ��"C��n��$Բ��C���R�Feٿ*�-g��ֿ'd�{�}x��{Я[vM�#��z.�Wc�oP��ǐ<ַ�خ2)GE ��^����ɲ���t'�����-�K�� G[WsU�a�a��o�9��iA$�"o��B�ᵎ1w��� EL65/n���-�>R�� ;SL�c]�H���Mpn�#��� )1��D�Ak�N�d;�� :�-��q�g(+�:݄�`��첦5��s���  �D��C��eY�M0�K�3[�|�Kj�JFH��`"&R;L2�S=9�e���ً��D�U|K���"�&`ߍ#"�k� 5/�fx]�ZI�͋K�~��T$�z��X���	dY�d8V��[O>�1�?�瀢�<i��^4�J�֓��E�۳����Nv(���UB�t��
���l9�&��J�p{{Q�z������moA�����߹���{{��~�u�CӒ ������l
�ctЁbTV�J�!����(�ä�˅Z&/�}b[�(���/48�@��9�AF6�Kn:�5ܶ1ň��jݝ�r&�i�*�\�)�@@_S˾ҬfB�.x���+��V[�ZQ5�4?z�`�W�f[�We�m"��Fbh����'�R#�RW��W��4�WgZx��L+�,1]��\5Q�fn� �����������=�
�(<�
��Y�bC:�($��ARP��>a��  6�}2�g�ߪ��Y�����T�_P���爴��qf�y#g;u���W��PB�l""zZ�#���@������ �VX1�Ɗ�H0E������$9�����%�nm�)3��)�(����;݄�+��TJ>��Pn���`k����ajs��O�69�`
��$I�������Uh��z���'"��>��v�j�h�Q��Y�me,��Q} �:[vC3�* -���4{i��87���&���T+b�&6l���!kG�PC̙^rE��P�r��dg���ob"������H�]�KX�����g�jr{I���@SJ�K�:a�ρ��Ҽ�\�Zn�D�Q��P��ڔkF�����{�ށ���t���:�t��A��\�p�i�6h�9�v�1Ѣ�ںo��=<KH���A����-]���7���m����Ç��g>�й��R&Tt�ail����?,z]t��F,���:��V���t��tpy9�e� �k���z5��i���/�~��z��|��xX>�M�xd㸮�W��-���>��׿o�]q����r���E�_ĳ�W΋��ph�[�~$*�O+�p��/D���ֻ{�~~�zh�z�S�^n�v`�N��<�m�:�M��f����Z#�F�1����8J-��
�{�í���Z�| \q\���@*wU��&����jH�Y���63<t�/����r`Bk�M������r�ھ�o��b]w�b�1��9I)�7
����k�0���Fq��t��I^�ץ��NF��1[�=�)Jp�R�#�iQv,E�R���b�ԟ���ܷq��x�L�fBB3mV񘀤�7U�?0ر�<bI�0C��Q���8��@F(�8��8!����?�{�S��m�¡4	�VGy�`����K!����A�hMOl�V���T�|���g�U��g$N�ݝz�9�F�C�ڙ�_~�?��#�:ܭ�K�K�Q\����c�.}����<8��"�Oai��j��ҳ��b�m~�����4�J�B�s�E*(��p~�am����'N焙KE��>]%�=k��SKM[��$ ��A�+�A�kO6Eg�G�9��@0& �/�"���	gC�NNb�j����A#�hS�:
��m��fN��Y�; F�v��h�g	2z%���O�r�H[�
���ӂB����Y����e�x��I��5���('���I�"���(hi#d��!g1����#U�矣��1.��k��cA�B�:�{a���B�c��/$g�H�w{IQ5�c&�&W���On(t����<��F�O��ǫG�ڎ����KI$e�O�m�㐤$��Ť����O@�Y�3��rbσ~'�hd��&P���i��1�{��9�T֓<��J�0i�MHa��7 ƳZC���2��Wv a3�\�>�-���iXt�dV@���1�?m���H��k�lX�w,�;X7�ј �'Y3��9�9���7�Y�J���
�>�<_�[+�hq �8=�U�k�޴�7����<9��S}H*��p�m#Ac�_b�כ^9��l�A�,��rY��S�Ĝ�h^�!I�c����j�]t�y��g��t6*n��z��=T��&Nj��N�+�;�_����.�Q;�z'��_�=��W�ǒ�5�Ќ�&q*� ��0q"��چr����$k~g��Ƙ�OV�T�ʵ��xX�1D��[�r\���-,�O����\o����O��K3ߦ %���+Y�̟wB�I��2�K�$�9���o�'��܀���\_hHKP����Y_h�H�
����L�,�|֒2`����c�������?@�;�Ϲ����L���t
�ˠ��
|�xQ�1 I�d;e�..+� � ����%��M���f�fҟ�\j���w[�Ǫ�>�~�a���s�#�`�֚,5�: �$�����8�R��T؞��YW4Į�nKA�V$���3��yBq^�̎g5v�=��8<���b |�&���n��v�j�[��f��$-y<i��5�j�5����2�)�4��t8�R�O����Z��ܠC��7�5G���|@5�w������Д'�ۡ��,��0*���O��#�9��u����Uت���y�]���xZjPrv�������E��Wށ��N��S2�էy�O��R9����[ɉzi�yD�oI��,�=�i��pD�_)���;����)OXUi �m���@)���g��b�����9\rw���y�i��ٸn�rSJ]w�����%� ��}w`�<�%���g{������K�|��k��ف�#zր�����/ֿ9�J������r��̃_+j�S}��. 1L���0���!��b����ib6�p�= d(�8�|�X,�F�ץ��mO�/�	���ƅ\�-Q @�ܽj���L�s��5�ǕV�
C]fNj?�}�UAe..I$�8���؉`���w�����TX�J�����[7}!�~Ox��J>������W�� *��\+�_�S82�1�S,(�����j:�Q(~V��h�cK���(�l9*S��J
��_�_��{&���;{KΪ ����zL�4k+r�"��D�R��D�#��;Du����4U;{g�eˉ�p��@`-�-d��G��q�[�䅓yj9~n<`gBO���X����ŀ��;C���|"cqv<<)��C@s<���,�B�\%چ\�Ҹg�R8'�����9���鮎�ءS7V�ٰ-�[�l =�i�61t���c�<fj�MՊ
�q$3P�P�-i���� J�Y���ċ��9Q#���q�&����������X��3�la������쒔��M{��n��%��+�}ξ�Y���X;q5c�l$�9��<Xa�
�џID��8��ľ�&�W�G�����jn�NAWY�ryZ�wr�����ILPV�&Pi���_*����R304AA�Rb1v�}��kڴ����L|[p9�"+�h�"&E��@e�e� �\��9�8�aG	�PL�(�H���Xt0�,��TẄʉ��u}�J�w٘��
@�~�u>	�ӫov@u�͵����)^]7`]��UT6Jm��`���Oq��q;9�PR�_�X�@�f�[�����J`9[�h����~�+�Ku�򫂬�bQq��y��� �����0L	���բF�����=�]	r\Ԥ���2���gO�Ɖ*0�N ׸37�7Lb4uj0��"��̌�@��1�"k�x�e���!��/�<q����÷hS�MQ����32"&4�`P�ծ���<7_2���N��Ǡ\	�(�]���B�>@�k|�� � ~���Ѡ�0F��Aӝ�c��9�~|�m_v,��^4g���� N��?��8r���1��[�ϼha;9]F л����N��/y�-<�[�Mv���r-}�j��a��[rWnjVF�oF���r������f=���?<mA���OL��5��ZD �s{(��LJ��ٶ������U���K�֍���|0[��>�v��4�\�ܭ��Ќ���ެ���R;^�)��wk(cܹ��g�l	��7�L��9�ϼ����ҥ���/�FM�0;z�����#��8J��d=�m�jܝ��y�k_3�a"H&-�fj�����1l������yvK����#�h�s?��nk���؊@Btfx��'����r�kc_��(I��Ԥ�ǇO�jqO�"�Fllf���?�L�D�Y<���e��~ 1�X'��/_	��"�׾=湭\V,��������_|��ᰵxiضR,����^���&(��\[�Nѧ��O�3�M6�<�_k]�4�+	W��&�׿<��xm���/���E�(Ϛ=��������|�𧦄S+�OΪ�ƺ��]�aSÑ�byT��4®�q�e�(�yu��>V_Z56�v=ڭv�H?�esQ|�`�+E��zɱ����rQ=�kC��������3N�2	�l������.:�����L�DɈm6����t�%[L؃�ؓ�#_����POa����Җ}�	 kL���KsE� ��7��7C�, �(K�`��jm����:��k�6ԘgP��TȜc�/�*���2�
Vx>6@���?�,�v�t�O9`��e<��WK/�xI�V�^0��R���ͩ�?������b}o����=SІv�W
S�Ŵ�ӳED "d�D\�9(q���>^i��HXP�H��qkh:zu�1�}d��+��H�9��̙�(<Nb��Z(�����bZ�$���z�wR&�i�i�t֓ڊ��[�%LU��~��*&�&04���?�2�ӖW�)�{򴪂D|�t�_��(����҆J�S|�;��]���f��Xtn��AS�0���,�����+�Nˌ�R~��N�O~������8�q�����_�"��K���H�I��`��ʥL>�10`<�AE���x,%�g�!�E#��g}��B/y!�挏�m�x��j�\��tz��u�t����wR��JV�㆚l��W�>���+��#����H�fz�r\Z�/Y� �m��଺P��7��m�p+��[�)�Pb�!�HJ�$V��Vk��q)���[C��Yl�BѸib�ҧ�(B�\t�3m�P�:K約��	��"��{>�kk僇Xq�(�ۚ{L�:���`��f��[h���A4��A��z�1�y6��J����I*o��g�fo؂��z
_[d��L�Zm��yj�b[��ǈ��8 �!)�=V�ђg8�)�p~�-���
�U�X�CA��<�n䚟��E�p-ʇ��В����q��KR��Qn,���LZ��bf���'�IM|6'ϼ��kPV*���%+#��r���j���6r�!���Qy��R|��3u��.3�n�2�nݦ@�^�U�{Փ���$v�����r&R,e��0�wD�.{��	Ĺ��!�~���{�ٌ�Z���9��f~c��S�~�-���j�8^���6��L{^� �e��ݡ���匊�;��N !]@�3Uesĳ�����k��l��4߬�ү���k]Ie�9Q$,�FSm7խ����`�~gtE�ׁ�֧'���)JU8ܕ&�lG�`�7��S��xN����j@Gbc��f
���9���h?�Yu�p���Xh�y=�rf	��m����׉��l���Tv�.�C��O<er�7v�s�ai'�Ì��<H- �����3���S�7�9r}d�C ^�,B|��P�����[�'Oཪ�rg ����O�>�~F�H�<�W�X<س:si7�U���z`%f����Vh�Um~Oʺ��(�T�P�!�e"啮A�BI�+��*���������KG��/Egψ��N�2l�S��1b�5��e�B���8<��ϳg�>����-�`	͹��v 2��{�?�=�ۙ������u;�Nz��h;���f\ �u��:x��)K��'ksx��p	-}�@�~N8���Y�5�rҫ����]VEԜ�5�?��c,��	�����Ϯd
~�܋��籋{�_f�H��Agb����iH�%�㸳�Wgf��Ȥ���6�v�lt�Ģ�U�{� q,b�zV�>ע�ݹ��y�� N�}��AJ�B��$/��`�])|��J��uzf���*�� ���LE݇L��Q��*�\�0���V,t�᡼�3��V����N"�;� %�x�*�oQ&��hֺ�.�z�ͨ1A�g�&�KS�vO�n+�nNd�U	�=��F�w��]Ҡ����\bC��R ��ki���Y�u�N�}�e%K�3t�u��A�:зj��ŜX�bS�\#��Y�ә4���������>��o����
h1L���Ɵ��x߫���K��-�5�Q��LA�����M�����T.��-|�(?S�V�f�vXFa�ܶ�a��e<ܩTMo}���k�3�GyR(!;�[5�h���Ap���V�G��n��)þ��_�2gF ��*��N"���H@:�-s�ʋ�iGC(q�c�v�Oݹ��	WmJ8���dk}p4�B'�!��11=p��DD�)g��K���'A�1�Nq��Ѓ$��a�qKM�@� ��[#��?�Z4/(*5��*��-�
VB��ȝ@�7�t�����׊��|��q��-�2`����`z�b�V��T�1��k��U,��ꩮ�]�)Hy����`�}ޤ2���Wkh���H���c�Q3V��}:��$�8 �@��o����CdP���ʑI�_oٽ��<���!�:|l�`����?��m�z��?�l�V�q��,�L�_
lgL�� �*�=��$���N��v�u��JdJ�^eC$b���נ�ף�|rc��48P߬�a;�	�u�[���{�{�N�j���ρ�l�G'��:����#׻���`YM�h>�ۋ��� ã�$A 5��S��i�$�Oǩ�w�0I6O��b.ȇ����10��%�'�����;����4��$�#��ci>-&���;�j.�fcP��+����j��yG�s1�a�[2�e	wV�O��7�(r�v��2�>�!��{:�B�1��;XDh�t1�/qI��?��@<���|"5SnR�e�}.ƱX��5�.�#��6�����WN���'=��XG��y�������y���W�u���eL��5�d�͠�4B�Rl��"�{^-��cub�^�Z��pvD����;�Jrꣅ�b����7��ю�!E^�h�%4s�4�P���~��|:�ѝ��ȇDN�[�x��>üߴ0=Մ�u�N�Rb����ek�]�_6e�BYy?8 #z�QV��>H���ǧ�Y\�`�M\s�і�?��9B���cӟM=O%���:;�+�������	�tPwI�s�N��au�{G�F�Y�.w(K��xS�����=��۩�L�T&ͦ\��Z�(�Y�V�� 6��LT�A-�x�C�d��PEJ{�,��YYLvQ���;��_C��Z��⣰2�����ɮd�2�B��z�i�z������gŨ9�����`��*^N�>�BCa�����qu��8#�y�BX���1��o�t���mp�!����KT�D���2��
�S��ة㰙��#�[w
 ���5@eF�P�d��[���0�y��\�P�Ǫ�y���� D��]�8�*>WK�Z�d2DU
Vby�d�5%����E=S�p�6������GK4c:�� ��+t��������Q����Ôt/���n�0�[\HN�s��5���r��7�ti�����R{��6<1*^���q�L��pg�2J_�����:S�ķҀ�L@�7�xp[���7	�����m'�r��d��LL��G�!�[���I)��DiX^��=�*(z�H\x���y c�Z���"qpLq���͇���������(���������&����<�����"��x����u�6�K�#�U�<!���(�eo�Z���P�����j�G&W.��������-]�w�ā5
�9�_!�����0%���<�=�Ԅ�W�Iؤi�����x#����`�VPy�~�����Q���!�YH�+Q�G�V��>j��?Bz����l������Q2K���>�17Ҥf��S?��*��)'�i�;0Ԧ���(�a�X�F�M/ϖ�C�>~	wY��$A[Fs!����+�6C/F��"ēdi�J��K���[6t�G]v��-q���H��nX�F ��E���A]�R���0D�	ؔF���RC�:Yz��a���t-��R>Z4\��T�"�k�आ�b^ps�=���&�(Ǚ�蚎�ӡ3��t�AU��S��i��ؿP��)�覵����''�E�\�vec�e���[#�{V��}.���-[_��p�Ѿ���;�K#�$$ET�u�Ԏ׸��n�J���v2���<�6?����d;;���[mj�.=b,�渘*�cN�6�M���C��E�_��2+��29t$g�\�/(�T3�oy��i�!]l�0�w���K��&3h�N��J�)=�yhc�{��W̏	���� ���'�X���hGoM�W�$����v�Yփ�*3�v7�\Lw�T?��D!�gg ��3_ύ�[���"}�M�����5t,fc�*C�>��Q��+�5D�r"1��#�f�|W>���JY?�}��VH=���0y�,�. Sb6-�s�03ޒ���0	�q���m���?�^P�N8N��t}�#R_��~�������]��&2�G`:���g��є��E=�rw7~�f<�/�j�l�E�L�C�� ꣅ���(u�qc]렪��x��N*���r`��p*�B(A���QƿIpN^ܪ���	8��S�� �-���B�;��h��(ǃb�d9Ή��@gokh{�J`����Ӂ�7Q��H��|�ۿ�E�fmc�֭�U���Zra�y��H=��]a�%<�j�p�D�ܻ_�s��ɏ]*���j���>���Q�tV,b����É:�(�?Ł�<r{�΢Z������ڮI~C0-ʥ
��,�$W�|Wg�Hv^�0�b�i�%b|��+��$�n"��2]��_�fY-�<$�P�͊��2�fPT�#�ȅ5#%�MY�s%��A��[�`�I��<e<m�<l��35n����<��խ���4Ȟ�NCˬ~�L�ET��X��vĤ;)6@���cxHr(�����|�A�(wK�Y���dhz�Ӗ�jX�L�oE�,��G���8��%h<�f��G��^-�O�B�]mz�%��Q*�A�.���a���-6��$��~ѿ~J��� ���n�g{���(/dj�@8�q������2����E���[z�-�d�m�=2�Q�C{�.���	��R����6]>�!2G:���&!��Y��֪8�R�|e�|ᮂ9M]V�LbƜ���Ʃ�9�)6z��Y��\/4;k�"4ע��Z)�B�����(&���E��ZG�
�*�����^C�e���g9�T�[��u[�j���G�-$�[۠p�7�z�EtH@�W�	`66YH�4�n�M�g&��\F�e�#��p�>�.íqbXM�d7!�obk��-r��گ}d�/&���msO��6���T
{�"�F'^#������
�n�l��sS�/ؖ��e:��*8'B��I}볙�x��I��Y���˰$���'�`�'��t�N��n�C�Lb<Fni3���y�N%�8�imH#���m���6�h��'?(�F��FI�V,G��cw6���'f�bA���	�b.L���>����"����	%�Q�b�L�1�v#�.o�{��D�ܓwT�f���uym��Lf�KRzzV�����ZR����G�#ż���c����x�3M'k�(N��u.� �Ȳ?�}�D�-�=�~"#w$���v\��W�a�16�Z{O���;_i�qx�G�
�]��2I*�+6�.$�!nH�N�#a��ɺ��I�P3��)6��5,��[� g�)�^;�If`�tB��߽@w [�"ۦEN9Q�!׌�m�oV�"�;�"��6B.�m�P1��|P/e)&�בMlx�ٌ���H�nP1�h�s�;o�m��9I�.����Ik�DX
S��Z乏��v.�!\����zpis��[[�'�ۧW�h�u&˸<lR�&�M�ˎ	��uTX�bAĵ����}�ѕA�����|܇��]�aRC_�h �a�NK�;�$�K=OOň%zb�r��ڏ2j?M50vo��`ڔZ������H��X���dr�`(����4Ce��rݬ6mD1GV������W�&4�\�T���T��3ID`8�,n�������6Cok�}����c��������3W 3�n`&��~��C�K���bLቋL+p���?Y �o�eC9��RO�xGI�x�vͶY�+M�\"j,`p �5��(��Ju"�3�H8�S�r������,��0�м����*y'���%��`�tcOA�@E2yE���L�g����:���N]7���3n_�Z׏q�~(���8����)6�,6��!�ʡP��4��Ԇ-��Z���G�Qwsf�yD��֣��q�U�^��:��F����W��G���HI��9 sH�j�
�Bkl�"��V�FR�O�6��Pp�W�����h���\3%yF�ʪBZ��'���D��I���+Ņ�8*��x��|{���GuPd��Xȣ���&��p�9��}��K/�&U�OjLR��ǅ�^c�9()���(}����'��?oD��^����j��M oE̝��7|��?��_^�����[_�G�{>OIfA߆b ��v_�P�����c��	x͸���.> ]����!��Й�4*Hb�P
TFQM�WP�����d�V?�P?��I�Cd� ��8)�ȣo��Q����P#%&'?����o٨P�_GT��`���(f�z�0�k���Uc�#M�h�<!��Z@&KKt]^����wer�i��,5Py�@���	_���:�%��]F�k�([ v��f��~�`���C���A����2�кL!�z��b����E5(=>t�J�ZV���	��Cݝr�:���]m^�Z�����6�~ ��4�?:Ed�=��J�#ܺ�J�b���8SkS]��ĝ��V⣊d1Ymۊ�u���F�x�g(���k���f�,���x �~=�(�p�F6��@}3��wF�x"�f����:�����P�|'�Bw��z�Zu��#��zZ��ΘI]FgAK�����؟���N�<EY���x,���$@ԿR	��p�u�1H�1+T~X�)j�D�t+]��V`��G��L��&�R�\1�K#"X��'��ka��s�\%�V�Τ�7�>%^G�����l��o�P#����"o1ę�K��Ƨ��.����W��;�km��~\��6�@H�u���!�	��3��5o�K�mcw�Rq���p����K�?�C�Z�έK	t�3�:��͡d�m��3AAdx��T�Cg1q�l�3z�>v�
��B)�.3�,Ҳ�n�)���Ƥ�Gn=��tE

�o�?\O��E��	��uҾͿ*#֑bw����KH��u�!�Ab��Q����X�_:�|�Iñ+K�!vp��@"h=���0.�v�2��zC�uU�}y�9��S�x�q��[DK�W(E/1�VAT�A+�|�F��@&�_�&����ꤢP3K�?��0/I�>�+�$�� �tM���/���g4������	��, �[�^;��b׼�m���q7�Y����~1bB0)ءF8ᤁ�X��f�ؾ�3����rSЈB���zt�fI%�@�m�o�E��& ��էŤ����u.è�K��:�)D�l�G�.tN�;Xq�n��؁��Wl����F ����+�8�ܣ��kD^��� 7�&���y�@�P
���L��g!��x_���@�z�nK<n��!G����H,����5�j�F��ۄ�6��,�<h�n���Ӻ�y���~�1@�o��8SNmOGc,��߫�߻�^x��ֆm���#IX��c��:����,sY�e$��ֈ3b�YF���m���<DQ�x5C����t,��K���o��.����̼qG�rRS�e�Ԅ�BQ��O��;�|��\TQP��<xks��fb`���a"��
]3և!P88���j'Ql�qa.�8�����3}(�ᤋB�
l=��s��[c?�'P���}Kr�����R[�-�eO~o�J���-es<����^]c�)�e�VH��(��D�� �"�� ����Q_3Bo]raGUb!���a�F��|
�LoI&:1׷B�A��*�(�|@<���V���	\m�ʡ�t��O�q�99}#��H ����	���z���I	�<|!�~���=�Wv���oI���	�n��ޫ[�� �2Ӡ4F��}�Zc� JR��3�v��\�.S�h-_�Ův���j�"�0���jk�*#��n��z�u����[Ōn�l�8��.j���x@m��(^ )ʂ�(�A�`ҋ%n�44\��,�n|CNl���3 �����9g+x�><�i��M �D Eʘ����\�"��_6�fB�l�]��¥��Ʌ˘S��Uw-�4�>��G)��\~d.� ���k}by�r��-��f���C4.�yK���ȼN�����kA���y�6C�<�:�&�0�����J���P�b_��5���eH�+m�N�uI���H�8�[wSW����Y��f��Nw��|���o,��q��AÙ�)��]���t8��a�����X+l>��KN�2���7�3�� ���TW:9#�8wF�s��9�J4��vW��	3s��CǭP{��L��\tu�*�I��~�����I��8��(�Z1F��ښ�?d�r(�<��2,Z��)C[+�C���=�[k���0�/3%���W��ɤ���I��Z����m����?O�P����c�����K�1��mv��Y{K���'���ws�C��ŏ�*ob�[�N,c&�	R�)���M~���J8{��Ϧ�F�B���2���=s6������ܟ�U3�4�t���,b|�'w3�����ݑ��o`w�oТ��Bᩯ��v?�b��F'��I�A�O��"�$��a�xH�RY�!����������?������P���G�<�mS�[Ǟ6ȕ���o\���9N1ܯ���:�]rP��3���g�*h��t4�����yn*L@?�"��Un��(Q�Oi栛g����̥~���Z�����J��뫃R��q�5�Jͦ�疌b���>��� Q�Ү��	L�P�Gߚ1���B���/���'�MI��b7��.|'lo�*| U��'�Z�I������(O|�=O��0$��!��?�g�=������Q7�0� ��e0f�I!@9���Y��"x�Ip�`ⓚ�/J�����X�2`���B-:��m������С�C�=l��q-!��5ކ�0��d�-�Zt��[��S�@vV|E�I���� �c)�4|c-l�OF��L��%#�S5��]u͡[0�M�'�KgǍxn�Ĥ��F�'���%��C�����d�~��Wj��;�����g�s�&6��mt�Z��>d����`V�6��v���C��_W'A�Rb:Zɓ:  ]V� ,��(�l�yY+D����q>�cc�����58XN���@��M�i��6J�j?�	s�EKρ���%�5s;i��n8��|�&���0 �ܞ�X^��L��v�X�ϖ��w{�Q�����݌��c�Ѡ�l�sd}[o�=�6�a�b�F���_+�K@ߒap�)m|@(0+�M=�F�`��:?����F��w�0!��	^�nj�]1vpY��ݏ9{����@���0���R��m-��d*�O����r_ MS�u)�'gĬjf�L�� �V�C�L�|��F�<�w�w�=�ר-S���)1C�SqK'��890_�>F�v�l/!me��Q�9�~�6rף�y@ZR�q�A%��<����P9��|�P5�hX��۽Q'b��Ϝ���h�xpE 4��k-�?Y�^�S��~��z�dV)$�aM>�a�J��i����ҭ[8�:�э�B�ccd>�t�e�9�|��������A��,>�q��9�P�-\�
h��wF�Ô�l�̿^84��`�c�q��ơ�i�VʧD��^E��v#����&�8���Ť����W����E�-JY���Bw�tBW��_I�9AG�xa�[�ƅᓬ6uߒ̗7̎i6�-����_u��Ё�S��y��,�����@+�hS�fԳt<��B��[�Cn�*��� ����	k�c[��7�"F˩�c��-����p�@�al/ٖ��J�M.��|�L�9lT��pX�'_x,E=�
���JyVe���ل��'ptg��@L�B?��� ��?�<����Y���yQ	�j���^�������z���u_�v��S���i�$�3i%G��
͚��UPxA�C5Cs�²I������f�i�Q�D��r�\=�ޓ[����ES�pSEzpر�15�X�zwpr��Q�vg�¢���]^�����!JաK.?u`۟����}aˎ��ŁV`/��=�.�MW7�i Й#7�x=<t��0\ �z�v���K�9��%�N���(��A���b�*��_y��o|G�v��T�4b��C��MK��=+�!�b��ۍ�$�M�w�A:s(�6��K���.�0��N~Ź��$h�B'(�^g���Q�?W�xq��F�:��Q-�������h���P��In��C�q"F윀��|�՚������X�!�$&��*7���D͈�?���K%,��־����/Z�Z"Ҍeս!Y�Ns���q����v�WST�=���q�B�&����� D3H��G��k����`:xK�VѰЅ��_�&Z\y����K�d�=U7�ew��N�P���^�c� z��t�	�R�T3̲y��<�ڎք�Wpj���J�ĝz��d�.H��_#�=��Hϳ�z��7q���L��M��WfK�{��CXp����NN�SU �_xxZ(�-������a*[f2������f�ti~������~C���8j'�^��(!��6� �&Fx�D� 6=���-7�Í{��P.��;O�˂z+8/���!����h$�ra�,AYy��npVr���6L�C�r�R���>�q�b!��촂�i�ơl�� ��4��V�
��y�w�G8��,*���-rٕ��(���9~��\C��_g*���^��i}ф%ҳ���X��"�J�C�~&-t�5��#xѤ#%&�U������J��$i@sg�����������Dh��ci� ~8�H�+[(\]A�7,�#(�,��ǥs#��#����\�5(!�X�i.�bj�(���a~L�Fj΋��������� -�}W�����=�M�(T�S޳Q�s��"�m3EU�+�غ�28��\Gsqᶇh�.zd�^{Ҁ
򝽸t�a/�	� w' ���B�"�׳t�
�4���'���Stf�W@f	I�^�aB��T+��VA%繉��>fz4����9��~|/@Vh�g"{Aq�$�7���E��(��M'CZ+ǷS��ڳ��JI�� 2Y���Ŧ#��@��mj�v�E�ɀ��`~W%��Bp.�\��TH��Y��F�$����36o�'.T���w��eak!t�cG<"(����M��6�З���[4�|0MC~�
!�mG�P�դ��Ρ�>�s����j{vd��H<�)�X8A�L!�$��Za��E�(���D�l�ܴ1=�j;���!P�O��Mi_?x���]�Z��.���+er5��$b�M*"mݩ�O>�p4&���t^��&�F����]���P��|�:k��]� PAE�7��Tvޜ�I���>
؋ �b=���h��v	u�h�X����7�	��-!�B��(< �%�K��BV� h:,oc�|$���:N�����M�Q3�D�[�}�ܬ�x"J�S�iG��n�4A�n~�.Zr�>F�����xN�h��jt�K,Y!QV>G�ƶT����2MC����;޺�3J�F1D�v���&DeS `
!�x��&�e�)�3P�!ti�������^�ol�u�Z<M�J��,0[��<��$��7�1�?�B����؃�,�ұ!��ᩴ������ �\�|������� jͮ��YVB/�bn�K+~4��f��ICBV"��"mP]]������W)�䟋<�H�K@F��e�\�.w9ʢ��ؖ6�f�1	�s��Q�f���V����S��]�K�U5�}k�(���} �K/�\4'D�ˉS1���)��ZH*Z���6��:6/-m����x�S��й���A�8*|Ơ�	�k!b9r}�S
�kRy�Y��:5�@$�
M]pݝ*��t+��l9D���#�?�߲"�<�w>HCW&��2��`(#y��!0Pvڜ������#�吵4���T�`㟛 ��4Ic�U1��"�l����/�V��):�r��o��K'�=���5-�*��m��a���:�@ˊ�5E��������h��{1�w��~@M,�$x�ُ~B �oT̏���0+
��Ո�_�`���M�2�5��7q�r�z	��pb��|�~t����p���#+�/W�@:�wG�U���J��?��|���h3|�UӲg�ߚ1�O%c�Oe�l�V�pCfQ�Q)��*�.-�pe1��ls�2+fX��O�<C=����d�<(���U�*` �g���'!�	�Ri��nFY�D�ps�s�� ��yf�Z���O����T���a)-jI�s�z�x�A.$0Rś<�-bff�[{[#WZ4�ĴE�R�q�H�gB�҉\9�B
(>��ȓ{�V�e8\��K�Gm�5%�P���G��)W�>�'�I]�A�n^�]�'���o۬D��c��N�c6v���b���(wє�3��i��LX�6�Dő�/�h����B)D�{��?����G��	��K�{�8'�4բCz>q��ٿ�� e�nk��l+*x8��姯6�)5-�9qulF��Kh��!���R�L�q���NO�/�6���9�V�m(�p�Sّ٩'F��8_�O5�M�j�/e���O�<�<�3B�7N���u!N��U]�,$ts��YD"N:���#�/�kY��֞HT�gX���g(�"�s{�&s*�k 㥵"��\KQ?6N%�^=F�� ,Z��*�����b,��t�& 6��������`jS���j\�'��W�7��,�y��C���k�����Z�%";�)�r>څ8���g�_YL��v�	�	�&f�������"�������jL��vr�����Rj�|kE��M�I��T��� BI��5�����GCE����M}d���H�&���hJ)�kuk].�4�Jq�ꔜR=��e@�ǻo/b}s�$��=�Z�+Ҕ��%���:񓘟F����p�u���>��7�G*���x7�Aԃ�M�c�����Ԙrm�������e(��C
��1�s@�v7ǯ�����Q��Y��Z1�)w�%os���1��m�QΑ�i8�v��-L�!qb�3��+p�g
	���0�Xk��j�� �Bn�������:_���nv��6@�����X&jP��3�.��)˟��9kh)�)���sSc���ZP����:6&��r�U�Wo����t湵ԓ߮J�����puq�ɾ��E}C�?��Q<
�k�ކ��F�u��RW���&���n����8�N�ߩ9/g�a�KZ��;I�˕7�u��	���v_��{WC��sg7OdW{�i � �Ή���NJ�bf�8��򢈙׵)s�fq��8QuC[�oLEg1O�]4�w�R�v>���9�����Qn�b��������+�j!�h�۞�$6U�,#�ԑ(@�ܑ�=8��Q?m!Եfg&��}F˶*�����Ҍ�&��8�H��"?]o�N �š�X�M�"�'�z
C<��D���#sB���W�zpV�<�B{���ȅB�u�k��;ĉ���f�׀#��uO,�8��E�/m�쬆����D(zY�o���TiX!���|%b��Os�~S0��6�Ԏچf�{�X/��L��4�T� ^��}�	&�Q� ����zF�vK�B��"�\�S��P�h.*��r:�,[q�th��A�S�Ƃ�B��eǵޕs��k^:65��҅٣�=���g����H-8�2ܨ7���3����W�.;-���֢�
*Pn��K�������H�J��.[�^�6>��I����]bއ� �_h�~�]��4�aQ�*\L��}�uV�6^;�h�\|A~�n���>�rN�*}@��Q[����V 
g��	Ӏ�ؔu�������nʕ-x�Yί�\��Q�`�ˀɃ9��\��ɯ	���Lq r�[̊�����S�W����6'4.�QTH�=	f˥֡����eut���^��(����mb*����|�֣���c���<4�P�8F��� �.;�m�yF ��3_��R\�����[��,�2䇙��@�b�v��sv�v�+�Nn�w������Ã:F{�v�5�{�zg�>�}��b���T�D~&�(C?��k�
�����tt���݋�8L�S���X��a>�na�-�:���MS��,��v<�c�aco�]*�����@���`R�W]��]��w��z��'��b�5�ܐ��!�>���ž¦ocv����|WՎ^�z�)llM��'�z�����8��l�qU���3���Hv}��ΏM�9��@��;"�� #Հ�7����B� %�nxP�����ˏ�	EN�������f���碔x(CI��)J���������(ђ��w*<o�����������U!�pO��aT��}]� w5��5uU�Ysiv/ď� ��n��1t*3>_�:[�\;��fK/-1iwP��G�� ��ݔ��@������FA�FL=$t~'��f�r�-MY��vc(pᬬ�8{B��I��)p,�̛��
{��]�;$q�����.;����m��F��O��t�<�/�O�*���`uhv?�(OB37��y�Ǚ���l��Khߙx>8���eZ��xJ�ٚ��l�OQ��� �(w�!�|o8^��ݧ�&�9��Mj��B�3�(d�˛*���$ >ぞ��_�A>�ۍ=s��XzÒ��ַ��I{e�X�Kĥp�R�ª��.��@�^�^M~�Ƥ��N�k��;�_�B�5$T2�#_���7�	L#
a$�`^��d**���4�L��{�Y���.���*��5�Ut0��? o���5ē�_�N��d����]|��F~
�ҏ��q�Z����H�l�p�p�z�ƝG����[��ӬT���EF�(|��h���󯛸5Rŉ���CwGZ��\�� wr���,=�W�"9E����r�\lP0x��.G+��t��E�%6(�$�~8�_K%��0�s���3�#\�s�����	��M���hy�t���&�y�Ș�=�)�6���(*_��9��R�4��h�Ӯ�9a��C���s�3�ʎR�^���	;g3�ZO�s�$�&&���d1�:����+L�\����5�H���lԔ<���
!�RA�B���ZC�����H�c�:�e'a=r��ԍ�wq"?��ۧ
��K��x)�yVU5W9�jm�b��&s��$�A9<ư5�/���_�L�:ٳ҈#�w�@1G���� 
�Ҏ��Z(Z�z�bO�mu�Հ�q,�C����=GuSe䧅S��e���y��Y1o/��Rn}S�`�&�y���h/���{� q�t�FV��Vic���[����+�?z�n���9¬������Pԁ����;��D�bI���*�u��|�~���ssl��.fl�=]8@V�z�c���#m�|y:e>�f�=&O�;�$> ��$�"Hesx�O�`�������� `��*��.�(oD�"5������D�[ca)���´$OB{9�Ө+��;A���4����v̀秽;�r���������J�R�lΏ��IG�ʈ�S���;�h��]��<�Ƶ���9\D5,aw���ד��3/��CL��i���C�q$pD ~��>�!���j�ŋ$޾i��@g��Ư�+-LН)��샄b�b����O\���&bL�3���!�)�
�9���#2�rN�@D��PK
T�84J�Vػ�T�����UM�/~��k�� mO>� �	�k�gʆ̱����5��_Ȼ�`}��ɍb��`�ܟF�̱b��~"6�|�� V2�ڼ���t:��151n�]S}�0�q`P1AP�G)%����M�x�[J�]��BE�GR�<���<ڋ������)0s���碃���YT*S/��Ȣ婾���{�:tbo�]��uZ�' Y�i
���O�y�&N4?�WeNISS7z����Y$�� n-^c�&�Z������>%r8
���6l��p���]�0�M1թBEzc����{��,�3(s �͆��5��y$*��Hy;����=�Y}1�����Ɲ�yl1�O8��7�s�'���&0x�҉���[��`;���!;& 5K2<�5E�ZKx[�;��"g���ZJ�����ݡ줸@�c�=��8���y�b=��l��O<Ϛp��c�N4Jcrv���2����qj{���J8h�%�D�����x�n�Y䚑bV�ގvk�CՔ|]�Maq0�>t�,�5x^"m� -����܌9�LLǦ��0��<�bl�I%C��~�tV���i�K���S�o�� k����)����y�ub�M���b�J���(ǪD�6;�i�h�s����UU�O)$�3=�r�܈_]��f�*�32���S+��V�]{PN�z��+��)��:y
j�/�-f�CI|e)VD	�4�r�"=ДŌ	�z��ذu�(���L@��\gԱ4d��[7"�Ԓj�E�����q�<LF�U��]世[�B�m����Ο���.`�"�;�.cjd2
��O��m�h/h�
���	38S]�>}�BB�������Tg?�}���)�9̐��������������vM~�lT�_g���Re�^֕��@���X�R�1����5�!$p�;�n�+{��]B6L�!Pt���U�T��>���U�1ui�`�M����3���n�.8�fZ��}�m=a���T+���#�����q�"�h�-ed�_�YA��ڧM��nI�&�x�ǦG���l�k�]0�eķ�h�jl��)ivw�U�ĊM�t"��t���vo����n�s�-.��-y mv�����w���v�p����_�_B�#3��a����S��9���T��N�ɣ.#�g�t�0��3��3/��Ḿ=�G�?���t�%K����=��E��%�.˲��>�)ۂQ��k�K�C�.\)]��x=�	�K<)$-2�J� ���:�-"
�>M�w3~=�B�Y]{���]�XP��f�u�°�߱a��&qq.iXX�״N��f��cs��@�e�P�7��nX"_h� T�x{(O"o0�d���:�@)��rC96���R}(=Ϣa���Q(�l��N�5m_Fө�����$� ����A.֐�̏ �,-q߈Y� y-򦫼�xU�{�0`U*��H�ol�#�4ם;V�¢8�%��Y�.�i��"���(19��aB��[��\�u�W�r����ow��K���l�=�7�l��v��̫'�$�o�.���P<�9֭������ 1��p�������z�\quB�������s�%���Nc\���(�����T����W� h��-��J"U����HM�ފGfTY��b�I�8��B�0���S�T��ZTg��T��=���Wwȯ��3Bʵ��C��S��X-����vg�G��?�0EG3��"�i�(�J���q��K0w�s��R��T.���Ĭ�F:�؉\�7K0�̅ڗ�X�S��?��bЅl�Qbʉ)?l�e'�ߊ���ADy���;,��c��*���{[<a{J�q]/�ݑ���U:��=��g�8��/k#[�h�X�W�RT�:��͚����"��ۧ�z�Vb��P���GkI���A|�Pz2�VQB�B�#n���4mvZ�Kz|�Sv���$�6��{�7�SD��;(����O�n���9��/$R�f:kx�l������v�:��d�;��,mNl����N�@�@�8�-\ϝ��@��r(IV��-�g���毇������Dg.�tG{k���P.^�������#a��p��;a�)�4K�gP�ג �(�ߥ)��YU��++1�ñ�Zp_]����/�6*�v��
|�4�Pro��l ��Q2CT�����rZ9h�#��͆w��L>7����F�]�!'�(�c�#L;���]�L��,�M��������|��*]���U��u�i�Z��u��'�[쑛4������~�}���t�Q�{t���[��_5�\�Œ(��槞�ưG���S�����|�P�[6�|o��LEl5i.:�פ������~��<Ϝ�8}��d�Z�wq��*e+0xc����_V��젲EŸ�՗T_��*�� ���F@e�{4s��<�"�D�yӁk�8��p2��C��Q ��R<�"��K�M�*x_��{�R�8����am�
� Ĥ��]�c§��s�lT�L�.�j�cs�$�,���_V$�S��ὀ���ػ��`y�pAT:>�mH;VeݲIBm{]w�GRq�����_m݊�}�+'�I�L^SO]�Dz.zf���CSOr�τ�l�4�ګ�KN��I�/4�=�����+ݴ"9�����:%=�]�y�g���c�k��;��W�b��|e�`�B*�
9���t�ۮv^�𪳵�,Sˉ��������X}�0�������HQ��!�'�_D��ZWх��91��b�ۄcv�g<��r�M&��Hg�����U� &��Y���t�;Hٔ>�8w��+�M �kid/sQ�v���=P�����1U?5�}�5�|��Ѡ4)����_}��ge5*�i �N�#HTcOϹ����ǥF��.I�5r<��v)�~޷ � Ռ�F	T�#q!J1�m���z,��A�H���a<h��5,BF7�u��I9�4�E�~N.��I�%��h�TV"�K����ً+[q%�lꗈ$Ɵ�&N�ꁙV�T�����< |�zG�1��/�ʼ;���.�O��ʯ__��Q�ڌ���z�?����9;b��Grl*���.&��Ѝ�u���9
��֢�_0����A�>ڨSM�ޤ:���H��K����G�0�rV��č}�o�9L���B����?Fs��@*����s�	
T�J���2��&h6������2R?�Ultk^��5���FwY?���dˋ(>�W�9xH�vI �����L��tvs��#��G$7��e;���[�ǡ\?�,3/�&SiA�_���:��«}�w�#ϕ����&�O�LXߝA�8n*������RG����T�4H�U���I�냎$�Nۣ�c�����e�"�i�}:TZ��YnBet�(�D�PqǮ=�w�Z�DcA�cKSW��e�5̱H(¯�A0���ƨ�"`Ii�`�q�ml�ʺm?%Ѐgj�����#G�R8 ��@���cbaU*�o{�h�)��;�i3Iq��_-�Z�.��j�`��Q���/�ފ�����B�nﮑJД @|Ĝ�����g�g���OtŴ@-2�L5��,Til7,6Q^T�xꅶt"�����
,�B_(<�!O��z�a3��'j���^!̈́Ik���J	Բ��L�R~�[���J����E�P���#�C�FI�>Q0��� ���ޗGW����b>�/�O�5o�������LJ�>ˣd�T��­�.��2��SR�C�$���"����ȏ(�W?W�*b��=��P�C��c�!�%sS����Vb�+�ȵ7+g?_ W����SvO�\h�/$F��j5�_�H��hԬN����	��h�F�k�)����H��]��i�]�Ѐy�K��:��r�Q`��,�?6D��,�jO��������MP4=�g֪/���۷g���l居.����v����լ�#�
�u��6�J������S�A0�G��l-��`�?��8�E��0T�4��_\��2�������ؘ-����1�sBe�e��#�L�şjh��2ii��m_L9��"O`�����`�))R�ߧ�Jn$�v�} M��w_����g'�����T ��Gۦ�5��GEGaQ���C�������!�Ry�q*؃��N��3�PH��;<# 3�7�k�9���������e �H�B(�5��A��h/3�w����əy�u����@#�Zn1�<tDL]h"+���VT�����
�ƻ��3S���2�:=���Ϻ8��$�.��$d�^����8N�Re��k���u�n�`�H��=�}���G�&!t��`	��[3�Y�U�4�i�!{�e��=���]Ї|O��*Dwc��R�0C����O���\��z��D)M��'
��sZ�7�Հ|����^-_$i�Vn6�%4\�m.0"B��3��\�<�/7��hFq�k�?xN���~SR`��M�+r2�F2�R/�/`g �/���1�k�������lnE�8A�p C����)�(�L�:�e]ы�D���8D��R�W��t]���"�[�d�%��K=��ԫ�c�;
�`�]��1/����"�n:UL<�N]V9��[��F��2]�����>��G��P�NϙW�� В��x6l|���xvY������ݩ�.����_�Q�/��W5z�4���B��'��U`�ϒ������,Z�ϫݱ��Ŵ����@����:rV��%/��X��$�YZ-I�k@����`f��&ֻ-������_�&�������6&`�Ƅ>��Lc �:��Q$��.)P�h�'�# ��ְ3�×�7*z�n,	I��8�G�>��E�������~����ƿ�9Ҧg���h ��76�U�8����>�-BH��4x�P�6��XA�hBb����<��+7�ow��?���6`J���p�l��~����Q���G����?u����E�����8��߆w:��8�������;���c@C�j0��]�Q/��>Kh���������?V�f�'1/-/�X����Ħ�Ê�5~���GTw33t�z��
�����s� ��
ET�������y|�/g��)��V��������F����z˦ﹳ�ȑQ�s �K��VJ���^�
�Cr��%���������֯��ʖ	�l?� W�n]t���5���&���0�,/��1�ݭo��J�hY�6�{�J�<�?i7t�-� (L�"| ��R�'bt������0�>���/��Jr�w�w�� dd��O>��=�#>�-b����q��2dKBQ}�ܤs�~�p|��\�%��qZA���vAQ4��G�:D��.�L�L'�r�>��[<�Ϊ#��|�V�u��D�j'�d1X���X��l�
�C��<G+�W�����0T���F�A��{�dv*��j}����;�r#p;ؤ����aj V�"h]�|-i$��G�����D��A�|6Վ�6�Z?��5�$-'K?��P�gm=|���g�I/^*@h
Е�+�`��K*������I!��UnG���V�t��(H�R��M�Ψ�9�)h	bLaN�*��q�震�t^��vsؓr|��LaD�'�(����/��_��7/'�3���y���;�_��e�_^ q���b}�9:�����}.#@���QM�_t�T�q/[�a�����G*.��LQ?��I�S�bT�*T����1w
�A��Kh�'l$$|���i�s������O$��Ah�@��c3��pAu���!G�qKք��5c)�s1+��,��o���7�m-|h�}����q��ú�,Ǜ|9��*����'
�u��9��]@]��O=0��h[��'���Dh�okؔa���l!:�u��^�&[�s�똝�L|Vq�&�Hw�������G�pJ�}#�{ՙ?��VrV[8S2�����TZ9�F�J��i�r�uv>�� �U;������# ]J{����E(Т��Jܯ�~q�ՌQv��< r�Ţ?Ҝ¨�NA�����L�OP��&dV����X��d���"嶗��L�Q��j�<�x��zK3V���3���G�@EF�<�{+�$\oi�Z��
m�z��6�ڰ�[eSQ��.2�䨙���P)T��l����!�i���4<KP\
+�6�׎I���J�Go�����;��հ���
v(�� ��l�����D�o����>�z���^����n�$��G� F7�r!\�͹_J�> w���?O�3S�)o(��2	 ϧ��3b������a(�XC�Ż�;��!���[Gk��t����/QSCꊾ��H�1�ҩ��!���zQ59̒U��er���o��I	��)ϷS[�_��4SF�=��¶�U:g(�0��T�������U�Eb��?�ߎT�Ze�(��d�D���E�?�C���Ӣ�C�zxd�"�溈���rl��S��)(�%��C�� #B�G�H=�#�6��!����F<��#�z�^$O�قjQ+����s�w�K�h/�a΀�L�����&�e����Ƌ=:,�]�:�P*�A��֠���w�6N����+���P+ M����5��p���c�`���V���v�;Y,1dr���E��f�څH�����h�ĮE�t�1��Q3��ys�<���ӌ�G& �E�Z�N�DC���c��bЌ#�A#/�Q]cW�R\?�b�������*,��]c7�Ǣ�*�w�{P�ş>�辴�E�l0]q��xOؠ���������
h���ER��J�Ђ��7�c�w:��=��~���!�-A�Ǽ��ޛElEzT�I�(�xz��$O���2�֥&�f{���|��i�����A��@f��"�������io�̦�*��)Q �e�#�GY3�sf��4О����ُA
�ֶ��RB9��A�m��ݬ��(x�O/����]k��6�gUɅ�<��(*ڇCH�rf�g�m{i��sD��U#�K��qI ��� �g���+g�B6�����C��/��h�\����k=�s@�P�}%�Ujoj�K3�!���bvA(�j��j�2��;��EM[Ҕ9o�+Jdi.`�>�`E��ё9�>SJ>i��T��E������$��i��`%����p�\���􋴵��t��>�.��z�}ڧ�]�!8�����S�j�5��4�Y~mF>�Vo�Q��t����=�;���M�	�
��R�QZ΄�n��AJ4��j��@��.ո���;�4U"Su���[U#=���?�c+""1��ܓ5 %:�Gs�: �A-21��	���Kog�d�+!;}W���aa��։�*���ׅ4�ƝF(2����ٛ�#���/��|�LN�M!W�$Y�F�#�g�b�򁸇�^W���L��\<���Br�˔s���e�S*�BY����P�j�>$��FRw��_l���o����7� �rkl�����!��0-�WV����˶�*ޡ���
TUY�"��?�5�0�6z�����N�r��n~�`��6@b�a��_�.�v�7��R�(L�������5>��n�?��K�3�R{�B(G��!ǾFR��K	��;��#�pB/��ǅ@� ��쐯�8i)��ş	<N�(���$6�Mɏ����?��m�3갷}?�	�������~f�9����]��LM�����F���v��-˧Izo)Ɇ��3+3��Ll��q	�`�xkw��1�TK�@)��TɁ�)�;f�U8�[[�B*�u(��BǤ{���zM�_aO�i�����}T�w+�t���@hӯ$	�lb	�E$���:�Q�+��-N���?2e|q��D�Z�%'J��Q�_ߟu�9^�����|b��!0�~������q�C؏O��2X�~�h�<f���:UCZ�4PL���]#[v�X�
�ߕ�6�J�����Z+��г�V�ϼFWh$ŴD�GM��cJ�F�����l�4�E��~t)UѪ�V*�A��XM���-h�{�ϘB�nEғ�)`��lr0�k�HA�@X�J����6+�N�7GtV;�*��E�@EQ�$���)s���u?�������h�1�s�H�<��[�-�m3`\�����l��h�
�n�4b��mԩWƶg�NѴ�Ib��Qo %ɿ^ٿ�V¹�4)|�B��;0)C�7n�� �S� �X��0���U��|����*EB����#�*$�iX�t��st��%���8�΁�h��%����P�b[������8�NLQ���9Bu	ֹ���\��w��sq�$f�W�D_+�>�5������2��k�wbҜq%�������.��S��|s�{ɂ�Z�fVW��ĭ�+��ρϻ��}�����+��C�4:T=� �d�'�#NW�(. ���^���܊>"��n\��[�m�
N�fB!`ޑ=�=:�֖i	��D�D�����X.Q�p��$2<���Y8^�!���Z���]v�����G~�#�<�2��,�2 ȏ���V%{��4�x��A��L�҅��5�|qwp���K�8vqr*��;r��w��GbѲ��H��zx�$OZ��#�v������!�Ë�M���$��u$��x�j�LX�`t��� �_e�)(�"�0>������=�s�����������e���sP��װu.(�WX�5��{x����"0:��_��_v������Ͱ���������G
�Bq�T�?7�V��df���#��4�0�~�h"?V�Q	�9�[��镛����5�1��;�k(���fY�93<u�� �bJ���n$$�-�Z����ըq���N�Bg	��s5�Z��d�;c��}Z0*��FYD#֡��WC����ى��dPBF�n�8�%��M�Z�l%������q��MG���/'(���Bm��s����!OIX6
BHe�J�KyP�����S�������D"��vv��bA�WW\�����	�X$�I�?ՈS�ѱ� zX3u�ُg�����G���zKx:R+_�Hkds6��'2��.k�1����t��t����L'��݂.S3tu����"r��h���>>���J;��9)K�%��J����D���j���S���8��Y�X��j��3 ���Tץ�i! �[��P�y���L���;8�쌵���f�h�
�����Ȗ�|�Nz�����GZ�߻�3�l?���P9o�)���{�XL!�d�A�w����ج�c0��r	�BU��"���0D�NT�=٦�bۺ��!�9����F4���}3����Qզ+v��ҩ2�>�<�0S|��m{���m�i��Wҵ�n�0Ŵ3��Z�siУp�~�8�e�ʑU����Nkx���	qKe��"8�QbA_4'��[�PL�߉t��sb�?�ɿ�����L-������^��$#��O�fV|��l	Ar��V����CiwwB�<������?qQ���1k�=��[��P 9+κ���Pm�C�v���8��7��1Ɩ%�s�ir�^;!�LL;+<^|=���0R�CFO�̆S��ɛ04�F�JZY�S�w�2zDnѶ�.���O|q�$���H'Z�ln|Ц���4i�^����^d�Xl,� �ګ)0z�94�V=��1E5��۞��3ܤ��a]�O��Ӝ�	L�\���"p�_8/!�@���d��Bj���ٔ[bH^�%E�/q"ť�%���Ȯ6v�v�/1��K��Bf�U����1�P����i-{0�qHLH�h!D[?���d��p��p���)��(��Z<� <q騭�0;bX�	+^�|(�Дn`�ۖ�t�Әk�l�دs���l��HIA �CS���\Pg.,�2��mty�S���>�Z�R�C����F�Y	ud��O��>+�-���1�>`��K��J�-�x�Fb6��o��^�Q��3�>:�n��'�o���M�O-�B1�0�{�2讵��ze�טAC��d����ǎ�'ХG3U�����ɧ�e�]R��Z�a�-I�l�K��J�R����M� �QM��yX�ϡ�i3�菡��G�����'>'�\鵮V�j4���ԶV���"q����ŏ	��b"O�S{,��ySI*��m�`�Lkhg��������~Q�S��1�d��R~5���q5T�l��-�uV��9c����/�9�F���DC��\Mw���+3#�@����y��Wε�8����d��n��W�
+��j�D�B��8��B��.{��~ᚖB���y��]W��(ѓ-wو,��6���o��g�o���KӶCС�+_ ��`�uI���P%�4E�k#�MX{�>�.1��Ee'����'7�ғY�dǺ4�Î��DVIO�¤�Qdt{E&g͔�硧-��P|�����h�#6!ﰃz'��FN�����C�t����*F��w-�uz���J��,��D��~P��.�Q�,^�սҠ�#n,!O�vAD���*_��-�/&�u3�y����8`���
V��Oh�ת�'�)�A����o�$l����j	��FݗX�����_B�DhRrrt*_Qxlq&x���<ZƧ�G��'�v���=8��c��`0_[uP�E����Z���4Y|ّr,��YQ������@Z��]U���0����X�#h�̉�8&̔����Xwk>~�$�׃�Wy0כM�4��|lU�1��!yC�w\�<<�����5�SF�t@{�j��2�ցW�#�f��=��cU�})��`�	�|��k�aS)[���"v_Ijￗ>�L�%v��˞9w�hp^a��I����\�4��'�p��Շ���HS=K�r*k��`6��<)�rϺ����S�{�﹡�z?����{��)۶�VKz��hP(���I݇��Q��[�@s+�f�XК��P��Ā�G#��>�X�#�~���YJ��Ղؼx���������4.���4	� �=���x�j���!ġdP����~f;�q���$����Z��u��`Wi��3TN�����q�0���i�@��%YzB����h�f��`Uׅ�����7:ӝd7.:c�)([hY2C�i6�R"� p����\{0�T���i�'�c8�YV�=�nɒ㧫\�6`~;��"x���(@�g�o�Y���5��oH�~�5���jP�����m5��~\a~3Ӝ�l:��j'��U���,���oS�p��>W� ��:��R�,X,H'��)��⺼��Ƴs�r��1}i(�����D�����o�ُ��$�x�����@ܙ+���r<6����C���Z=2Y�@�8�l;!�_��9��7�5LF��`gCq2T�d�[��)��19�^�9��4���K������YK���d�v��RZJs�~`�Z�BR��6R�t�a����9C6���t���7�Ӕ�MM����>�.���p�\9����%����쇽8��Vj����+�Z������]{��]���j=����^FB~u;B\@�8]e�8��jX��8���F�ņ�/���[���F��M�2�/L�*�S����^�����L� �b^@v	�θ\�˱����D
��,�EH�ؕ ��s6O�dV��O���dgԞ�J���������Q��r0�	�*�nr�!����*�m+�?h�:��HƔ:,��J�Q��`��F=u����geѴQ��mDY�N���߻Wu�C��+x�AP�݂g�3[��u�0XK��;N��R{ꎴ�z'���{�Yh�t�&Zs�ų2K���������<�nY��+��R�����raaj�A��i��VI8��R�� !'x!�hX;Ŵ*�^;���]�X����H��$����LP��0\�E5��2^���x�Š*'�a��4�,8�8�3CЄ0˼&��5Xˌ ��;�=�ķ�(Џ'�R �ǕF�<�,}BGR\��*�͌eR���n	]f^�|���9z���	ͱ�*��]��:.1Z���Q�o���eC�ȃ /��X��:�iT���z#e<v�oi=���h�R�(q�uW�֩���9	��|�l{�&Go���˨�<Ɔ��rd�F�=�3Ekꢏ�/4J,�ڗ���h"�����+����?�v%5i��#B|��8w>���y�SR}(�ߠ�p���ؖ�����d*|�-"z�&��߻M���N�F���W��i�����	t�gG>B���ctX��3���!���:�p�z���Vl���^�vg%i��CZTgaQ>�H`��h����(�u ���G�}�\T�T�k�N�:����c�����Db�/,�z�7�	�٦m
�Ty�ɸ5.H��6��0��O�`n�N^wU"�7�?�k������z���u]�_��4�� �,A�"C�gҾ�ƯRw�Dþ�`�����;��r<��uc*Yf3���d���I�Jv��h��7әH��9�=�c�iL�y3���σ�z,o��ؒ��8ш��ַ�Xr<ϖ��lr���cn��<B�O�u�l���
<�B1�}j1�����	�$��xL�
g�H!^�Ӂ���Y�m�vyv�:��z�m"�s-0F$���\7��T���G��(rG�R,��ꌬj�Y��|�q�,��MX[�:y��H��\	�>0�#��Qzzy��f/;���35�!�t��=in�8Xi׶?J�����a=�s��;���p{$��4!�l�/�a9�ż �P��e9�V;���rEn���F	F�`���J���6�I 7e'6b�`�)�Cz�a�^� ����W��g�~�e�:���(c�y�pmQ���;��=��'���gS����1!u���E�0�XMvI�=E�T���h]�"����t�@?zpȈ�C���\���:ܳ��,�Fi���&DO��R	��;��"��$nu��%��	k��|<9BNh Xw����x���v���ǝį� ��
}���/q�sӍ�'�G���Bh���{��=��)n��b�F�&�n1_6� �����=��7�?hu������Yq��p�Oﹺ�L&�K�D�9TŉN��v觗xCP�|$��fɪ�Z�g�q�_����6�Ai���?/�Iڂm��X�S_N�����s֒�|�UP���<�nDt���/D(�p3(��}x	�/K�K�#n��-�3�^dF1���:��#_�f�åЈa�`�D� ߡ�}�L���7�d� �9�̶,�tֵ2�*���E�P�u�L0m���X����T�ZA>b&�����\PBM-ݱ����pwCX�:Kop��hf�`t�����X��_e��X|n0D�%h&2�Eެp�g���J+
��O���ϟ�ӶB�$sT���"Gm[�c�A�5,(�DY� <�$�i��g�A�Bue9&�W��Z��i,�3� ��5��L��T�b2\����W��Л�n���"\��V�[z9�l%7��w��y�0���^L8��p���h����_t�V��7�t:=�	���&о%��'����2�,�˅�>ɸ���!�YG\ Q�ݥ�Ś`{�@ ���>��91��y
R�:j.4�v��s=�E� d=�)z6i��4g�ܠ��v�P�ˁ?Q� ��h�ߡPG�Av�U����*�ᆙ���B�A��l�ц	C| }�m�k�Q������ex���R��D~lws�s
c������$��ӲCG�+�N".����f9�N���ҳ����'��@"&�{.tGBh���I��NŹ�k�z��&E�𔟘.��	��;����,���W��{�)�B��+�c�؏銰��|���Qh��4��u�'�Fk06H�$eq���m��t6��˄�[���JT�2�*�ؒ�Cg�����5�r `�{1Zs�Z�{�D�V���^G����$��^��_�X��/菛�����66���#��!"����O���z���H[y�zrh��1�/!I�=���m��:�-����7�`w���}Xg�Co����o���;D#K�q#��VE ��e�aDs��.��p�&U������%	�$ǲ�ȍN]hq��D$�C���GU��OH,D��{i-��ͪ�"KO�$R������ʵ��{tc����s�a�
0�OP���x�&7w	w���`S� ^.2+����$�vZ����`�������{PV�4H�fܲK���i�|��ĸP�g���mf��-��[�z�����x;D!�!<.pn޽�|:/���(�l`�ϳ���05j=X7l���vsnN�-��*�������A逥dH.�9b]}|oy�U)��K3vE��dV쎯���w#��g#!jnyߤ�)y��n�;"/���MGj���3"��=�c��Qmq|��X)����
�n�N�f�B��P�=vnJ�\��P�� ��+mȵ��%g�R�j;T�qO���s	C֞N���������*��Q��� ��*�?X�Y�;ޥ�V��dY�po;W�w���b���t;����8m��0~5�&��� ���L?4�6IE�9ߝ��m|���S�?��/�--��'�˙7ظ֪�t]���M�0�[��L�����mB8��%c/�o�T<���W�?�ݛ <:ax������OK�c1u�3\�ͱtE{��J�L�Qx�!��J^0N����
[�#s/��>�C��s�n���t%�!�I	��>gj���bOi�OŸ�����v��)3� Y�O���7�]{�}q�_��k�!�q�툤E��kl��CϏZ-�S��[�@�nݰIl؄)�2Ϸ�w�Ɓ��
��|�<�?m���otm�ߣ$;.|p��=�E�|�y�Mz�L.�lZח=��b��<<Y7��lN@�v����|<9�,Åȸ.̳��V���(w5Q߱��8<�+*!�*��T��G��f�v���=����O��`��gb����a@����X�)��:/C�B��E��~DQ]�}f0�����M3�\`�Z����E�(�H@��$�=�q>,Ǫt����B":�(�d,���M����TbG#ŷF�ܐٸ�i�؜��"�{D�Po:���c��0f�-�(Gf-�xP_2��~����|j���p��~��m�Xv��`�R�7g��	�T� ��shôw�Q(������}�!Ɗ{��r̶�Up[�ـ��D65zS`Y��D�^U�&$���Rz9;��)s�����j�d�X�*��r,�┡S25��2n�ծT���"��]zRMbHz8z ��K)�9h��z{'<��8�xvm���6�XXJO=7����[��y�VD�N�ؔ�St<7ݞ�*���2@�J��&H��Ke8�v��W��������#�(q�Όo���f&���(@k��@�՛���sK�;�����mT~�_�ҰiV���̶'��ϖLp��Y��Iv׻nB�z�J�=N����PZ�`GC�c`5PKh�`w5��;�IǬS���?W]%��։	r��g��}Q�^�ٕKa;�U��7�9n�W
K���4�ѻg���Q@���+s�J�k��U$S0ş�硷��[׶�2^�&AR��jO&�j��~�$Y�]������f������3I��
�b�H�=�O{<*k����ཽ�k��\���tlm���H1[o}�����X�����>
�w#rH�
��O�5�oK��ŷ߯tԮ�_SO�`̷�*Onw!	�D3���\��t��]��jt�R���A@`f4T�2������B���ǹ?ܣ�Ǚ��`�F��?d٩[�.�&�%}����0^���&���@����jG����(�.~(�a����w٣���tt�ң	�F[�-�Ӹ�^�И�52�t�(�[�yI�
[���03��V���-r�f�uQ��Hh��`UOh�I�(\���s̯�3j�XTʞ� x�.(!5s��nRNb�57���.ٯ��}��J�س<O��f(�+$�˅�߅"^����g���4�:f��׹e�����Y�j��]�$L㱊x(��_^�F ��ZG�����E|"]�+����.�ϾKZ�q��eq��hAhi��C�҇n�z;e:�\	�'x�bZ�C�#�p3�z�-��0L]��g�`�sU-�>�fHVn�W��j���*Շm��P�2Ө�H��@V����ad=�%0{�F�cOE�V-<�R��?�ڳ���x\�Usd�EJ�h���ߔWpu�7eJ���nK����q'��a����#�?B�G��,D�R4�z:�Wu�^�l�����󨌊B�o���\��b�������_�K��E>�'��׫	�ݐYa��gJ�������U���$ښ��_a�{,���+�6��ƺpcna,�aɥOۊ}0li4�k~��Xp�hUr���*���U�Q�
���vz�wI�%Z�ޘ�����u����^�^9��R%>c�زx��<�zeo���������88ܞhR������Q�7�Ą����Ե�Iܳ#"`%oq!=UT-0�^❄$X2��+R`�,���t�"?�I�+Q�C�k�w����� ���9�Uic�y�qT�A��d�<k�{<��t��B�瘚.l7bތB	F˝�)��-{`������YAz^Y��ދ���P?��o�A))ظ޻ 4L�M�R.q�?J�������'��������J�!nF1<��z��*w�#��j�c�+*�9/3�!���W�,o=C���v���^�ǎYQ�����@驒}�����������'?����҆���V��I鴷*�y*��1��j[��VR�s�[�aJ��D}��R:d�cF>Ue-y�#����MA~Lg�-��)R?N�n�Wʪ�"E��iB����p�sE����-3 ���@��}�K����*n��#U���X��u��9�f�g�LM��s����4�a����P�;\�&�q�4����"䈤��_;K��q��;0F������&����V5���#��jhR��ߪ�KW/����g�.���X�	��oc)}��L�K�Y�4� 	7��j6���}��،���j�Ց����1D]�Û���t��QY�2)�P�o"��8��;���oH{���,Pf�����;�w�ox;��KXzĻ�R�["������p&,f����`G%ϿC�+~���?�H��8SX�嘊1k8HH�-���*A�:�X3$]��;#ċ.G	)W}�n�&B�x�Y��ٌ6���� e�2f���K��_�nh��am��@k/U�����Z/�g��~�
ޕ��������� ��?A�k�P;
 '|%�)����^4I����E�}�g
���τ�P�qt�Z9�rw���u�.��0�=����پ�)�.����8.і~�%O6OӭM��C_J4s����}�ٵ���,�QIdH�c�����*s�t\��e����7� �*]��@zA��1	HFz��eD���Jo����,\$��qY���W���Ѥ��x����%~c\�쩴�p�R��yp�*����4���_�!�
���Ε|{������g`P���} ��=�	L���m���/73�đ"�'�9#&k� �'�<�5�y��z��l�
ݲ��: &��B����$&Z��b^|^��ۏ�O�r�q��s��C�I���N���P�r�%��Hv��wގJ��8��h{-����'�'<��V��pY�:��7}}� ��ev�Ϸ��j�@��׏ٍ�s��$5����=W�2�a%�%T�<�(��s��6pN&^�/�s�U���,G���D��Q
!{��[�^=�9��cZ��`�jEB	L^����&�;~�UB�A�!3'�mR�h�7�勛�����
�P��0�K.��QK����ɝ|h]f�}6��U_��Sѡ�A$ytX̏���a�����,���bz��(/�����1\�_L�ͦG��=��,�+'a�488���>,�Јh�t;�o��uu�V=f3/K۠�ѯ�#�Ѭ���B/�[�� �jnښ�3�F���؇��7	=.?����0���ɭ!�8�$��LHYp)�^��\�(�>��dr0��c���9�X�S�=[�c�b�����o��9��?i.�|	W{�H_�H<i�Te��	�n��}�~�-kg��f�ZiT�_�9��d(CC"�󴉁�k�3	n{�UZN|����I�p��Ӭ`ݯ��]��ap�Vg0����m������M�1��O�5�Nei_<d����H�=�曑洟
�-!2&�U�<���.^�)�=T�\:����a����I�Z0�O����(�ql �]�"�%'���w��+!;�ZT}��G� R8��G�
���$�H���YS�)��}�V�R�rڧi�4�<>�s�2&YH5��c��!%�4�]�F���LM" 	/��b�8�Pn�3�E�6B�]�ܲU��YcPl��#��T;�t���`�]��:�;���>/����Ա��=dRK���;P�6�؇U&ɕz�}�?���"���7R@2��ձd��,��i+
A��d�QT��dS�����H��2�����,E���q�#>���W�\�}'��P(wx��m����~"ַ5<`t�a����_���존��:|^?��窠�Y��d�|E
EP�CY��I��f�t3�Hx������}��s�]9^f�k�9����,*6{�������i5�	�i�;��2/�8	���8�-p,"?3��Csa�\l�T5�C������/��'����Xm?Ф�ڠ]�swD?���#�+i�т��?�Q��B��K���Ɖ�wve�w�!`O�7���9Q��`��8�F] Q���w9��,b��;�z #X��ɚ��Oy�g�H�;�~ɦ�1��@�vְ,N��Xy���ڸ٘Ҹ�����9b���:��1;�Z�ITv����K�aF��5���$���;G��L, B�%9��L�ꎘZ4����/3N�U_�'�3��0�`+E�Ќ�c��Z��ޔ-o�� ���1��?�'F1�Xq!0���F���\�~4��;\~3u�:k�(�6I�����������o�{�p����oG'C��h~��tL0h*�&���M	�˟�D�N=��=av��*���Z��jzox�;�x���C���e��;uK�L�� �LiJ�dd��9�Р7��)���a��\Y���.�P����_�UOEOX��͠��2�I|W�>��S���EX�S�5(����9�r�mjF�N��:���Ūer���pi�+���Ʋ��>{M�P�m���6��������bd���&=	�ݰI�����^%ae�n?6�@��V����୥��{���<Ǟ�*o>�f��i*,R�v<��Q���j�uN��\B����XOzWN?,����Sk$4j]���ɗ�v`�n1���=������(�78(2j�|�
�T�0�j3�@c��;��r\2��e��3H�vKy-����� j��I�����}��ʾ`VUʳ����v�3[R,��&������M����9���I�'�yЫ����4#���o%�;�5��MV\p����(�����uYK�q��U80h����Ź�diE�t<�*9(h�ۥ�r��d�i���F�v�&%��@qk�{D�aP.�R*���6�Nywf�
j��Yl�	�]��h�9�_)T^�x�y4VNY+�Ho�y�H�Ȓ���~�.��̡�����h��H�U(e/|ӣ�<�J�C݃=(�ܳ�3;�����l�:�W���#}~Bz�6ʈu�t7_�N��b`X����s��l�M�RUJ�X���(D*�*
�14I����|��u�6�	H���j�X�63fAl9aN���uc>���M��;�Ty�� ���?nn܁Z�;���Rn���G�(JP�NL41?�qĐ����aY�"&�����ո��`=R��o
`*��b7x4tR�����ԓ���Q
\�2b1~�[�%L�����dh����!ڴ�t���JC�#��w��+N�y���I�>� ˣ��\ ���,:Ic$�I���)֍�������gp�A]�4�7?�y",��:�j^3��[��w��TUj	��8���(�1�$�f'�y�6:)���H���_��y
x$��-��C�7ԧ�B��&e=9�e�P���X�0PO�Bw�ؾ3+�+��Z�mcR{����ť�1�XcrU�VZ�(*���j�<ȗ.�B/��o�Oj�$W3���)� .ye�d����g��U���t����[�~WՌM3�/�i{T�M�G�><1H2b!J�p�4��9�|*���ÕikCQ�7ߍa�#��g@V����v�9�9�ZKg*��+�a���w8�����E^ה/7����jt#O%M2�fh���WH��&V���,��p�yj΄Nk��r�ĺ�>
���cԧ�Ѩ(�����_�;.��5\�J��B�(�<�@�<W��2�����~&­Oƛ�)����V�M����ed��q����2f-�C<��L$���M�� :ڌ�쐿���Vg�$�;�rב�,	s��\dD2��rOF��O����A�{Ӭfw[�A����.�׊W:;�܎�+�^[�L���7�3m]|��!�ټKX�;3��x�����E{����*Tx���o��4� �*vw�1<�{�%a��4�E�(ox��3���OWCrM�
�