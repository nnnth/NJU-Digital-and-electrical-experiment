��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��>%����k�ջ*f�oE�<^M���2�j`(w4Μ�Gu>��C�Ֆdu�p�t�,cÉl���& �G1.�Lٲ��0vY!��|D��Z������{"�3ug�w����0�{~�p�����7��[�[dy5@�~�qQr�!�MvЕv�C�m2Wѵ?LK�?#��¦H5�o�_'�Y`c>3C�	@�K~��6���9��'�
�A�H���$giC;�'�C%�#%0P��_���l��Pw�)���� *�+�Ќ)B="�w	��}fFlZ��&���_�2��-t�h�6���s�꒮��	���SV����n��$,�zݛr��_�Q����I�Q��J�U�RX��!��_&�sN��+�(��g��27}&��]�p�o�}��ֆ~{�����:
E���J�����jZˋ�T�YQ�I����?�xma����n�`m�NLv{�@*�I�6�}f�ݭ?V0��5k�L�l3��nВ(۷�D�R����!{GY�F���ER���/��������ru@c�ӆ�/25���L`��� �L��M㗕[o*r�x;��
�P�,�4,����:�W�[�2�]����Id"�w=��Fኟip��T�q���čB_o���	R�S�D<r
&�#�w�(lݳ1�߫�Us"3��u�,�jŪ�>y�kN/N�(�C�f�O��/�~:J���%C���qw�D�5UfXI���E��:�y���$���I�>�~f��@��a"*s�đ�R�"#��z�����PMY�&�ra�2E���!Y����`vh�$k�sԿF�E2�T��}��̙H�4Y8�]2q{f̪o��;G�%v-}n|sk�Z�&�c,��H^r]k�x�]QR)�B��#��P�2
� �"V���Jd~��[s�26 B��;M����V���^�����ER�Jd3�j`h��$sz��n0��]V��ub�A�]��~��y����7�s�/�����,Ē�?[��j7F�(��0�Rt�j�MJ0�|����ez�⣹�H�U⺌�YOǺ@��N�l����6iO���#�����Z����R�?�Lύk���+]�����ַ֌$U�I��5�Һyn�4�,)��Gor.�KN2(%�b.0�Ro$�؁u'4� ���}��x	��+)� >N�={���5��LaVԧ���(3X�w�Z���!u�-�8�d��� �~���$ݪ�Ԙ<�O�iqK&�t�Pq�ԍl��
Wj&���+G&��j���n/�C��PL����C���>b*�� !e��=��qǬ����6��f7һr�F��t7$B6*�|%6��'d���-"���b4�P�к:��q���v��|�.+���gN%#p�4KK4*�e��}~�) �ե�UH�^���������NZi03v'o~ZY�كT��K����2�Fe�vs55u���Ә3ધ��O�'6
b>��K	�y-q��x�N^A��eQg����$@7�E.>E�'u�:�/�"	�w;)��g ő���T�ъc�3�Ve�UN��sZ�IU�Rm*�%��Yn	�9�\Z-�_\'=�u,�S�?z���������^�1һ�/�<-^*�T���[UU����7�v�mJ=�@9�x�F�SM����WTg��b��ؠk�Z��JO�T��)�Ap5�6�dn4���p����u���ᅹ�uPq��h��}v�S;�2�o�ށd� �B��	]H98��!�� �BM�;ӌ)S��O>l3ūj%��������Ҁ"�b��F|�}g݉[t����@���l���o�;�ZdBG��Tꎽ����(<�d�@5�����f�TQ���������\F5��PSpPE�f�/��c��N�@�{�ᘑ�crs�����x �fs#t�O�t*�'Z&��t�Nt�f����!��8D��?^�E���4����Dڰ��o0+�!J1\�$�[�o;��#�|�N��w�mg�kL����^[�K �Q�ҷ_d>�x��`�%���&��k��X��,��qr� A�Q2���wC��TQ5x�i�?�M���φkiO�%[�ER���?�,,���o�s&�{}9#��a�J�v	X[�]]�%Z���٣�	�jJ7��t��m:�2���-�l�_��E4B(4���'`*���b9*(�M�s;m��j���g
״)� }�|��g��4��#O0����l����^��c����91�g���&�L2W�������0�!7��[�e�;�t%������
�+C����/-�nA�U+�����y�w(��xb^�=�Z��Ƭ��"�*�KR15M�����sa���S��.B��l�)�O�f�Y�Hy����!x��P����:A�$Կ~A�tw�K�aH֤y��L�h@�w�yo����w-.��zJ-��1���׋�������g���×mR�=/}�!X�Y`>{n�p;�<�#(�fC����g��S`oY�����'�2�O�A��џ�$5�� d#���_�8�-7ʣ���M,�?3&��N9��(�LD�U�l����0��B�,�f>؃*�)�Ҙ�����UR�c$�H2B凰�R����_�ۤ�e�T)�J�
� ��ӛ�%6R���|����x7ўW�ou^�P|�ϼ��9�w���\�ӗ�o,�y�wє�U�:�+/6ؖ;R���A�������$����)���s�Ĺ�)L�8n�z��,e��w���r�F�Z`E��&�wS��}˂:����|��_���� ����k�2_D��:���bV���
u�O0֤�hmHX���L#q[tLK��T��k�.V���q�6�5_(KS,�	 �I��;I�K|I/=&Q֧�
q�^U5�)5�B�D�@�_T�`��gp��;�?��Ci�7ߴ�
��J��\}�W�Rκ0����T�L3���xu�-�1k��D-�[���0�G��!��wp+@�=s~퇿�l�������X��EIA,x�����}��T隥$��O�
wYZ:+�b�b�#�hM�p���cQ�.����2*9`��r��U(+�~WvM8Y|�� 3��m낷E�}� �/��uL�D��S���x�}#�z�@��5�ʆ^��l �cs�S:c]��oH�F�0P��8��X�ޛ��H�끖PA�_�����QV���3w�w�ۚ���y�:�&���X�g�nt��Lˆ\O�����v�)�P�U��	��ue�k��w�)O��?fO��PB3
�Ml�I��,��U�eo�%�O���Z�j��{��2�0��'����{8����cCVה�z7�³x���?6���\��w� �\�3y"�H��S��lv�A]R�0��X	�tU�[$����z���Uvzsݣ��0HV�(�U��ڎ�ԃ0����_;�uI���#����DB�_r�����𯂠�\�쌽!�K�1E�}���N|)i�o��m;W��LF��b�c_o�Dy2����"���$�9�� �ֺ�<�ÒZ�̷T":lٟ�0�m�5��?��o���1���[Һ�֊�F��NǮ��+To�������i���!H�l�~���ۄ�h�\��pCK&?��nve�f{���pz	���l}Ȋ�C�
&�!�@���A���|���=]d��pJ�Q�H3��hN<��ۦX^��?�J5^����m����5���%Mh���9BR��?�$j�2^��{q{�����Kz��T~���H[��L���<1�x�~r?���ɴm��,4�Y��UP}P����[�N�õ*~�d/GϡGtE?8�����1&�=����
њK����ʐlp�U�_�-8k���ؐ'�B�*�t�"��!G&�K��h��O���<�Xe8a�[�_%��2Ѐ��p�]d3FN7�9si���E���'���jT�-NR2�Juf��.�|W�M���Ʈ�)�ȱ����u�X�G�%�iu��;�"p��g���NT�-�g���6�\j �$=��u"F�X���:�*v���i�Edt*��H��H˽���#�uc���}�����3���d���\�BC]�������8���rEEҎƭ0���4,Fҕ1��H٫��J���7z0�6`O�
��]�����c�l~����bg��BR�jy�OY��\�]T�8�t�����4��4ۼ�e��|���k�-���Ij��d�%R:"gL�k"�:ΊEyp��
NDq����l�`q��3>���$)�������.�����^��G����kP.�I¯��#��iQl7a�2�7���X��AP��1S5z�;V�ҧ��<"A�;�N;�( ~���5�߳�:�yC�z�榚��48F	��Ej�@U)�\��#5TJg',�Bx��H�:���#���x�j:8�!��[�l;�n��7e��I���eZdF���`,�:�����x'wGL,\�����A��B����_U?d��(�(�d��#yQ�z�ݏ�΢Z�m���G�-������Em9�_�`��i�ǅ��.^#l�0���_��۝�Y�D#�'�sͅ��E�r�O<��\{�y"�0��y����<����K��0�ڟ� �J��J��-$��&��,�ct��23:s����5�0$b���|J� 垵�Q@�޹���� ĮL^-t��+y}*���5Y���<@Ǘ���#^
�t?>/얪g�51,�5H*�����i'M}��?G� �_�ao���?�)rߒ���a�Ų#�l���ӂD���׊r�fp9\kur��P����S*��˪�[��F1��0�Y���
�ԙ�->yE���1H��KJ8�[���j��*G(.��2-�,�a�)j+�"�@�[3�$ȧ���
>Ƿƛ�!ǈ�L
��m�g�c�	Ӏ?:XD�B,�Z�iIs%:�V�4��>��/�7fB�#���*�����P�����H�l��rD��3�W^� �i7�"���E�������M7#Q/�;a�0���nh#Fx������.s��c�Q}����  ���F���t�����~f�,L���i�	��l�\��'?yb‮%V5Sx�v̼���7k�m�4�~�<,�b��!�0���KXp􎽖�ê^���S���u���ӑ���5Z('CUi�J��H�)?�Ύm�f�J�9_7஭��;؋Z�:s ��!�Pb�&��0�M�éFoaN�O��^��qr�#&�N�N���@�.���W0>�'��}��+s��r�4Рb�u`@n+-��"Ny$�^�h������2�n�Ȍ��,�쨣�"kl��Em�:&u0��U55x�9����8�����PhÄѕ���H�s��\���9���w����<�˞�T2\�������G/��l; q�����}C��]?&T��")� igҘ,���Y)�j8A������~���j e9㈃��l7N6����1?����I��͔���+�﷧�K�*��T��{�.��pJ�Z`C�����Nc)x���OyP��ub,�ow1>�b`�Y?�<�N)��d�r��\H���+�ֹ�"%��(��HD'œ�$���2{Auw�'=����B���P') ���˓X��p�q�d���X���K0��޼���6����P�B���$y����.B[f� �95^�}�Z�!�-$�$��I� w���L0;P��Q��4؟
��₀��6��m�=n��g��!G#��\P�G��άvq��$|�Z�0q8J��W_c�&Q��� �������Y!�:��k�-=׋�N���B"���WF��#O����G�V�9��h�%��#=`pv�cgއ	���b��@oh��qv]a�6Ʋ�؂?��Ņ�'��8N&�m�Ms�5�O�Y>X��\xSt`��Z\�dG�~�n�J��f���z��fc�i� ��o����@���`�`K����s#PZ�s��P@/&�ğ��ka�5J��>��U������S2T��A.�����N��_���a��{x�U�
Q���@�h��@�~��Y�����p#t��Z댞Ӗ�$�X��Zx�Ƶ�8�A@��j!z{��j��2 �f[P?���3���t�ى��iA��&��Ͽ�`f�-�$-�ߗ�-�&�h3X�
�E�]�S#�fWu�`�R��H����A��z�%�8v�?[g(���B��[�F�*��0P����T��ዤ�&P�����M
�t\R*|�BQ�8*�X��M���&��M�T�J����]���8�<q� (A����餛�o�dD�ZS�����k<~����U��C�,ye ��%R)I�R 첮�Ԏ�� ]I�32_g�:�|��Z�^�59�C�qq��.��X):$N;�rF)C�$�Ѝ����͟��]�&Q��HlM�,�K����=�7����6ߑ�g������R��� zI�zB��M!]+Hk�_huyWh@$������,���b���FM�7��bl����o�/<�'$�Yn;ϋ�v8KI�܋G ���U�)꡴��\O1Q4t�.c�Ǔ|��r�oŸ񘈿����+����m!�z���} à�*�z���h*JS�0މ@&bu��A��>��,W*�ϱȑ
.藥�n*;��f� }��OԾ��b�C�g/2���.��}#�'Wi5Ĳ��&O|�5�Rz�ܙ�+�<A`6TQF�N��j3p��lv�_bT�^��i��g�hp���9��f�W�#�t��o+�=0�H�z,}�@�OfǙ�Z���ӓ��0�d�﵉i��`���6��U��m|b�G�.�?\����m	�톋��л��ֿ��a��I���K����.�PN���o���ތ���~�lT�����p��x�6���_�� �.��/ky��2����������2���R|��5~T���9�.�IUG])���- ]u������Z�֔A���]:����tJ_�#��5����>$sx�/��C�W�M�)�e��2��'�${����M2�ߟ���W~ ��C���s��a�Y��`��O�n�V��4����WK�I�G���
��La�P!
/�2z�vl�y81��a��l��eAj�-W�-V�ҳ�3�ڍC���3�v��� ���v�.�	�`�
����J��*�Zî�O0���ʁEmu��<z���Ѝ�I:�e�&~e�4u����B8XN�\;q�y5i=�P�!�f���{$�V�-C����[�QC�P'�J88_~8�%�k��$���ol\���VBd�c��5mϩ��?�&�{N(�oݫ��W�{�Cj�Xxƻܩ?����x:\%�d�S���g�Kk)�P��{8�^���J6���^E!3��3Tz�Q���A���6�R���=�
9!�	�����`�u��o���*��oe5�C�i+�F')(�Ｋ��e7�_w�<���F_ֹH<�R��N�TyR�X:ˏ/7�C���*ēK쯾0��R�AjI�m �g��Nh.�p|����I�z��;�ݾ4� y���/��L_�c�v���U�����,�t4��@�������7��
d��d`]����ԧ��c�D�hh�Ae�����)8l���L�(1�׬
�Z��Q"+���)o(ݹ�{r�<�N5��r��l��x7�wiB�ԫ�CK��y���=��@���b����1Z���n#p��4§$��T�TrP%F)A���5#R�g��O�VV�9�pe~���ΏJ�0)1+�<B���`�yӽ&��Q*5�+e��h9aӑ�"�{�(m(菩ը��2�E�H���ͫ��C����N�7�M�?��=�΅�FOa&�������O ���C�,v]�_��J�:א̉�>�h�D��T�.���i����9j�O~-n���.\G��=��顢l �M�hGuG�}���V�8�cNHs���~	)a��?FC�aV�T�8� �&i�9F�Q�+�#�����!�$:���܎�
�^�a�Xs��l����h=uAV7��2:y~0H�.-�X�:��<�^ R%
*���3ެ8Ub�7�ɞk37�D�oBSoi�ѓ7�Ďu��}���$���23�Մi$���I2���zL�����	?<�$�5ii;�Q��B��lVKt�N�mUeH��,��4�	���TRTl�7W,0��~����/U�@
�n��|TA*��A���4�������S��H�5q���d����syc��(d��� ��n�7�=��g��5�\
�� \H,�݌a��g��{�����fP��
ٶ��2O�A$��t)�幐J�R�8.��IygF�W��n3����������e�{wݕ�.�;�5&���X�߄zm���Yif�ܽ�����0 ౺�L�G���:��o�7�C�l���[�?��X�A�����<Y�`ն7�]w�u��B�"�6彿�vĤ+Okj%w}P°cn@{W������>�����j��	��2�Jdω��V;F.����d��t��5�7����	Jg3l�Q���b�r������w�ɀ��b'Tz��{��#�&�>���WC���u��u���͐I�<EӶ�_:��sG݀���Q�y *PL��P�<Ⱥw��-�tGڭ����r9&�!/\�?;�G-� ]'F����oNw�#�kki�譿��#Ջϱ8�b�f�I^(�#N���/�N�/����V��Y�#��Ŭ Zȅܣl<�T���� ��ۇ�ֆET^��1w������w��0Ο��h��~���8����Ϯ�3�[�/���=�Z�R!��_P��j�g��0�����˷W��/�-ge9����]V�n��\eF}KV��~���@����1�m ۞��Q��ւT��X�+�(�@1Ʉ{3�&�r�������ŧ9|�p6��~���� 0R`t��Fe�����74����%���wt���~\j�#�d<��@��s�q�C�"�8���t�v��ݳP��t��ƃ�hbh�Y��k+�(X�<��j���OI�2�TO5Ƥ�a���)[8k�%t	Y���d��!c�J64�)�q!��K��<Q�nԪ �u�+���OGq�?����do	\�E��/s`H�0���l/��Yk٥�K���7	�A��G�IuU��+-}��>��@Y�p���4D�Z��J����wl���ǫ:�B*�]����^)n�D�g<��R{���B�\�J22�������B��L��k}�<#d*�� p�2쎳R�t���~���E�?Z�tСI������(>O�{8n��Q	�8Z]ܴ��W)��2͉���{*��5�:���/��*@rB��V
�\V�o5�1��-��z�e���K	%Ww?ҕ�a�xƮM.�l*��7��&G�b�)>�f�0X|Оd�S�bj���s(q�+�N*b��|������k�Wx�= �8@����}����
��2�3�O�4r�m�S��AT5"��_�����^���"�;�Å���N-�S� %M
� ��ꃦ�];y(e�m�Ԛ�q������BL��5��x9q��9ƚ�+��oG%3�?W��z$3]
��T4���N�=��g��2B�S���O6^\�n��2'���*��;����_7�6����/g�B{[x:P���ȟ�@��Ĉ��8�F1���0���b�r'�΁j�Eq�\<�?����9�4ob��^P;�u�ˮ�#��+Ë.�y*`�;&ɷp���/Nyq���I��ivPP�R�\�@�X �����kp�@� ��Z��
�J��]}�{�b(`PqڽaUx:AX�\+x�G��Z��O7m���OY�
����;|�x�x�A�
<s���1�2w�e����ڽ�G�1 
��̴1󢣹�2�΅^�3���Q��������/���{3k��)���\9�Ӣ5Cg�Nk�N�L+�·��P�6R���s�Md~ty�9����Ò9���K�_�@Deme�XV��[m[�q��,���42{2D),x����3�$���4:�pG�S���
YS#��M&�8����n!lڂM�,qſ�p��Iԙ�2�3�.�4�˻��j{��G5���t���z"l�3����W���B	�؟�$6�sڇ�,�;�y�:I���,b�+�l;�V�A��ƴ�à�q����g|��Y�H��&m�
�g����K�
^) ��J+�Kra��gT�D��$�ѿ#�ܒF8�A�V	ɕ�ڛ_䜖�Ǜ�m�ۗٗ���z��<����ZŻ�F�;8F�?)���n�v�=��U� 8�j���A+�y�!n��l���js1q�;���{�o�9Ȥtxע�?�eU�@���}���-X+�7)`�u'{�S�=BK����	W� ,W�ō
� ��Q����)�=������2UeXK-�ɟG������U��X����ӈ�wf��7c�
;���vuq!�E����?��WZ[���(����k�)����u9 �x[��ݏ��)���ol/��}���6�)�||7���ܰ���l�����o�+U �V���h�>M��j
Gǜ��"�g� *s��/�+р��B)q_Y-�^��Ҷ/^� �ȭ�'��C6�Ĺ���d�P~��&:���B����b��P��}'�a̎�#;���]��+w:���e`��~�&�c�n2� �����LO�����5�����=�H�w���J�����%�~$����d*�c����@���LHZ�i�):��]�˩qmm���l����y��3\���Zw\�%��]"�G�"G��s�ñ<��-!�]�d��&�Ez�)fu���}�i�n��q����KŶ���VL��� b�Eg�M �6��_kx� T�9����ʥ��.�
���Q>0B��b4��J�������!��.q��-�j���d��ew��8�P��5nmq1�����*#��f�51���g�W�;6�c���>� F�\��f*9ok;�k҉55{β'��n�����z��,���5xl<j{8��lߢ/���w�<kܠ���bB��J鵴�ϋ�c@�D��c
]=��`v>��{�(A�,�Pa�"����ɰ��@�vg�eOs{�>��B�{6���\��@��9ۚ�YL+��dܑ���e��c����~�6P�pp>����7c�a�Bgx����@���N��������n��h�S#����U���p���T�Y���ac�I��b�i]b����%��E{��7C��P�LU�X�u���'Ub��Wd���k���U�$��u��Ea����|��#��^���ͭ���E��"1}��k�m��N�ұ�Bfmr�5a�e=,(�Rx�����5�N�+��٠q%�'D�����f����;�M��N8��L����E�u�����q���]�&{�]N�ăd-'z�n D����8�s.�pY��u�P�� ��۹>ϒ��tjB;�$E=~�7x�1O���xs�#q�ɐFp� *�fz�Ãe^�ӫ<kL �����>mp�Ĭ��X8�'v朇�g�N�	���0���"+rٗ#p���*�$\�h��TofDLj��6Ů`?�^���4�l��M���~�'|A��p�2k,|E��ة_E4)�o#$SB�� B����A �/�9�l��N��$�l�.2�M-��V9��(�o��DV��I<�`��8?k�r�^��a�;��G���QG:!*U�����:E"�r�lR8�KOדl3�&����3%�AX�Ǚ3��Mӓ�ׂ4C?�omX�e�n��yT�sR.2�5��ޏbU��d��{��/�:�^[��Cw��h����f��G���w)�"@ɣz�E |܀��go���LЏS�r���Fԧ@D�q;�P��>I�!c�Ǝ�-ߌh�����+��_�֢߻8��޸~	�l�dD�����Ā,�K�����v�Q�y�u��.�t�$[�S�[`�kd��q�lt@���]���1:2�a�� 
p[�=���z��YT
�[��%�z�r�}��?�����y�TإT_���i�����.�-�Z�i��T�W ���V%��<`p}�����J�΄���f�WfY�res��i���Qr�za�!�*��F��&����::�1��,��$<�U��Ncf�z�A���R��CM g?]	�:#�h5
-��~|�(Ph��i�`� �m�6��}6I5i}�s��8*�oq����n'��%oX���:&qg��'�p2�����5��%
��'G��n�#yȩ�V3�ȭ'�dB0�#�~;�3#b��U��>�1�H¾��]�R�N}��M�\[D��p�О|��@�5��M�r�o���ޮaf��UAL���N�v�J2[U���x6_,$4��K�d*M�$��ODl*�[]��.�D�s �)�D�Azd�B��8o�4��;��⋘�3!<6��s�#�H{�Z-�F� pr��G�ɾR� �b��nDF��߇\���ȃ2&Fm��Qo��70�]v�]R�}��pEέ��Lְy8�V�����Ӌ.�J�"�;��%��O�Ȇ5Dy1�����"H���p�S[_���,�p�D��w��#)�|V��զ�䮬ٌ���~}C���s>k���k�0���_ne����X���J3V4MC��d�jMs�K������q��[�z�
����tY4�*�hǘ
l������/���V/5-�'�c5���e�m9����T� ,�[�2eZ�\�!E��k5f�>B���_O�t ��B/��A�,�]�2T�ā�9-~q�Z �~�Ma{�85
l��������;8k�da�w���B����<��s��P`�bq��K�STM��������]��r��(,�h�	�eK�.����Y7դ��W���q�cl�1(y�@m���-TI%5�8��WǷ�'DJ������F��0�����t���w�5�ahv��ER���P~2]v���ʒG��]�GqEʔNxN�;��:��*���)�IK~���j�h�ۡ��cu�d�`�	\����'5՛*��и�����U]�}��N�?-ss��tVZ�H��wo��E��e���y�<��e�cH��?�����Z	�f�������=@�rC�~n�J��S6w4�����/C��
˟&�����@>"nĜҵ'��G��;�@�Z�@�Υ"�DLZ�{�١�%��^g���<��席-����'��EE���Id�2Ud5(�np��ƣ8�BC>��ꮮ'�Q� �0JI)ҏ�!JY�B��8}�6h���	��C�)x٤�Q�+]�:�7�I��"EXb��T�
�O��0�~��b�՘��ʢ0��$�Ȓç&�o5osԵܜ:_�+��=�yZ�y��� �٥C �Yu]�~�-��s��`�}Y��=!�&B'��|R�,��'��np4�GQ��M��WVZ�UN�c,��<���!�O��B
k+���;��7A2H%�֜�.RNױ��������ߕ��m0�1�@�ˏ�\��'ShKa�{�
��H�j�d�� ���1�<h�kΌ��DOQ,x���x�ŴJN�T[:pM;{,�|d���~rͣ-�bxq����C�����V�F��[�堿B�m�Ϧ���w�]���V�o��ݢ�72�$���Ig��=gJ�0^����%�K����Ŀ�� �^j���nY%ȏ��EmLľ�KE��os�R��q=X�*	~WB!�Y������E���y�
ZZР�W��b��#"|(ml@�@��I�@n�?LRf�|��hW����f� P�C�p���5b�'@kjˀߠ�*
S��<������a���<��ّǋ��6�`�5�]cN�
h,�Lww�I8M���!�|0��D.	�" C�j� ���?���=>w�bI�����H���"d'�6�L�]�I��]�rB�2dy�I�*mxdG
�IC��Ѽ�ޓ�>
d�I��[�L �Qh��,�	��Q��C���Kb�w�4��{�RB�4�%Xt��� P�M�1���'�/�Hh�T;�7�
���I����G)�Nm!˭K��X1ͲD#w��+�n�/(�+�T��1vO1��˞'@�t$�F[7����J���bk�
�����{�	��/���".��2d���x�?˗��k�_��g�㿰�b�0`���`B`}�i��_�m;�3sz:��}'!� ���0����z�7�d�����A]E?��dY�j�}�)�h����Ʃb�Z����ܒ��tQ{J[ܷ��Zoe��f��g�FY�^NM��؍����PPF��3)���]����R�%�s�ǋGe@Ǩ�w?&;�Ji6vj�7q��r����i.��1�n�h�r�Eb�����C��R�K*ۃ�g����T{��C�n"%D��K�[Vnǀ&��+QWֶ7���e�kRm�R	�yB�f8$��!����Z� p����O��nU�iO�	����!9ù��.�T�:]h�Y;,U�#�F$%�Y���9N���^�ߞ�l�aI��1?Yz׭�^2�n����	���B������B�,�枪���k�>�4��.��^ �ɸ~��=�������6�p#f11��/a}��9������br��l�w�7�{�&;4�,<y�~i74)%~qLJ�ýH��[<��ID}+�:`���M0bDB�k@���rd�qo{�e����#���&� W�|�0�������= ڹ���Po���t�U�N�!1>��Z˯2�h9��5�	�>��3i��;�BAJF��:9 π�X�18�C��\�ES0��zP���}4y_�=�]�y���Ys/AZ��x�r>��V��с�	�ʻ��6��3C������N&�0	�$�u�3Lv��6��Xk��־�l$�=xW�����!HQ�sB�y�$�]�Q'��S�N�GAӳ��o�U�]����g5ºn�I����n�ڑ6�?���!+���B������i��&�:T��_{)-��T;Q����O�9��-aB�j�/۵)�c`�I�a/�/���8D�8�ZS�����me V��;u���>���@��B혷@��^G��KaR!}Ve�O}�����S8Ĺ�J�A�nSm�eGk��ֽ�B�1'�P���S��dp����D�^�� ��6x�d�.�~@��d"������`:�8v`���e
�	8f���4��:��%�Q�߲���*��p֭I?4�1'B?t1^v��h:Ĳ|����UT��Ӯ��:�@��9�V6�	�X�w�~>����99���)��B-����X����X�5m��etפ�b���?h���3�?�o�;�Ӝ��p��=:�(�#S)\�Bv<�;�p{��ÛZ�����6P_��;ۻ�� ��hؙl��υ�������S��^=o���K�� ���II���v9A,��� �xD��S�x.���p['&
0��@l˘/m�V�ެeR$�%CmB<ƌ7B��9�\��*+K�.�**�]�X�Zs:��r9�]"�n�N5�CVpg~�Z�Yh�n@�������ۼZ3�{�fK��>,�Ta�eԃ��R��>.-�-��Ƨ(A"q�Zg�;�0Ұ1�Ep����f�l��.���V�58�7��'Y��b)&�4��?� ͏�-��b[4A�&��*���I(�zZ�����X*Tx�ԸOU���%�;j
�j�ei�/��	`X��X�l\�ܴ�ܸ��b)�/�u
����I���U=Z��I.�O�3Z|����D���ۜ��kPT����e�k��ĪL��So��alO*z�$k�m��h��J���%�o�x��ز�c$���PϽfˋs��ЋTT�¶M���A��R��_����#�$~����V.>]	�N�1�����h�[he����Ca����[fG�?~�@_{��\�C\��6��S$Θ��'�Õ�z��1/�&�vd���w�m���f@��T�y-Ǜ��[+���VW�3��,e�&;l�%�С~�d�W��XL�����aK��:�:J��O��o�2V�i�~^�\xf��Th@_�����27T�/fr%cn����U�$4^�@�+QU!�7� ���ß�g�5�D���'4��vth paU��Εа��S��۩�*�%�3W+6�
ᎃ��өkU���͹��J�n��@>z�_�v٩��;�5�,��Ek^e�E�}��^�;I�t!o�A�p��%��5u"� U��|8Ld�G���3�S���a��v�$�����=- ]�BMK8�pr��jxza��������5�Ʊ#K�������(,3�wݭ�W;�9�PA��xs�˔tc�|�{�"��j^�>�_A�`��Oe�S�-5fD��7G�A+��N�J���p�1|�����/�Z��My#��3���<;kr�l�� �zM:P�C�സ����� �kRq,���o9�� �MN呂��ܽ`�'1t��*�/c���x�ϼt�ְD\F�E���$�Ӓ���ļ�Ϥ��z������^0j�a���뉲���`�c_�%�������������ߦ�Aͭ��H6����%t�[r��w�|��{�.�t #QP<j�n��Y�!��zF�5����>?�ʡ�lc���h���L񷽘A@[��,$D��<��JAz�S�>��H�P�����̛'�k;*�1��Y��G��oֆ�j^8�S�M��A�lo��L�[�c�~*��,m땽�[��:�h$B�4x�����}�L"3Bo	&�@U\;Y�8�B�"U�Q!�UK�&o&لa3�^��X�΄DU'rD�W����b��/*B� o��'����e�&٭:-V�/Q�?��Htۑ��j����q%3�'���'7�3� &mk�_��R"y�M�b��Vu=��p�kg�^�&�Wv{�5¬D��lIZ�0��c��N�|��ۼ /�j;@|&�1����RhVzL��H
�)i�d���j�{��6�~���x�� &y�,�e����:��xu�/���%���Lg��kb����zb�]��N�t"���?e4Ev���� �p�^�$F��	z�̟�O�SЯIK<���r��*����S��%��ކ77�4�9��󻞏L�+����7ϗ�>�#O��	�I��I*y	B�Ӻ�`����F�5��1����O��mp�rF���5mܱ��L��}�����P�]6&)2����������b���l,	0F����h��,-��N
W0����)�� ��Ѿ��_�?>)��5�9�:\"9}�:��'�SƧ�-L/�&�0Z��E���gn0{��x!Cw.;l�P_Vc���V7�;�VH�<.	���0[Š�Mww������
��IP�*�	>^P�Ł�`���s����i87�l~�������0ö���W���~-��t@@=��lf�+]f2��2{��CU D�&�" �g�V��a<�2P6��{�e�,)��G�-PQ�z�Ә& ���R@
&��&,��]=*��͌奟�����m9𖝄�\�� jc�=B� >H��/.��S\��ɣ�Xw��{b��sx�oo9�1��:7j�:-H���aD�ǵ@�WE@(Jb�!cS,��(Z�3��Nי W"Կ=r!S�� ��Xj�ո���l�`��ڲi�t�8Z�-�H3Y�p���K��.v�������¹��̖�b�G���y�g�D/�����W?��\b�P~�Lے!FB�
̵:����]���ah��=ȪWu��m:y��B�U�8�^W2��Va�6W�K��Q��{��G	|�0��V.�Ӹ՞R5��q���{�,���(��o݃��dRE4׎�\dU�z�3Ň�%��0��bQ�vZ���c����D9e~�l ��cn"�CF�Ӄ�F����X��'U�����~`��?�Q�%S�y�87��<��uI=�h���5�5=�t�텱�\�E�� �9&r�KX�2�b����V����������k��pV�M��e�@�>W�t�سR�-5|k	�����;�N�J�x�����1��"��n*���M��4M��6��r�Y�Jn�L�6� �|��p��2\�c:���B
�D��!
�c;���<:��"�m��\���5�؏����7�6�z���򘈠���T��|�C�5�k� ����%0ƽ�Gt-���lm#�C4bE��#�����*u�&ī�D"B��(��ܡ&r(�M8�T\�abJ������/d��)L?K��8:},�~��<>V��JWx���/�.vi�h�v�_�2�g`�8ٵ�9ݳ�e�� ��QXS�����0�� �eH����3Ι�V������	�(*�i�o�e�0�Ly0�
G�����wI�T��v�7!+X�7{Q��<	o��ւ��8]�[����T2����~ ����Zߖ�b������)����OϏV�ї"�����}��}�T�d���h�O�Z�h��jE�������io,�v���4i�\��C�����G/�QV`��$(t%p���߅F]��#3'n
u8�	���o��e����ۗ�rƤ�����nk`����W���f�%�kkM�G,P��fT�����4Z]ˢ�'}�gR3�"��L�
������W�������ia�𩡊d0����:v���\��;���W.tH�/A���E��g�Mmr���M�N*�5�3� �>oK�	���f�!�O=t�k��n�Yq#��}W�dU��=Hz���@���a���k��7+�[֏�ER�U|�/�͘EiT�ˁ��F��(�P�������_�9��*����cw�g�񱺓w��R^T�+p���r�Q�$5�vG��e���S����lD����R0����v��Dq�yt��w^�ޛ���+�$�����{�O}m�z���(�ʂ���Hq�k�v�XV�]'C�g���^��{(�HkN�<��3��J�m�0��'�X�p��I�̂9k���ɾ��V�����ـ��V�"�i���- u��q*��Aa�Wi���J�P�KlC���<q)^S]���=-O_9���ƻQc���b�M`�p�MS����X��f6��P��h,L \�MO�816! ��x͖ؓ|6�>b���������\��Ӣ�'�i�:<��B7��zr��h�rj�B�j��u[pRF��*�4:Zip���v�iRm��=�O�*�u�^��e��
��Q�l�ߖm���b�i�sxu��
ݩ��]�gs������Tdb�W�����!�!��6Y���c���T�,�Jh^'�h�p�=)|���,�A���|�~�8GLV��ZN6��D��d�W��<(p66B�~�ßh��2�	Π(��I`ۇ�y�ɋ(s�s��p����$�(��,�_i֏SLk�US��_�}�:!��2��5���j��dh]QQ9= ���61ѿs=�Z��	�m����&�ӄ-u��S5��:�o)è��J*.N�-�5)�P�l�d��ۨ���=	J��~2�*a��S���lؖ��M9�&bc5H�������U�e�k�������"u��9�Q�e̠�bx�ԯ�S�z���3�nF�6�d[��a�i��A����(-���#���A��S~��!��Ff�Y3x�j̽/[����	
�/U3&~�yWuoјv�A�������y"�J;l�����Bx����7��e_h�~�lI��M��1����&�A�� �d�x�^l��������y�}v���G�/�w%�ˋ<2����Qp׼Z��t�5c8i��Qt��k��Q�������?�/��<L�+д�p���)i��e6Q�Bx&�3h"�gC"�د̍?��}GR��3�ϼIYCnc�.M�.U4�1Sc^��AR8��O��!8L����W�W�"��cQ�:��&b�Q�7*�o�a6���=���S�-��r��PXd��3����8?P-�+���j}��,�����6�jh�Yt_��tU�#r���K��@,������S�OXK�[`�ӈW6%��}��8u��sCDʫV��<v����x ��!�AKi�e���Q��.+�U�q>V�tS�"Q�J��$G�s�L��q=o���m"���qi6؅pk�q������]���a�!�?:4g����$#CJT�i���G��V|�Ü�f�I��#U�`�_��7�Z��`�1ɅO���]8�sF�"�E���p�$��ti��W�=�dH��ׄTSm��UΤ4�����]�B��Lm�����M�H���LV�ԳB�w�[A�޳+���>9^_�#�L�{��{�8��[��q̴Ԅ�"���C<M���lS�?�������'z�RIu����VǩK�e
���q�!hXb���
n�0��%|&/�V:��n�4(��a.�Ê����)�O��Ӷك�' ���y� �o�}&U{���w��u��AQ8Oc�:k����`oCt�ӫ����j��� %c��8�ˊH��(pLֶq\yU��2�<��ϭ��((�c�x�r�D��"���?³]���������ԢeR@T���9��	����VʃC]�	Z���;n���y���K�� �( i��,v>ԭ��#���]p���y��HA]���톲'�'Z$sn���,��:����Ξ�՟��i��f�Q@l	�y�|�sv�I��wK��:��k^�OSY�p6&5J��V�~�C����3�jO�P�e��o?(���22��CM�����h���S��
����ӵ�k�;;��M�7�������{�H�0���^�oE.����"��6Xu�$�h/��q+���u������C[ud'����'�):�\M���$����,XH�ȶ�(����.�/���8v�J.�j��U�
�L�z��,�m?�>�SO�]u�e���
�$OƱi�?D�B��I��g6�_h�Ç�ȩ3��Q��lCc~���{e�ܤ�ҁQ�:~�m���%�	Y�鱁mxs6#[n!3"c���\���腕�L���pfF�'O�dpz]]���^WQ�,;�Sr���Ko�	T&.KVe�n�0�>�<15�N�U�'���H"i������p�|Kw߄)#z�)} B<�=���x�e\5���wzn�=�oCo,�9]����|/��`+HH��"����k'��Zc��Gv����?PM�hv1s%�?/3m�s�\>O��5GSj�ܵĈ=@
�g7*Yd~>�#������q1{�U�4�e���/s�B�KW��u]~�̈́�h8�`TmNB8�,;��{���n�u��_d�q�1��,��=q9�3�1�Ѭ���B#]>Wc�W)��X6��0�� �ɱ����~��7$�"9Qu]�N؉��$�$�f�Z�bAm���p�.�`���Hl>�H4<�
�����VgN
���ĵ�{�P��R���8��w'��g�H��35��).D������S%]pF7ߋ�gp[��=����w\��/h@����=�_�݇:�l��Y2���IG��PKG��j���i� ����E|��f��J��)��	�D�"U�Ֆ` �tc�g�L�J`3><��U���%��z����4���/�N ��!�,�L�S�/���՗��)�.�LY�����(���\��;��k�B��b�C�\����@p����ǎ(�T!D	5wN����Ct��17��ǅ1�|����!`{�$�' �pz&HL&�MI��t���;n��:du�a����#3	'�ڶ }�)ATۙ}���da�����"�W��	����:�wsxy� �,�Ѳ�4��Bi�k�Ct�Ah���KRg��[� �&5MhHK X9�NFa�Ŵa��I�3Hmm������a�����³1���`0����D	�'��)��YTlZ��	u��7�w��