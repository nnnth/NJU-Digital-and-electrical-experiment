��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�E3�hoA�zFҿT�,��/Jۭ���Ab����4y?�;�GU}R=����ā�`I���u̭��-�ߒ^Z��^Ha`��4�M���(ilU�+��!i�]�đg^g��}�T���gZ��5V��DekJ/�x�z��/��c#��Y�@�J͐:���}���Dc���#���wcɴz:�lέ���A'�2���rmoN�`j�X]t.�$�Pe�MCҐ�Z���;���A9ά�8�{Cj؈�g\�d�=��?��A]l�~k�����������_	\a:�sCg�;I+C�o��Un(�I��WU��J�_��7��}F7�O�>D7j����oG�M�k��:��N��U�R�/���H�
"�s6��U��1��4�ׅ�>pt�8��Ѿ�ZR���0���}N�V���v�}�lx��!>r��A�-����?��5yci��6b1�M��40�*���:��&�����.	Lf�D�D�x�~��!�J$cm6�b-gMofX)�f�z�'�U�1Z=�[�<v5L]lc�ؕ��h���>�yC�m�e�]{d�����h��c4;D�<�W�f�鵉�b�B���"^�y]�Gz�.�>����R������<�4�Xբ��
��*i�D��I��y5m�4���mՓ�f��=m���tJE�%�������*#�m̴�y�u�,��_���lݑ�F_]�0[>P|���I�v|�+�H��F`gE�˱J �7�2�x�*�w/�6I�B�f/hp��
�O�
�� ֺm�5�x�~��84&ɞ�@[�}���j�`��Q�D�8�r�-'^�"Zl>ToW\�)xI�}��A��rݠ�wA5m8Z��#����{�>��~h��bǕ��YJ��)����g	z�v@���pBch�-0�et���R�t�Hʑ��8u%0c`P:X�@��Mg�d��'��j��b�9����/���_�,��2���)a�$��5;�"<6�,����w�T87g%������zPG8Lnog>��L����>QN�h�>Mjý��@�}�žz�v^bA"�t@W} L������[�Ք׍w@����^��I٢��Ƅ�qZ�N��I��\�Y�;T�'��;���Р�52��-���i���D�K"���$H-�X�)�%����5��i"���3#�~�����G���&��i��S|o���D�����$7]����+`��[�������e77�4dԎh���Q� j�ب�H�e��άROe���<�"٨2G����ϼ;؅=}=�{�Y�s،�����g��N����}�l�*u�t�
�?aK��g�sFsSF�����\����BJ3���˪g��i���G�"~����]bC�Qδ001� �a:��a�����hD�e��5�ћ ʛ4o��a�l�_�f�գ��h�C��o?Y��[���<fMe#Y2i�3d�ᏇuQJ�M[kB ?N-���'�!��C<�i��L �<̫ `�����D��jc����WDPX�,�-'��+),C!��i����ս{��E�� ��NH�k�W]ag<�!n��zF�n#�*�q�'��L����]���hq�$�Ew� ڧ���(0�y��+i��c�.EF�i�X�O�2���/��!��澜��P�K|��,m��Iu,�!$���-�:*�,�K2�����\WO�I�8ap?�Dkݤ'�0��{\P�Pݶ���.c�@���,�eL�Gc�1�G��r��\$@�+e�Wz��
�,l�SS<mHU��|�9b�}l��<�2[Ӌ��fH�r
�x�2���<w�.���j�.9�=�����X��0`�U����7�܉�\.Z�C�YQf�3#�y��{e���5TA3����,�攮�8�"�h<���>2by&�~X�V}�F�x>�%pSJ�9�
���	� #���7Z����\�cPjfJ숊ȓ�+j��,;�::˽��g�a��ygKj�TyM�M�����������ӈy�� H ۳8^�"�Z�mW�����9�J��X���|��c�!�p /�A*T������ 飝G��V �ľŌ�Z"�]�|���4u}Td�.��e֥���K�v� B��iM���Lh�n훑��BD#8��`0ń���Y�eNZ|�,?r<[R����vDKQ5��7����}�Z?��8�VC��Fw-��?����L��U���rZ#d����Ǐ�&��)$-�4ue��q��7ʹ���_m�-\��	��p���c��&�� ����~\V'���/HŪ��HD��)CQ�F)��FX��#�2���ץ�*,��q�n��ʮ���T<U�r���E��ϕVcmn��B�h�Y��t�d�G.���&����fIgq�6<�h�_���ܻ��k�+��}6����XS��%��vZ���7�	��QE����E�UM�Y<{���%[P����cPz�����2�r|g�o�d�#���������"��N+UfB/����5ȧ<-.�iY��#<ķ85�w�'�m2�? ĄdE�@{u
��Է�Pա<O�`�s��t��pz���`�D	Z�qQ�e�r?!��ί��3��:����^�2�Ft�{���C;'���)���ǌr�@�G6����vd��z6Ԗ��ml���?*�����1��V.1ա�׃,*�W�t�ӝ��HEn@��t_�"�v�]�5�{�+��¢��+*��S�\T��,��W��*�vp��9��vc�ꯅ:�◪����Ҳ��dˀ��fi㘍Z6�9�����'���Q���6)��X���y��$�炉Cӡ[]��6����˛ Ѵ�<ߦ�)�^�Y���'�<�KJP��&"sF���6?X����ʈ�	1�����>;�;!I'M�H/��!�Ff���A[�AH�Ș�X*��@H���(EƱGA�0M��"u.�'Y'�#����e�����U^��,u��:j�`�J9��M�<�8���ז��w��`dg:�M���	�MɥY@P�@�:�f3X��V� �C�e�"�ֵ��G\sDj3pӌH�'>���m�N!<X,��1����G熪�o�g^h>eBE�w�H���w���/�F �?�+Q�2��(�9X���}v�̂X�iĢ>���)��(��;��B��|o�p�r�Å%JL�H��,�	�\�����Hi��SF6É�0"i��d�S�45���:�����dc�YK��#���|_)�l��[�G�ڼ�c�����<��D]w=�Z�G�t�'�Y�p_vq@HpEm��饬)�EWG�B����
Kթ^M��:��.��L������{�ζGj�Ti������^�x n|(��E�C�)��Gp�)O�0�c�q�
�0�s>�.�1��U�=� �
Jz�"d�M�����O�*^��t���$S�54�����b�[�&�;�P��I-vO�����=����h�1�j`�02r����x��9ł\�6ڠ��wr�S����ǟf���T&Wr�{F1���ܟ����:��)g�Ӊ��|�$f��0XB�q�F~B�ً��P��R�ـ�%��^]�0h�`h5j{�q��k���KB�鸠�w��̳�����6S|�a���lI���W�Ճ�/5��X�TW6��u�e;롪���,���'b��.�e�J<������u��6������Zi��c�<����+�����\�E\S���Ðy.�Y;l؅�?[m�^���w� "�r�u��
��uߋ���7D6o���9�l}��!�V�1vF?����6B�ï3���D�9'�Ķ�B�x�D����W�\��:G6y<�nP��x������`^�i=�����Ķ �(�$�s/OBDN��K#X�5{u}��;!���t*wE꠲&��K�"��/vs����$�v�ӼIU&�8Hc϶S�}yv?U�1N�3�Ey��ve��0��l����f=�@�*�t5(���u�8ǿȥ��Se;�ˍ2��ڴ�Š2%�og�^�����W���r���z��>�2t����n���]�}F:���f�C7\b���֖���\wMN��&:�J�D==vvŉ�1��n>0�n�ɱy�K%���3gWND��(o�ծ����_�;g%��m�U�`dU��*볦J�O�=�GfΣ�6N(v)E�)w}�L�\�h�ܧ�7�|D,��_�[m��\f@�1c&j�r�`�uH9;�t����8��<Ba���Q�#��"�*��9��X��ܪ��d���vH�o��ؿ� )z�;P�{|���4ؚ
cfΨ�%�td)���y���^{6 S�l�|��T���8z�#�����c����_��F{�� >8PfifR��(��故vpqލ��0Gi���y~����{�ܚ�WH��,�F�?���®�L�������y�7&۷�zGy�g��(��T촶�e�}my0�ʡ�D�o@,�}���8���KUW�=p�jYV/�&�74�b��(8q`��+�Jz_�G��л���oEr��P�$�K�G��_Ŀ�)D�Ofh>��ُ'E."~����
��^�{��l;eE_l]L����x+lRc�"g��h2�AĞ���߷?�����7�AdN����x��
����UXAPń<���j�^"[�&ۿ&G� ԾӞٓ���d@>6e�FeXt�xr�����˥�����]������h�j����u@�^�O&L1"�'ڲ�֗͢�}���"^��ota��� �ȸm{/6�!���=`M\Ϲ�6𩞥�㐷�p�<��8^ف)zqv�e۵؞.��V���;���d���e�! vI��,f�v�i9{���c����,�_?�Kr�+'�z��ÿٸ�l̖�s�7.�D�Sǲ�&��P@�5Ԥ�lr!��ygmq.�X�FVi�nz�iE��H4�:�|0Q6)�h���}��ߒ����`�u��DDU�������f�yp��&��dї�MK6<� ��M�Ds4����ߔ�S-��`�`z�K�{��X�����v>O�]��:̰	��8�%��Ό��p��lz�������T��c��p@G×�I�h9Y,e:]x�f��0�h���7�K�b�\�@ʇ.�`t�}���C���Q9�S�����$�ܼ�A���!T�W�rOt$/��L�g��x}�3W�R��̙�zy�.���+���I�{��'ܶ�K����ΚAL	ޡ�b���}��GX�>��E%�;�-�Ų8Y��6p{I�u���q���R;Ƒ�P�Q��_��U3mMkj<$+[1����Ȗ	���sk�%������:�S��U���(�|/�{�T�a�]��B<�����2����ێ�#�[3�!�o&t�K<�t�x�������;��b]��֠����#���	�c�'7��e��5b�I6	�KZ�1�bd���o��e�KZz�$��4ZK��2Y�R�$�bI6.���\�@���0{W{x���i[�)dӤ��\n���`<(�kӘ@�4��	Ǘ�_��z�r&������,���F�'�ܳ�J��܉h�gC૔��>��5Dn��#����v��`���1y68�F�jJ.x��i[Ѓ�����<v<FU����H��	���7EXd���O�l�o��P>����k6] �Sm��E2��GmW�1"67�)�,�K��>FϧUi#�p�ݤg!el���F/>N��@�}�!��c&ةq�B=�}���}|��F�>���R�$�( �kdD;�!`*�׿7M��T���~�hЙzⰐ��M�J���X]1�~�b,���!E|�%��m�Sp��>���;�۪q�)�U~��*<���r2��b�Q�[�4��}�|^�󲤡�A$��6�������٠Ȅ~z�L�X���y�N\�f4��ڈ�?���4Z'����o��-��_2�j�����$�_�^��it0#q�����^�y�T��p����Qw�L�r�}U�S���ӌ �tz��t�>�f���p���g�o��5M@�(MsL{z�/��2޸E`�O�t6�� *�!.����D3lq��1��O�
h�p6h>d<��b�W�#� n�������T�4�(�8�y�kc�Hf�&��mt��ܞ'���1�8�˝e����m:$+�ʙ�&��{�7�+�Ö^��h&ɓA��³���?�' ��ފ�����>��MM�U9i�@[$FEK6^��[�kN�5��Z�W�Ӆ���G����$d����Y����eSހ��kq�i�4�Vf;B��`�B{��'+k+6b@���?�[�Cf.��*D�8+��A^4ks�̎!����}�s��څ��VHHf�g�ty���M#b$�P]ti���f�\F�J��	�U��&��T��T- ̠Q�Z�%E��l����3J#���/8�˂�z{�l��{���HRҿ�$4�aUsQO�=.��X�,͐-ؼ'N�d���d��G^�7-}�ɡP�fA�41�������/�g��ٞʂ�XXvx�0<�ůz��y����{���f�����G��|9�H����]�K꽙�n<��:�Cw�\�� [�0��'���]t��b�G,�J���3�<�jKB�y�o!T8G���!)ONH�Ha>#V�g ��J�w�5"��� �L}��0��t�Knuc�[i"���#y�LH�N� �Z)�RA����F��ڜ��t����}��1�\�H���LO� ����b4�!fε�^(+�1Հ���^�YYF���G�x��9!���yC6�gx#�����f킫��fUb,����8��	������قă2�b������z�z:CS��a�0tZ�W-�X�]�����7���$;q�[���cH�KP����@�~b���6�<J�O��a�l�P��	.�ۗD�k���T�!gg@�ն��w|��,%i���ċ��&�Ӥ�rf��+3�[A���hn������i�^�~#�4ݚ����L�|번�zg#=P �b@���������3 >&\ע��5��Os|���y���	1w�z��	ԋl����r���Q[�kg�ɿ���)�DJzD�$KE/វfjd�<z���ﵾ����^�xɖ�؁g���,Iu������� �/�����#��P��êU�=�K.c�ۈ�EշSr|j����U4��������U��������Q�˚a`]�'/����/]Hr'�$�gH� �S.;>�ӗբ���g���vPqM��\[[F��)�-ۙ�WS�\���1䎂���ɗ��n{���6{v���Yy��r|��ݏ=̋�Ķ���jB����iǸ�I�^&���][_�*����̙�$	\ a@m}�ǿ�tM�m�I�0՜,;���:z�ρ��o"}��<+��!�^ū1t73B���Nf�B��m����\�-�.{�՜��|`��1�T%���gc���K�GH�v��h�3K-d�K,Kc��O��2m��:!����Ht�`5���RH�lG��'%agKYpn�ɃsP"�0o¡��)[ә��4R�!�9�dP��u���wm[)%`Q�s�z
4����r �bŔ�l���r��C�����Mhq|�!ɱ��L�@1]Bӱ�,Y؏3b[@��ҥ`39��\��U7��
=L)IZ���rC�Ds
�v�8t
ǒ�F�8�KE��5��6� �_
EV��nCN����B�k�u`���{e>���q�Z!���s�����.o3ұ�#�HR�[�It�v�`��93��)�	w�f��'�������O;��r5<��+�x2K��^�ó�[Ic#����+�����+��!#���m-cp۾��5ZA��z}�ؼm��9y��Rw��������M}=���٠������}o�7�WM8��Kѩ����C�I���*��/��;�%�"4i'�l�j:�.��\���x����]�!�l4?���s�nUl�L@��[�uooC�C�a�هlnO���}�O���Oh�icm=��&޵lk���]#��H�}����&������Q�c���$�>��瘂��+�Td�uX�����OJ� 3��o5�Ъ֞b��_���!M���z����F�����q�@gi�g�3�
y�JY��e�ǹ�I�o
7��c��Y��1��g/cX��E�4���JQ�Zo"+GR�c<U3�1�q��j/���~T:�O�B�u�uĂ�6����wT�����
���ş"�6�t�u�b��Ғ�����*��DS��4��A̅ 3\�����V]?M c4�蜵�BɄ_����px]�¹�D�Fu���n�I{ޛ0��rf`'�F��#��hοHt*#;��p]���A�7���|���R��z��#�ڸ�.��P�G���k�g#�|���o��h��c{���0)~�䘭�� ѽ�1����nh"-���>$�Tk�SRJ��ᝡ��8X{����F��>�73�7�n�,#|R��\C���oc�<ρ[n�B���J�K/()���F�qoT���YM� �Xm�\�	z1gu��j���XG���G��	^9�*��Ct:��7��#-� PԐ��3@>�ήČv5GrK4���Q�j<�.tג���8�#�FF8���
���p%a��Ko�~VI�ex�;�y<O�U�
d�����c&��W8_��~���;`Ί7��}-h|UU
��O�%��Q.�-)�U��=e�}D�L�\�^+z�Π���P]�ޛ�q��0k&�/��J����ݹ��Qj������n��1K��o�S���I�W�q{>1�Uƪ���	Ǿ����!x"����w�k�'�|������P��+��}�BAձ�K$�:
*����0�k�Vt��d�y��ߓǗP��'�T�S�r����kc�T����w�Ќ�#�t4���0��sS�퐈L?f��	��Z2��ذ��]��ΓLT���A��f�5��r��%�Of�h�)�ܰ lɒ�)2&�5�fxx�t�6!�w9�e������g�LD��;=���h�ۧ���X���?؟��si�;z���~�)f����s��c}��a[�'�wu^{���mJV���pܜy��i�ְ|�v)� .�͹���
#�h��^�o��(O-غ�>��r���3X�p�4�-j�BB���܏H���������]:�5'y)��9�賧u�����_�bR�3=���p�UO�W�Z�M%`E#[Q���ϰ���8���nQ�A^(^s0�갿J���j�)+DC�d�ڧ��+�e�yB[c���ěbl>J�r�Q��(R�����S��d����u�}m+����-�ȷ�4�K��4\���ky��or{EHN>���z��f����K��(�!�����E�����+D�ZpO	`�S�����ﴡ�훿}�w������>���Q��oh��=m��%��w�0pS]	b�w?J�aU�4���Dkv)�z��2�RZ� m=߃���=|�)E���t�\|E����x!(�i��q�~��F
�S�N�x6ޙ�-���
W�CŖbrG]-ec oQkR�m�[�ј�1����L��O�{�%�+|���q�m���v-e�G?Ǝ��* ��-a�¥�������A3��H�:u�HEL�T�sԒ��6f'4)t��00U��&]Jё��ɗ���,�X�J��	>���^��.ú�Ð�˥G�WN�ָ�p.F����:.��l`��
��"���m�BY�tD%�,l������v���0�Y�u�PA�t� ��0d��ZT���������~T����M�ke:�Č@R��H�G=�qY�$�S��&kP]��97�"'鸵A�A��W��� $�|g�d����m{��+��w_7��]i5:Y���*���ei��<}�'ي(�N|M�15�'kƯC����A��v�+�,#��K������on��Vjڒ��Rt؉�$�p��:WJ�u]�@� Z~������R�SF#�I�a��C�#��o����[�7�X$�072�0�V�k|��k��'�d�#�˽�x!%STA�� �t|5�0M�q�W��jV�.�x^N���	��B:�#Q��~���"�8�m���X�rz@���V��0)�o���jkxh���QQӺ���Vk7�҇�Qܛ�������n$��a9�o�����dYÔO�e��^/@��Y^]�Us��l��m�o*�5��]عAp�� �.����[���/�}��U�j��U>�֟�aG�eb�� ɕ��c݃9�����h ����zZ�l���$���#��b���֬���B�f B0���Q�־��&`�3�݅��yǉ��u����$6��fր��ޱ���=�Hs(��j����e~Ĭ��2�F��#ϞG13t�?�N�qaH)��zN��/�+Z2�t0��
:@c�0Vu�c���D��g�	�8��Mm�Vu���YJNm�n?r;��V�i��jR���c������~��6�ςn+r�i�bK�&�_*0>��Ǐ�!:� �����
�מ9%-�U<!�8�I\MFW�m��2*YD�)}$��3t�͞���C+:��X��1���&�������]P�v�Вr��uӫJ�\�z+�<3F�֐�NuF��"��-�O�ldvv
��e����>6�edGV&��l��K��vV� x�uq ��Ӫ���ZY��'�M=U�_�8Fl����Z���Ґ]B�u�$� Y����5��I	��΍���
. ��S��x@sr&�����9��^��A�������3p$�M���l*�?M��{�̮���������9vj���&#�/WZ��.�a�5:!P�E��#*"h%�	c��S�*���T�t��Q����&?�\��w��y��4������XB��>��A��q����.�1����](r�4_*m�{��9��lՙ'�+$$��;��#+ �0ú��=�.>���~�/��s�C��Q-�Fݏ=���e�?��W_��;��p�}7�Lt�K`�6���#7���-����i�,�a��cq )<��ur�N��'v|�",�Ҁ0���7.&܆*N􉆞��D��!�t9�K�^��f�h,w�sNZR��j�Ϯ{v�̡��`��&`�!��p�)L;��`)=;��5��aIԌ����X\�~g��.˛�� R�,D�lzu��0Z��"[�kyEo��g���ǣ�m� �h�˲�����<~��GQ�P��HcH��Z!��^�Efi}s�X�sBt����츱~��%�U�J��������Th��>G��ho*v�x����ԉ�
fE�1� �&�������D�!j���-d�vt�Gޏ�	��]R�Gv���r����M��{����g3�JKwX"�3KG6h�)��-�PBY-Î�ma�9�Fw$f|�=l��W�	xJQ����2ܓ�h	���E��d.�MnD�����^t
�GJn�>h�@׬ۼ,�iXAb��	��o����],�k�~�亜<��_6�$ȭA��#�<��w@�o͹pG�XZ��lax1�A����-^��[*�|�%=�PS��:m�g�Ew�b���������\��	B*��4@��>����B�]��
PWDH`�<[ûo�:��V�X}�����E�dE��<%3�$�����}���?��ɻpDq|��;��OU�g�3��8����':Vh���*z�,]8�kEk����y�J�Ձ�"�n�K��v�^�ң�ٚ����;���L�ٕ2� ;9֝V2��H��/���S����I�������}o�Q�ܮ�#K�'��w���X9	ibb���f�GY��&�~;X��<Rд�|O�و�w�+]H&�#ӻ���?�K����"$�w)Jʘވ�I��=��D�����d7�>�;�]��
�$�g1�l�t"]ܐM����6��~��J�9�0 5��?��V:� [ �ә/�_�w��~���3w ��b� �0�:����nρ�z�"��
*�l�Vm{)��v���#9�P�����wA#��5�R�8��6Hql���8ͫV��
��8e��p���5��k��Τ�~��n��w����������5;x4&�*JZ`��c��r0A�!!A
-��E�g�?���p��)m��LkZ��7
�I"<�D��B�P����/x�����ϊ�2I��B�:˷A��
9����(��hs0d��環�~c= � `z�&w�G`ü;��O�fC����o�������jM�bG��r[P޽��gbpE�K�����9�*��,Xu5Bg,]�d̰���ܡ:�[��==O�>�W�n;�9z輑�
�|b<s�2�uEn�mV]Qgڒ���t�4n�� qO�Qv��M�o�R����D��iy��#����ˑ%��?����r��7熈�����ں���C/�I����
�ʆ}�I�YW�t�At���a�OT�j�V.�y_�l6Z9�'ӗ>��ևC&(�ݪ�l�3nP�� �V��O:��{x�✻�Z����O�O#�e#�Y�VJ���<�TR�U�D}J%�Q�b|��8l�hZ��x�&�yf���c�]qʄ��Z� f��|���T\��6���!��Zٺ��R$������$:�)>����Ė�)��^e2YRq6B`?�j�1�,bY���N�� ���!�A㾱,Y
Kk������#�����*����a&.`z�qc��dh��?��r�vc.�� ל��ۛE��N�ctW`�0���W#�2�3 �[ժ
4��  �FE@73��-ˊL?�E[�����k�3~��o�DSt���`�{'1�x��������&R9��vF{��#l��5�b��L�ۭy#�A�5F�dc��]�����t�7����@T�(�p�L6���&M	��Q-%���Yg��ǩf`ih��3B���4�������{���n�a~9�Ȋ�׉-�|U[K�H�;[UJ��~����̱�_q�Nr-��l���[�����z�_UZ�Rĸ��f���ΑȠ9�
���z%xJ�����Ӱ�LL]�����:!�������Uҍ�;f��L`�Rk�F���N,"��3��D�Ln�:�N��3�������B��D��UDD�^�#S�׎p�P��C8\u�JQ���_z��ཱུ�BS�����a�d`�!Բ���k���ncW���T�2�6`/C���q>��L;:���Ul�6�V���.}��g�@󺾾0|p$.E�qNS��m43�)KQ�Ҿwp�I���w������v�0����b�'^ ����u89@,�3�h��ZaDR�D�3Lyh�l>���d�����iT�8�����Ɩ���?���ՍNPC���x��@�_us�qG��u{�F�7,":_����c���5owO���W:1��g��
�ys޾Tn#z_J�drN��9���U��D��υ�9�E�F\О��[�a5ft�e'ަ�d$"�T��A�Zw?y~t>\���7Tݿ���k���:|tU��;u�bÂ�����I4n"�O��E3�O�|]h�-�|R��gr�Ev���Ʌj��	��9���k�$�]DI�+VpC���Oc
B�ut�i�	[JN�O	�Xq��)�+�T�	���d۪,J�O_��Aq��6u����S�e��8q�h�f�n7>��I'��h��� ��""p�(o��U�&��H� �J���g���[ٗ�ur_���3�(�-��D�.$�&L�����v���)v��_��.hz�������s�*����~��q�N�9��L������0k\���k]Jd�ܯ�+�o�ޒ�Ȧ�Y@!�٨�
Qa�A㪚Vs4�����)d�daX���+NP��>o� t�{[��=�ӛ��c��T�x�Z�;��ZwW5����n/�m��Ԙ����+�Se��T��f1�\��ܫ"�;K//"+��(E?�u8��`����NS 9�$1�d�EZ�݆u6�:��[����Ȇ�!�KsE�Lj/�y+L:����#�`��T�+%�˲�Gt���V"R�/s�ݘ�y�� =���5$>kfՁ6���[�n$PF�F��hb�"��L���>��}Fe�����*�Y�ɛ�Cc�����SVpe�*ɅFr�#�n�0��� �9|����[��Pl���$���6�]ڋu��戟�-�KB7YV�g��28�1p�1AF�N�6�_/J폴�&"�d�"kp�[mKn�(�JY�=�6����-��Ϯ�f����a�Lm��j�  F�Np���1���ܛf]����íw�Ӣ:.)HA�~�⠐	~����|�ȴ�\Хhʬ^@B��@�at2�`��6�zm��4v�>kr�SbB��On����ٺ��yQ5d�O�>�8��e����ƶ�%�;"KY[�^�8�u>h�N��z���Ԫ|��4��d�B��8�m6J���O���� ih̻�V��N���O��"t}�5��"Хt|b���
�#~�ʠW���PJ�h�f�����Z��ړ�O���җx�wK��F��m�`�V.�./l��P>���-=� ���"H �K�Z�_#���	{Sg��K	��a��o��4ԤS�*/p��S��^�m,4���ޮ<s��i��w:6q�d���9�'n������oѝV�V+lN7�\k{&}#e��i:fL�jO������Y��2ϝ��;�Z�����:ՆJ�/�=��#F��h#����&�*r�ֵ�r��b��B[��99d��駕��?��V����'1)
4����[y��3 ��_�f��LTU���-�2�v�*���Qr��K ݇��
���k��1�"�7�����2��Q'�H�S7Ao�o��:�'P�AU�`%k X�6����(���?�z7�e88����=I�;�p˷z�N^v�lZ��Kb��TVot���l#0��Nv�0FΟn��FFl���!+�;��A> ��8_x���?g�|ʭ]}Wj����썚f�~��+�6��î�5���S���%�D�!ϳn)�D������O7j��&� ��x.��&�v����D�����}?IW��K[B�T�q��.xV�͖ j�c�z"����P��0;,��²�I0��W�+0�8�[��ҿ[[�\^EP&;��������#�FLfݯ_�Ɛ���_��I�H��h_�Ψ��W�	�er}Y/�DC�Xܞ:h�q��i��^aC�#���q�F�*�ܴJ��@����>>����k�;G)��<�ٶ7�"b�@m.K�Ϭ���	���ED༜JZ���Uq�}hqd�x� �g	��D�^�-�� T�}�KTܞ�sJca�ǷUbO8:	���U:��Dׇ�5j����+��}S�}�hh����\���Zq^Ω �\SU!G�;�tl\���(�^P��o{��?J<�`Oq��z����ta^~��c
[�^<��Fu?-{�U�[��������j�%�Ys��������{1`�s,`(4��\�Hq�AAu�D��aǟx�Ýׁ��8W��'n�Y1���c0����6䉏J��L�nO�"Yk������Q�i |�Zx�h���A��C)�=�4�ߋ�"8{��ϦO�I��%������1�'_��Q_��Ln��yo��7��{M���>h��U@�h��T"sT1�w���o��	��	Z��hg�B��i0���6M�X��Z,�c�@��sP��X!��x����kG�<;���Ԑ=@g��r��\��
�i���+w��ˆ��Gؤm(1v�CcM��T�L�����X�4T�K*����N�� ��Eq��`i��,⡜�V5����$��}�x�K�ݴ�B�=��Xu��i���4ڀ�t�+�4<�Ч#�]�la��Һs�]��� fs u�-ʌ�,�+��λ?Fa��J�/.qY��e�����u�g�P�}A�j�+
��k�����)�n��IkNĖaV�z�_V��UBNv��ge�n/+�_f%a����ԧ��L�[����%� -��F^/+��[~J�E���f&�!O�!�0Z5k8R����Ɋ׫�������Y�S�:_trϨX� �9�,ᄕԡ'�Q�% ��urUU8�mA찹r�6�3�RF�^]f5��f�9Bw����rJV.{2=�R�����߱-l�pD�<Ij�V�o) .����2-H��2��F6�Q��ҏ�S~8|�ⰼ�m�rׯ0:QIl�!��I�V����ۼ�����-����VcC�?�~y������iى4�X�I>�;�`#��E����\	>��&�֎�Q��ŮqwGb�e��]����|ڛ �<`ڛwHӿ��Au���Y�����d/�F��E]9���b�p 闕��|#*�����θ<|����Q�ɫ2,��ߨG���6�'#$aࡀ@��X����y��Za"[!aS�5!6��qˑ�G<���9II���h��R�t��f�-��WF��AҘ��AA8���'�F�WN��ԓ&�@j�K�+l��ֻf���6+-��A&J��@)݄�N�2@7��S�ecޮLP���Q�\k-y9xS2�dy�D�䎺ޑ��h��+��i��p�1F85w�
A��"`i�G^|k]�=���d&UA�/���� �T�c�ߒ@$鑪����ג���+�4�c[}^�҉mS�&��g�}�b��Ɨ9�e؅�+�?#H�F���6��H��8�1-����\����#]g�u�� M�ٖ֝� q�B�u���36�}������R�I#�;.>�k��Y_P��"��f��Q�~_���v�W$7���=����ޏ O`�:k����x	]�N#����LB�|��us��֎ $�6*-�3��Qt�.8��o����� �"H����i6�K����M�B$��e.�4�|�@���Kً˲DD�=r���m�q�{F�I�T%5�=��=[<�q��+	_r�zn��Xn������1_�_tȻ�F��"И�I��986����.�z?'�Q�L�_<˟
1���嶧�rh��0�JY�ʎ�Y�^��oϒ
VfU��[X5v_��l�ol��5T_�9?����,�+d��
u��I�%��2�m�X�-���;��+`�;���h�R]���^��<��i�!T�sW�td�a☀U%D ��X[;�$���yƴp'���Rv��|<��b�,Lu��md\�DS$K����ݕl���y�?.�;k�U����*%�)�E?>*9�)��P7�C-�YRcu�x6��?�i7�紾q��=t@�}u�K!��c;�V+v���(k|����U~���O�"��Ze�����-��ɐ��_Št؏/�|�p��n��Ȁ�х�7)o7�q��{f� X��ikd�������1��o֏h^Z�6C%eZ2��ڭ�_}���\�<�l�sf��]�^E�T�a*U*����Kr�إLfĝ�^���CJ3��T���c�5�3�� ������/��Yqo�k�<�t}��@�չq�qƪZA��YY��7VA�՗t���tʴ	9b�kj(fb�S>�)���`��!�rY���BpM/�yWPq�NXh�CH�/D�`p�aH�YFLN����������2u/�}� ��<�}�{�^��'�t=�/-�l�I _�d�N�
�!O������V���;xI
-2B����z���i��~���*1�,��aj�O��W/�y����	fؚ�2�[�|_�g@�P0�rI��{!�W�?U�L�p�����a���ޝ��Q�	������N`�S�R-�P�d��qv�)]��V�j����?���}	WTRA���t����_i�\�\M(���]��� ֊4[����Js��t���o�'�1�Ҳ�:�]p��;G��Y���z_�!���>Rs��~�;~*�5��1*�V]N������f���@OjtHQ7@����kj���Z���ܤ��� ^�d��՘�ls�ʐ�d)��h�Lj���8�r^f�q��"1L�>��'��I�o�4e��zf�>2�k}?ivg��/t��t?pp�}��r��z]�s��.���Y�d|�¡7�Y}b
����Q�$�RϑKGC?��Q�ءe˱�5�:h�6ņ\��3f� afuO}+���0b���q=�d��|c���BƊ�*
�������8F4���)�CF����dŪ˸���q�X�t�[c������'j�
��Rɘ�m{�
�����b��������0��iN}9A���^�7��F�<�.X��7=���ݦ�Ǒ�ｄ7c4���eme}�(�ۦ�
���QvgD��*��:�sY����{ź�̈́%=�����U�Q��N�x�`�eU�GL.����ٕ�P�R�"5��>ɩ+�������������\昚<u��P5�M"�9�0�D�adx����p��H�tQ]A��T�üFΜ&�Fs�B,�p$��L���4��"�����V��Z,�d�p��8b!Hz'�s��b���_B�5!��Al�t�:�w �j�|�;������7-�����2<��4Ko52O���fH����r(J��T���<��5#�>��=qNT������f���i)��	ǉq&������t�[�ܯn�%��L��v.�%G��f�bO��ώ����m�!���[��Apd�Kn֪��m�
?B.s�Ţ��Gu���&�M���-����8<l����t�=pU�a_qv�jH�h�ũ8�Aب,is-@�> L ���ɯjjl�874_��@�բrG��F��xX�s���Zo����7�ji?X+5�،K�JI޺�c9�'�t�����T|�-����+X}����3��!��0J%%����ƪ�ߧ�$�_�?R��ղ؛ׅ_�(ƻ3i[��oh�CӪK�u��wS2(� LnD�?N���Y�K��#�������. ��eU��asQ|�b��<"��U���6�G�rJ���r�#f����xs�1��<0Pֻ�<	!�Rh��`�b�t�W���n!D�i��ѥ0ga#���K�� �����&+N��zN���i�D;�C�;|����V�Uc��kH�8��V����X!�7���S<UAI<���L[q��Q��`�0O^�G�^"�ӷ��7��v����9*���V���!
��spV̍���R*�om��z��T�Դ��i��h�M�;ت��~�����Y��||x|,��n�ɬ�!�rk�.��V|Q�ߞ��H�B����h�j~f+\�M�~�1���-����\��߂�����S�V�,�d��D��fq��>��#��� I����������1�f��_�RxGl�e�^�#�R���g��͗[�x��ا���.`�50��쀍 ����j��K��I�Ʒ#�<���+^`Ը���<�i p��܋���s��z�[� ���'i���=p��f�%F]u��^�}ѯt!�*I�;��xJ䩦. 4N�L�:�)����9��hܱ�q-CV���jB{�Y@n�*�des!9���Jvـ�W�d/��8�
_`���sљ>B�9~������N�ev���}Gʮ�?|-�Y������QL�Q%���>j����_`�wx4�Զ����>}�^PZ;��`$w���۽LZ��QV���G&`��9�[���Jί�!�1`���{컫�ǜ9��X_<�Qf][G��*������q�%�*��3�SH+�,��,�3�5pML;�������t0�э�mP6ҁ:U�����@S�U�2`���̐C�Z[�k�U�3T�c.)���Ɨ|�"/-51�v��hp���j�e�F�Q�ծ�_��u�x3�<l����WTQ�/ym
*2�U�t����QԳݽ�{OZnu��XJfno���bh���e����Sg��n�{v�Wx�2�ʤbν�N�;�@]-W�_-?,�@r-|�/ y�R^.�B��H;���䤉�_��D-�	��@�@�+�IQW��r��a<#�>���/�
����@䁿�#��_��JK�E�p^(D#}Jx}�[O��E؀�1����׈�䭍�"j��^�C�n�_����������ճ�F
'��	�1�Q��dJl��u}�n6�A�ֈd�V=̳�{5�,Ŋ�)q���r&�PTepi	/	Y��
�g���Kn[L8>u�ps�b�.F�d�MɃ4�����9�V�j�����3�9�"��ແ�~`Q$�]qb�������p�� Ŗn�N�Rz���?B��ҡ�hϙ�-p+vL:���{G�+�0���$�Ҽ�
_҈.Dԉ�O�k����@O*���Nl�9�r��w�7��
}JF8n�_���޿�4G�[��3�oO)[�������
S�m$�.�iF�xo1�	���%�Z�|qWx�c��5d��3WӔ�&(�
�>v�|�~^/��U<.���/>��d�h���~�����Oτ!�qs� �N�#!�Rƫ�U���i	�;�F��0j�������N��'�~��`�N+?��c�ą�����z(3�����uM��{^���a�]Z�gt���e�N��c�<����$]'�SK�ǬϺ_끑C�Ͻ?{���w���MU��n���W((��o_)�P�3����Ԧ�*�3����=]�s���!��B%5a�hA)��e>s��/1Kw�4�7��SN���ۄ����B|]���<'P�D&6t2ؔvm�V���m)��%��2�!���e�Q�;�e���wj�wM}�.xsL���2� o���K���SZ�a?iԵ��z�F�a4|"�zSt���q��@+�3ZL_*_�� �.`A�d���:�z2��:6Jj�%�����c�����>F�Щn."�����"�������sp�%Zİn�W��2�!�)�˕U1<&܋�������RE�'zaZ,�P'��z�W��C�!qpdl^:��KZ?�(�l��-;y�����h�w�� @˥q��+ G�R��u��VI���,#��$JZ�qB�7y~�z���t�{�lE�8m.������%�� �F]�ɣ��l��Kw�̖e��dG�:QIS�V��i��;���k�Vo���HX�)Ln��a���b��F~��A�"$"O+�;'��1��yd��Uyo��!n��g4�#1���GGr�a�'7�^�w�6�<w�2�k�sy�T�̙v��^CO!]A���f�.	�~,�h�T#P+���<�>�I��H@/��j[��ȍF$�r����zIvN�!�^xSG'%K�%>p�@z�l
� h�HA~�����Q��1d0��T���ot�fF4�c�P�~P����\庶�X	�]�9k�nꈠ�Dr�G1,W��b�d��?@`ּ�����/�^>��ru�	��?�ߧ�N����2VП�!��M����X��ou"ܣ����[�(�~]ƨƭC�)*�m�F��C�9�S3�H�p:"_����/�Ϗ%O���s���D9���4�]OO�@fM�[9\@��ƥK�\� �=�9���sd�Y��ſ�@��^��Yp�`�)�Nr�b"�b'�M㾛� �+��?�� �����
���2s���S��d�&i�-�ȋ�d�+YP�tw���H�w'B�Q
�m�n!Q��MY��f�)�h��-��le�P�<������V/�� b����Y��8xыo+������ًws�-Tv�1�ݜj�.�W����k�~�܄E��J��a�eYj����� ȷ���)	q��С�mks;PsM��Fv>�+�}U�:�I&�2u���6l������V�x����+�<D
�8œvPl��:�J�nqr�����I��Sݭ��o‰�b�s�P�ȷ`��dc����rp�ۭ�8�6k��F����<��������	!���ĹM�7:ѕ�O��.�VB��1S���I１�st��sc[�����X�D_�BD�ɫE#Sx�UMyP��XB{��}�����$-N�)zO���E���"���	<Ƒ�X�.���}S̥�4�6X�:��j+����{�C��kC���K�ŗ��y-�� K����(��2�A!��,P�DiK�r��������ub�0mb�Qoέ�X�V#�]D�w)-�����NS!�(�D��4�$�\���|��.��D����S�)���䪈IP�K>�l6p��!�;�n�Y���}ɑs���[R��
X��J/^�*.sE��پ������ؐ/I6;��v�r��'K�� �b�B��^�K>X�M�Vֵ,F|/�Ul}ġ�^�k~A}����Dׄ�"y%�m����w�l ������Yǫ��F��A��3�|�T�Ѧ���ϵTc_d,L�{�8^ʻ�3�;;~}J��#�<G���XDb�m��i!T�b`���=)5�-`Ϋ�qڞ�2��֥ð�%�!%�	�� ��>�Ơ�: =��s2l��`�1�t�ی����B��O6	e�>�Tv���~j�A��|�T�3IJVF�G� �,���l:\�� _h��e��R�s��s2�/��R:bH��CO>���a����c+b�#�hO��ݖx�Q�6���`�C�z �cn�M��_��B"���\u���wE<4ጣ!T�oFb�-�����
	��3��E��O4Q�;����;}��2 ��`;���I���"��Ep�-*��qV�^n���Wǜ`���̿;���f=���m 񙌽�=
��u �x�c�)P5f�ֲ�ɟ��OmBZe��=S}�w�Z��3�P��E캿�L��^���0Ǿ`K=ç�/�.�pu�J�v���8|/d����)#�F�f�	�f��o�V�$�#$�<�>	�_�K��c��nQ�o�E���Ղ��يs=�SX9I�6�=�Ù�3�-^�%���t�[�Č_{�[���KZ�"�A�����@�w��?�|!m�Y
��ˍ���&N�An�zA�!�W2_��VfRi�֒�k̍~b�ey	|p�����ԭc7g������U�]n�����2٢Cٗt��7>K�X2�¤�
�DG�sPK!u��\L	�꼷��k@�γ::���ˈ�>SxV��ay��c�ϟ���~#jl��������@����C�>h�&�)��¾j,�� Bڏ�d	�q�W�`�3�}�����蒠���!��ҟj%4�#�R_>B��jz<� �U]��U"��_ĪtV�ڌ���es�u6X�zy+NP�ƩbT
<����~��Q�a����� m6I��F�|��.q���r��R��l�X^"�aM�V����iIUI�ݍUh����~�`�HץͰ�<h���	g�ڼ]� +�G+�iY�`H,.9VH!�*p
J��U,��e�1���*��H�4�']"!�FA��[+���4*�`�7Nu�}�/�Eb�ʣ
��n8�0&���Q��!��Bx�V�/�|��n� ���
\�Vql|��_�Xn���D��~2�����ь�F$�v7����@�ulv��$�ߘ�D����u()�qB���?#���:Q���আF,��\�p����eu�\&~ı�g�sV\�91�d��,}����]�?s"��#��b=��%���`�V���f
�u3+�Y��zؕ�t����F�&;�D��O�0�i��Lx�g����ؚW��(.�e]�PB������/;�"�/��'��.]?HΝ���O\p���%]���iȁ�OdY�m�R#��}I�p���c��u��M���D>,k�^�u.�6��	ؼ>K�� �g��M�\���t�8�mr�e)t�".�bQ�z���e�b*t=.<�dθeJt�`�W�C`���APٍ,����Ӷl㧞��3q������>3Ԭ�iܹl~rP�'"Z�<�Sp9� �O 뱏ztYn�E�ry�w6Q���|OMѢ"��oH��o�e�#���i�~Ɲ&|�da$M�W��Mâp�0c��m���<=ޒ�v����.̊�0{:�4�6�$��Tt�~0'l�Җ�����[��Tm((5�O+qEU4K�F:�ΊD�}�kO�&�n-�?8�������Sl�YIspkT��J��t6m~Z�3�3Ҝ���l�[Yi/�|�<s1)�Z"e�{���[S�ܛ�;���>��V���v^5�)Uq�և��饽�̅00�I'T{\ ��HX�o�1N��1������pT��W�F��%J�)�\j���x/b܂�(� �r܋��6F����x��$n�[���7ZŦe��P1VSII�խ7A�s4�F�{Z�u_��.ڀ X���[@���e�xx�7[�����ٓ��۟�E �Bp<$מn�E7)���w]?�<R{��*��e�,|bv!�i=t��I��D����4}߻�\�k����|�g&g�8a�Z�S�,9���_�aN�)m�82�z���/e��#Bv�m1]��uf�^k� ���H|�A��A�Tr���EFx�lyU�_>Msʤ����k�^�e�D���qfcv�Y¥�Є���."Yyt�
�\�<6�ja��v�<^{���i�?:���W����)x��\0�^�:�l&4)����M:���]ϳ7�
8���t���ߔ�Ξy�.�8xf�����˼�W*����5��˶ܪ�W�z�������&�ͻ�	rQ>�g9�����cb|�"I�e��Szb�md��/��JAQ�����D����ʯ�A������ď�w���$���b絕e\�ox]H�7�LQ:� ���K
/����"m��Ҙ��6	vZ�t�m*t�Cv�㭖o65��û���U��C��_6��u�2o��	;��\�`��4�>�h��p׆"J��\����%:���C�D�@!Sjni�9T�.��W�����������u4	(T<�-p<��!�,�x�������fp;b}��T�6�����v	�(�V�n�<G4�X�8����^K���j����[qKK�5F'Rj|�o8�I�"�Pw���%�G�>'-1�e���J�r��UX���A)���Y�n�UR�����T,3��q�[zE��r2y�è�;�+i���1bZ`��g�c3�n�Ї��M���?gި��uqg��w@��_��F|(�O5�?U�0�6)J����<v��J܌�uT�(A�x~��nyI�+ y��<X�ؔ<�6:B�۪���_8����9���<�<��)$ѝX�����V���
3����t�j�t����$�0�1���ڇ#�m��l����Z��9g�>�+ر2�E!�LŮ�R�a�0](�At���ﵢ���r��9ݬf|':;H`/e*��0��,�@����Ȱv�)Xd��--�Iߝ�@=_ ���6��a`a/�5���<��`BD���)z%�1���V�ѧY�.��a]�)h`Dp(���0��L�97���*�R��]����z����c�M-	)�p����,~�Q�
���]��Lc�/�3�<��]ڨ�����QL��@�8��H$���Wy��-�����}"j�E��&%�0�p��Ե���@@���-��/?��_Lb(���?��,K�U��Y2F��?�Ss5���.�9L	���YЬ�y9B#���u:gd�xu/t��B���q�|��!6T�z,�$�5ى��Ja;¨|c��>]�~lz�IM䫲�o��&$�5��2��oW��x`���kF[X?���\Ҥ2C�s�\�ډ�=O����*&�$T��{ޔ+�J����W�v!��O�k2��N�Zf�	���v�l�S�!c�#�$��n�W�c����RhP����!��5,��X�2��M,`ߌ���ݦ��fA���Y��2�E��C�[R���&�R�dR��˓ĊC9��<~�9�Ւ�i���U�+��C
Ԑ�Q�x6�b�"i<R��\�tMr�~?�V��~����ʥ|a�5�e�ys{��� �C���G�a�u�%V�9�wC8�#�N$OД]�	L!q�W��ߧ�~��4eǗ��N���YQa$�]�U\,�'��@ �4W]Ͷ�� ?�ᢥ�K�GnH�Ű7�d3��=d'��������OW��V�%wq����ak�vL��AB_�J��Jh �=��2鷽F�އ�f�;�xrHj9
��v�	َ��*9��Q�a��мg�U1�&��|c&I]�ByߢP9���8̘�Te�� Z�ʜf�0��w��
�,'���ɪ��e��U��W�3z@���Se��m�Y�e���Ƹ�m�V,]*�C�c�~��w�x�p��� �UWd���Z�!�JͲL���5��˚��]u���vǑ��̬���Ӷ �j����.��)=�*"a��2-�6�����k��*��n=$��xQ�䅾Ͷ�/�!�;�����W�HP���>"�D��#�1
�	6�.~���gz�O%�k�����W݈elFG���p*J�,%�e��ӍK	�rn�Y�7z�'S���-���#.4�n����x YJ��y�u�����k˛��B�c� �"�SՆy�gb���m�T����2���ql���'��/HY��?40����r+w�y�-}|���48H��m`ՄdԐ� EG鵉� ��D���u��֕�R�ܮ����9�jŴMl)s�-�h:�0���hr."��3��r}[�x4ca륅@QO���6�B��&�@3������޽���rX��1�B��~I�(�"����sڮYC�*Klv[1��}�z��T[�'d�Oh+�/\���%ƲC���5+aHi9�I��z;�f������a��_�y�1LvH6Am��SW��j��vֆ+79�y1���e��!���%.ڨ䠕�	�#A�����j}F߄�՞@�����'i Y�L$���e����- @���s/��y0��&�����a3����59�Yf����/��&/˝��᳋Iz�B��F5�`o�=���K����6�p���1�"�e4&k�d��r1����.<o@��;���kk������
4�%MUz0��%5��PƐz��?��E5LRo��� �ՠ�Q2�TO�^=!0�����M��l��Ю׷�#k¸c��ז�T����5�)ϗ�[�wp�	�?&������8/�R�&!џyg,��qO�7>5�9Y1��?���M�R5�r��������ّ�4��e)�\쌳�.+����J)8���O>Ȼ�{֗�3�י�/�o"f���z����a��	;�-��as9�N:ޱK��X:����5&"�+�R����Y������w�������&��F�g�(xbO��ūNU��b*������V�����+�{�so0&��T�6W'���E��������8s��?��?�V�P��l��8D������
�HZ%;��G�tg\j��k��k�f@��iM5(d�+Ef(��I�X[7�U�x�ķ$�6C��Cgq���v��J	�=C�6^�W|����ȼ^�[���s�1�m=1z�nn�	��6�V�� ���#�p�W(�������ה3��p�EY�E�B�&`	eL1R��Fvѓ��jd-�1BvJ�_uW]����`Zs��@������fB�<sTD�H�=�p~�g��* ���7���I��ы+BQ"96��Rx��(e���ܐ��$sx&� �Q�x6�gvV�7�3�\� p�h�B�9��tiQ8�ŉ�{N��=�5�Ag�%X����~p:�g����*��D�i���E�"����e�1�dą%�5]���;mV�aE��tF$m�to�&�~:8>�jq�K��:�1����Z;G��	��j��ҢmI&1��&$�<A�KZc�5\<�j�!H�ˌo%�Z���榪�N��c-�ۿ���dI�n�P7��>C�5��iǟ���%xH%��/t��� ��.7n���İ��C
�r�Y�,��w�*��e��g���<� ����fL'ƶą����tj·yn͊uc�4DJnT�s2�?������t]c�&���sK���V���Ρ���Ag�UE{���Ւ,��RZ��W\��P�96�FV��-��[�����rQ�o��ȁF�&����Ȳr#����7FJ�����E��f]�?'g)�@��"'Ў�쉜�q/�8:�V��wI}�_��d��@[�+�[?k�o@ȀJ��%��HfE3�$�[4�u#u39�}_d�������*r��h��X5�Ҧ�]�d�?��c����cl�U��Sr;��n%_�W�����c-o�lB�3�ZNwj%$6PX!�W�Z����p��^�tvk��M��eG{J�}�}�Z9�&^#b���w�nW��������Ϝe�e/�]F�C'�ߒl��⨓kdZ�R�X)>��
�T�dm'�ہ�7�E�݋���$�B�}��,�'Zۉ���Hbxh ��;����IV\�%���'r��+Ǽ2g�2���	*{!W�Q���\�8�h$-�����%!I�G�r�d�93T�sZ��pG�K/�9�A*��1��ő�9`_��Xn�w��,��BL���`&)�}�_Si�HWqq�0/��2���t������a���cZ�w�oG��E��O��P��ב�S�?n�_��5Pv_��W��[tXr��$Tw�~`���X4�(JSm��O���9��ݨ��Z<��%�N|*�d��gԣ����g�#66�d���3���ir�|`,��h�:DB&um4r�Kú�u�F�"i��],l�N줞�4/:����܉g���O��J��u�����"&xs��	�����zwG/��5�"�;*�O�'��D�̬8A��.��N�+���eۤ�$��������[)�!Z)�9�3p��o)�^�#lq���e�ֹ%���>���0�ȉ�䍸�s+JP;��q���"B2C���$��!�Oլ�T/�A<�bR��AsqB�Ta��4FA	��J�^�c�]]�{���1����!�kP�y�-7Â����N�q����Tž��4�əݳe�����D�h��wA���FO��s]B��(��&1Y�j�g��b��\9�aP����ځ�	5��]�{��V5��՛H �,;���p$)�I�_����s�R�jJ��^s��$� ��N'���؛�L>�`��N��ר�5i��鱕���j�K$���$��"7����u��[ī�����`��@�Lİ�]������?�_�C���Rǟ(	���3�k�(/<����ڲ�Rӹi�C�� �n2z�����p`�8	
��7[�s_BL�Mt�iG$�V�Ǹ̀C ��@T�=�y���+yl1�unQ��G����
׹ώ��.����1a���^1��9����rуp�!�ݢ"	�/���w��WPPm�"?�f������Rz��J�����'�X}x,v0��㮒�{j��V�?�_&��ޔ�Jayf�G�!8�?v���3:�!:���^,�d�,����t�(^�^�V�j[J����j[�Xq�Oy��)��ך~�C�S?[.N�u������nuԴ�� 8J�7dz�Vz!���v�x��@��	�y ͱy(E�d!�;`z���R]���փ��J�D���>�B�&`�<�<�>�'Q�%H٣��5����� ��v@�(5"����ppJ}��YB޺q�0ͼ�U_���4}_���ೊiE�iYv�]�`�ǲ�s�zvF+��u�a������#������f�t�{?�p�ӊ��."��2�dYw�S�h�m葶R;��Bٯ�f�4|2��{��&p��MX�Ap��$�k��p<.�N����J�N���<��^���Po�S�6�$9�}��E��28��k�2{ECMB5s.v!���>Z��  #l>}#r�0�@��C��t&}cط�R
־�U���F��F����n�̞7�u���|oTk�˝���V��
7P��/iO=�C(�[/D������V�(�f:�ϫ�f��/Z��lՓ�ᦳH2�	~��0V-w`��3�K�y��!�M,���:�D�I����������R��w�j����-�a��a|S0y�i(m�u�	�+��E+KR\����@>������{�%x�,��:c�����zP��
J#��K��* Rj-���Հ@��(�����:�q�,V���'�ɒ�z�����T+�}4q�w�����֟C�N�XMz��g�h�%[
go)�˹C�<ꕖ�L~���:����EE#o��+X�ty����e8�{�O��[T�?�$߁���;gS����躁uo�f�5ؒ�2��%:��ȯ*��hAL��u�MBЫ	����Z7[��ea[wK��)���چJ�f���iXI+��V]x��3]U<�ɔK$��s������� �Mb�f�Y�����2����ԯ������SOcl���/�����G(��	��)���]E���NGa�w� f�>���Z�=�KioeD*�T�-4T$�$�G�eݣ��:��.�s�u"�B*F�{�F��B����0����O5����������B��.�Iۻ����,��w�y,��5���է�È�l�)����������H����h�X�~C�p��	gÿS�k�'�X#	�Y�?*I|���,gu?����s6�i4���z=�;�cT�M�l/��DI��-�Z����r)p��}����1oC;��������ٙ�.��Sv��x#��`{�y����P�A۩4�E�:뫟2PO�/�9����^-@	�E�N�H���g�1ˉ:t0� 0�.	��m���X��O�!�R�����3���kܓ̳Quٚ���x�9δ��	r�Z�S�'kQQF�n�7|���EI��I�V��a�-V�C��im���h���K�"�&��O��m
��ḯ����,��U���r*����]lޞ�槀�(a҉F,�|��J�`���"LL�z2̮���˘��C�l�޵��s,�#C�7��;����ժ���/wp���uʖ���q{�0�nbx=f�yp��i|��w�Q����
)�.��t�0��.n,!t_�w^��6;�YC�Oמ���o�!���5��bN8*T�nj�B�
X�
j.k���/��6�>��p����[�����I�&]���n���Aԏy�!�_q��T��fi���#��T/�K�yL ���H,���Q�&t�A:VZp��)�R�����!��lC�f�
��6��+V'��Ii&A��+0�Ee��#|0��F��HZ1����\D����8�OP\���z�k�,��Z%yul��Eb��i���r_���Ir�v���G �T�H}G
��D�폆n�*�*� sM���m	ڭ���v#�g-����f���-��P��^�_Q77��� �@|�}�Ғ��v� 0zqr�t<��c͇�x淎Û:�
W��(SP�*K��QWb{��ۖ���S4`q�F/����z ���!DígW�an%�G��:���"�t#�C�7� m���&b�׹Wh*��9|W��Iq��g��2P���(S�9n�z�&�ȵ Sh��A��؊�/��J8�FQ ^��4P�����QU�8t��?�Si,�L�Q����Q^�$��}��d�P�#_S�`v+1�4���c_$`zM(��Ӝ�k�bڊHO��B�5��o���*-uM�(�/�����5��{�d�u�� �E喰R����̔,���]A���d��:'��{& �<$8����jӤ��0��i�q	��z��b� Ă���Ә�)�H�� ՠ��$�.H.�cZ�
��X�������2h+[&J*ē�Jn0%ןΏ�� L�0�eH��ѡ�l;�E~�����9L��S���Dn=!Ϣ�H��HŜVG�$[����b�9�"xX�7����4H�o�c!*�F�/Β&ǎy�٨d,�Yn"��i�y���p����J�~���D$d��j���?W6L��M(�fk@s���>�^E�{mV��"�d\!�)2��L ��<hQ"S�0���Xja���p�N�OL��])��$*;u��pFVJ�� oNC�E�=�����u��0���u�rz�8�k�?����E���m���@VZ@��ec�y{3P2����]���N[�����g)��,Y�X�qSS�whϒǀ������%���2���h^<P)�rW��P��q`&���PcH	�{�L�IЕ�� K�LB�ӗ��&�"c�������>7"=�o	)<��a���X��5�Գ���2��I�>B4zu�1fᥬƤ�<ܕ,�0���t�*�7I{�t5v�A�c����9)z�.[{�*l��6��"{́e����|B�U���ݫ�	�ss�>'�;xx���Am=�-�Vq�V�s���N����qS��׎�s��	 �c�Hn�ֵn$�řA��=�4J�M�&�N
t��<���[�޲T�2x;1�@��>�O�՜CCAqPƇD�@D� �t䞄�@�E[P��6��X4�-���rT���!*~�a�ɲ/��%D[8�D�\��:Ou�Ƥ�j�oQͺv����P�����q�9�g1A���	:�O�������c���X2{���@�)c9�>��~,,�;���L'D�����k�e�����{^S"�h'�F���=��j����})w&���J�?bA��SA����?�J����A(�t�<iՙ\.~�9keI�V�j-Ι�r$�s>+�C%�}t�/����G��?�o�Ҵ�� ��d ��rM�a"�t�CZ��cs�;D��ڎ"Sl�tw
����S08�x�)o!
p����E���@nm��;��-��+��Xz�bg[�*��E<kJ~/b5\�sW6�����pp\R��G�g!^q�$�8�ݺ�Dun7���?�h����y0�⭄D�C�/�1��k������ʄk���¸u��F�{F䬂���s3�<�����ǁ� [F���P��gm?�.*,�Y�7'�cZ�mmFd��m�e��r��][���Y��3�x�J�nS�����2gĔwo�t>���<7���7��d!�*Ƽ 4v'�P%n�K�cI�w`)�B����cp�&	����J�����C[��4 ��>���S�b���D��L>��:M"],�����O�F>M`�|F�ƌ�am������ā?\�Ѯz�\Ĉ�mU4�R�'��TF�����:���r������+nsv;�4���OOdM�m�,:l!�߁p2k	ْ)�A�#��C�'9��OSu�ĴK�,�.dJr�e� 'm0���iwD�|偊o���f3���B$���W��d�lT٣:�թ�Z���S����V�@6�fA;Q���$1�u��ƨ�,)�81V�]DWNN��A'iT��m�X�×���W��|e.T�N���V|���VU��mm�-��l'�����l)��{�� �����9�)���}��1�prHi�*������ߐ�����Tk?�
�84w'�h��n!��Kk<ջ���ɹ����,;LO�)Oh���;�"vF�y�#���rٛR7�+�6g��ꅄ������~j�3�?�)^������"�VM�{��'z�	���U"��c��+62��R�%�Aa1�	)��ʌx2�,�� $]_2�5�CF����]�փ���ZmPL����`0~'�S��)�߹i�7mr��r�M`��w�㗗�Fzc��ىZ��xM�O�^X��m�D����Wtt���?%"H���t��Ʊ\⦲�y�J}��_�S�$�Z��w�ߥ��,��\,v(,�HjA��A{
d���T��=�zr�x4��_�1�X����!�}��ϣz���A��{#ak�uWs	o@���2!<�	t�o���f�G��э-tygd+A��|X���Եn�����-H�M@̙�4���S��[-�	p�"^�%�,�J=��=X��M�z��D]`�L�+D���.V�eH�%��{�y��O�y�WR�P��c}����y1^�<*% +�@��[_�ƣ����ܼ����3�D� /mݔM�Y
<C�_ō��8��S��7�95�H�%�-�V�[[Y&u~B�E�H0�y��f����Ty�ԋ	���e~���De7�>�a���Ծӥs,���t��"[�\d���7�0e���2��'@�٭:�Mz�.:��~���뛯��z.�����H���Z�_�DI����5��(���2�ݹ>U'c-!/�L����U��|�t �/�Q��fȈ������1P�F���	��b�d�E��10I�����p��l�������|�Fg��L'�.$���l�ʿ�X"�6��E�
�#p�}��]�`⥽�gY�㸸�6�8� �t�p>�	���{]�X��
>�@�y�	v����YE�e����y��H���9��1[g|��T�$���2}�ǎ8l��o&���'��a2+Ӿ�>h�did1l�}��� t揊^���I���"q/��{�����,�o8�=d����[��K��W�-��o�����~��ԍ���n���⡗�fo�ˇƸ&e�9��0f@�i����G3Gu���b�*=z^���EI�i�	�*�~��2��k;�]��"֛r}⯷�`�]Gp"�����qȼ�e�6
���X�eŪ𺋂;`L[���kk�8_ P�%?�*o�ŒY�U��L0��O�2M���v�&��>�.������c�������]5AZ���`꠪�5 �w�w{7��*�5i��	o�ހ�}��$��#N�H��U�Q��OVN����{�yO�M��6{(B]�����5[ޡ�/��d�'z?f=�.��y
���N���پ1r��f��M�e^ݹ���8�=z��X��N�$��ѩ�J�H"�4�ˇ`X�
(�V����Q��I��I�]���	
�Vm��bH��2ۤ=���6:;�Dbp�	OhRQ�M��޿�K��S~H��2;W��)9��W>��EK��4p���&C�ǝ<��������H���>��}��s��,��6��؜�FS(ARG���|�i��C����@��������� �8�'@��9 �@����C�jh-S �cf�@��;^����� ��9�Lba��ƻ��V��=j5ZSkCA�SOA�ri�'<1�L�#G1��sL�m7���O!1�:,����a�jVY����	�?�1��j������1���h�޳��}����$�R�XN�s{�Gn0H�n�Qo̴��n�:j�����������Js��)H!�6����4�i�ދdqB�T��'!����u*� sQ�����<�.#k���G��
uz�h��Nl8�p,��!�����O(������$��G/�
��&H��Qf�a�x5�
|��<`SǛr��lH��yN�E�v��QaW"�_O�.��x��{��815uLzF����'�-� �"��P��-�:??�\w�u��
?�|H�����g��G��	6w�i
�˲,[��G��oW���!�j�ן��WdG�F��7�<��Z�D�;a�����e��8������.I.�w ��f F�j�;��:ijs/���ւ��7�G�EK�0˸7$��Ϊ���W���U���@MA$dP-�g>���/{C�/	G�~3����	�S��HH�$�۬>�˷�B0.6�)�"�ld��	��}�n��U��r���~�%Mw���y�Ѹ6#Q�D�����S��m����rN9�.�5�%k�r�e�BJ��j���H�j��Tk92�f~%�F��6��xi����1S@Q�R��4�~�o�Wq'�J+��Qt%�����������D�^<_�8|����:</'L�g:��`�-k���meK,���a��3�k��g��FiT�����W��2<NE�E�P����K8�-O�rt\�����e>��#�ח%�����P�ځ������z���C�V ��]�:��8m�8�v}f�?b�!���T׊���_d}�=R�l�	�7��[jL�Ⱥ��d-�k
��E��©��ϲ�D�����x��N8Y��#x�qa�[�*����i,%�
"��2M� �uR��;��ۙq!�;�}�>8Z�O�qAf���|dW����+H�t�~I�f�6gǤ|:����l�- 1�l��]\� �M��Q)pu��(��я��^���X���:3t3k���m��.�0H��"UT�X����b&'t�I�TӰ�f��"5��ЬFn�&e�e�t;�UH^��k��z1������7*R� �\�1�v�W���a^��#��0��T�bFB߄�j��C������ŐtH������d��5�#8��/]7޺������5�u�GN�UF� �@�X㥰��3��U,_����H�'"/ӣq�6|���9I�a�ر�X��G
|��S���w^��pd$)ĩ#�&4A򝆊 �i�vN)�,���l���y̱��غ�|L��~�|�}�v�6G��t�-��N)o�ߐ�G ���.�]�m���7n!��x5��n�ۻNЌ!�D=�nuH���֛8�g��zÒ`Q"��8�ƿ��m\�)�3�l�Ba�˽����n�L_���X:�~���>�*2�9������\�p^��n��d���o.Mk(��D��ܮ"y��\V/���D����="��~Ō�۸�}���T�;횧�8�����%��p�]��_��Ep�)M����E��s�����S{:%�n_���-~�qG��Lp4��*&�����?�Pc���r��Z��Fx�h��j�5�����kD��IU��6�Z+xT��ܑ��_ħԩvf)�F︬k���WB�o2�9܍'^�"{��:x��͋Z�`lKT�Zs�ff�X#M����h�:��i��1P7��x�u��}~SK���M�Yv��o�m��e�?M��uIﰳ�P�.\�V��@@�uQv����t��ѧ��s����*ٝq�ZA��%No.d]wN��pS��pP0i�ޚ�.�+xx_Bg�&� �%��W5�2���tHoΰ��h�G��qT����J$��u�d5�Zl�槱2�@��AzU��e�d�/��S��Lk]8uj�-���J�B�qج/w�H�VU����W�qt��g$r�[,��V�H,S9�Y/<�~�4�>��r&Tt%((=��n�lqⓂ�/��h�_��5O�*���n��^��C�ꆽ��� �#n��F-��"���ב���*s��W4�n�=�auhM���gM��i0��BG���uā-�!%+�;�Q� �h��݂���K6Jj��dǭ{��z�v��87�h�v+��̜���F����\NWi�8�UF����o�8p���� @��`��J�ޯh�z.�LR��6��p~N�[�jp��,���J��'M�O[�v�DsT;U�2_��y~_$�PP �,�F��பc�G+�Ӎѭ���Fk���s~�&���F�%���[?��Љە���,�!{�R{/j��($ ��/fX��Y�
�6�wx|�W���~i���
�Y`���Ka�s#/C$�ӵ���2J�ك�������#�S��̌���t�+"F؂�ft$H<�b�G ��[�*��j�:̫���=Z�ܼ�90M\�����w��y�\�"�[����r��S"���Q���7̇�*�]:
ЭT4���A
G^�̏%#��k���+��NXk�U��PS^�`.��B°b!x�T��U#W�1�)��A�������^�K���!�I�2�i����S���0�����6��o!����Ƒ�� �6nO� �;���H�,�Ŀ�?;��z;˹F�6L���$���c7����(@͓XJqyWY`�߂,{��m �U*Gb �D�%�]X��7������q�	�S���YE�?$�%c�������g��!;�/"7�H���!�r����Ao�;�L�X�b�=p�$��w!��Q��U!7�RRx��c%�`�1{������Ψ~����@��!@�͍�=s�O�L�c�i�|�¹f����_';K%0�����_C-sB�&���d��.ks�.+���N��WP9#O�� Udf����t>jg�y��E}+bwi�p�щ��>ƺ���L��/����O�59��)T>\�\M2[5MگL�W�BԆI��
�~����T����P�y+�9v)Ƭt\d�M/PRj�If��0�������V5���|݄�5�[o�a=Ѷ|�<�J�ˮ����[c�B҃����M����Q������~�(�UN��̡����Ɯ`(g�`����#��J��N47��� = ,��Ķc
��]㖚�ܷ3�D.7]a6�r>S�H�a�\��>ڦ�y�%�?i���p�w0�0�h�[�k��i���5�'�[S���.�[��Pj��˸�R)疚�$�m����n�	��:����B͙`�>� ���ҋ�XF�����`���a]�yM�D��)�wã�~��೜�SYGO�Cg#{�=�����R���n��g���U�@�*��gi�z��`�j�f!�k~�%�톧��ߥ��
�(�k"�j�.����Lh��Ң	� ��@XbV�l��<=�-x�hx�Y#��꘰CR#��D��H����H{tQ@?_	����%�HZ���>;�̼#&eۆ$1=�+HPO&K�1��Ϯ�U����`�*�h�9<+���dY4�6|�ӝ&�k�y����j�*�7��H.�i��&pf�J��s��߫89�"�7{N�h"~�l��=��=�9���`� �~�H[X�o�@�<��]�co$��ć��B�W}�k���Jr#}������V,��������M!O�v�J a1�U_�о������@Yߪ헤KC���V��]�u^�\�Y���{-�({$��3-9[P��֌X���)�X��>�O.=�Zy�b���1�����<�x`y}�v`	[����8Cj�@���"(]/�r�n_��G�E�
H"�� �k�����W�����Y|�HnN�ۉ�i�lH娅+�}[4(��b�[P2��Y�(%�1t�E^8J��vߕ�luL�!E^�O�\ �k77r}����C��?�l���5���TY�t�.�؃vCS���pB4���L�X��ۢ��c�QM��瓗N mYWI0D6�:��=�<]�רw!�nMа� À�kc1&>�
7�D�eI�F�pXѿ�V�~]����$��h��ȇ��|�o�鐾"#��5m����xx�\��Ԓ��8�X!A�$���=>� S3�
h��8�ߓ||�ʺ��������ò�k��% Z�o�'��-!�� D��g�Н�5��;���Kj��ǚp�[������gQ�p���e��f��M���0���7��ĩ�;	�",-�K�s�`^^��-(L�)e�Ņ@t���#ƿ�jRq��1����P��/��9�2����'8x�q�V�s0����,�G�L�^��ʄ�]�$m�۪I�n�o�\��)���u�I)�	��O���g5�����ӣ�W��"�ϰ�ݐ�N��.%�k�q�A؏K���1�V��>��B�@�I$�k!*h���Lz �E,7���kc�!K�Z	��q��gВN@??�>m&�E0���>�6�`	4cq�~1����a2�B0My s�6CN#Q��[�(E�{�U�LE*��EqB7T@r�篠�?�a̸��"Hk Ef�`F-�����>/B�.�B���$��c�ix�1xƣ5��j�'pQ"|1��1���^�y�����ͺ�� �[* ���1�JF-9^���OW7����sxӧXqB��2��?6�Π��J�?H֢���W��S��D]��(	ν�����)�o��	���0)�����K������]\� ����ko����q��7��F����M6@��U�_F�R���{��"'Xc�T�M��Tb�e�F�M�jM��܂���
��H�w[�=nC��y�hu/��.�3��Vozw�CrWEU�x!����d� ��V`գkNY]��B|���k�ghV6l��~�3�W�R�G�9����8򰞳�`2�K�:����	Ģ������S	�����r�a���w[Ղ��`OI�!9㵖M����z�����
G�jT��^&����_��wWu�P+�y�*J6��d���;x؟���󁛲��e�m X��p�*f�`�4>w��(�k�(D6�?�N����ծKK�i�.y���s�=¡y[)}����.��6O�ϕ0�N׋���`�0�Y�2���[�rf�D~S�m|��h��$�@�ubEV���<d �0`��� YGuT�{F�I'Mb��$P��7�\&Չh�������p���"�Τ�.���`����ي�>w�5F��R-[�A�[u@MXۓlg���0�^k�D� �Lj�1��ۼ]5����o�v/�-��tT#�}����"n��苃|�X�kL����Ux�O���o��H�'T��@�w|p��+����^Z��x=�G��R�EꬰAB�5�?
%����<���0����oeA.p�&��o4V��J�^Ģ)ܾ��m�t��s���f�,�y�b$C y�%u^���:h��&_�g+ʉ^o�t��¦SC���Ak�,�% r�rG�&��\o3�et��T*�.M���R��Q�S�F��C�E�e�{"]�A�H93��,J�K�|�?��������˰�O2g�  �M��}��{�)�)(�&�� z2vi����o�I��+�/���v~WQ�F̥�G#~�}4
��Ug[�,w��\��.ˮF*y�z���` ��		jAֳY�#o�~��<9��I#킫o�� �	� :��H--i�RE��]Úfw) Xbp=���s	��t@8_N����4��e�r8��IM���ש�#�S1 �łlw���`�T�Bpu���24�oΦ�F%/��Wİو���>l��ؠ��d<�
���~o㦀M�Ј�|\�hܓJ��Kz�f�OQ媿��!)R}��s{
�䶖�H�Z�6� 8��S�:�U�t���1�-��>��g�|�}	]o�<���Ϝ�9��y��{��g��]����[��a���-	�������s��xr������6���e;q6ʛL�fu�+���蛆+�,v��I;��:� ��8��^8-{�����ր�I����S0��������<s \�A~�,~�96��qD ��>��T���z�L�^*��0����Xh��+ A�������Q�T�oY�{"�:4B�[�o�*�cYnđ�ɹ,&��������]���ZVs�OEqO��b${�P(����F5/�"&FC��z����w��6���&�%�(�Ԃ��`�Ήi�4 ������) 3�0�i��"�5ވŃXR4���C(&*ش�%ѪC{Klٖ�������� f\�o3@�q�����qwJQE~�n�)
�ѶŖz*�K�\l�!N�%����>��#u��#�0r�H���"Ǫ}� ���#k@�l��n���ŭ�ma$�F7n�Ye��Q�bd�',���+4
=\��d��n��
�-_Z�P�B�ڋ��!3�A�����qAT��C��@�4x�0}�a�	���a��(��<����@�������X��/���v����X�������NI�? g���,t�$����@�D�uX�P
cH�e�<��c"{���=����Go�����o��7�V!Z&p�7��y#��eʏO���KmU`� �ܼ0������Z�X����F�)r4�N��)�F����~��M�����`�� ��|u�E�b�v����U���1V<�c�c�p"0d�w�y��g�sL��]	�"��p�E��4!�n;�})�\�(�~M���h�d���&���V΁c�v���0���a仛~1��< A#�n��� ���J��k(#}��'X7�(�@r8�^*�"0�b�SlCNȈ�9�;d���n��#��(�3���d��k����a�WTJDiD�6��9]��ّR��9�-?���I͞ml9�l�lu�\��-1j5��cGƓ=|�sT��%����;N<���>�3��o��{ʄC��iNAmŇ�]u�#U�X�t��7�?'8{�������˺;!�$>>S�ԑ����y(bO-���	��f��A1�h��}�3I�<g��S`�]�)>D��ݛ��V��N�����r�|���:��C�3��ݐ	,�upDn>|�|���� �|�V�.��I��r�X�8��׷�SO����Ly����(]��6����hc��
��_��`���0�f&�ǘ�+|ʨ�;����GQk��N�5�=�����Z������u��9���i���.#n&�
@iz]1����.��i�q�Ts���P���ܺ���8N����W|
�����3�����|i'~yA�'���2.^k�u����$y*�:�V3�oMI�̤�'۠d�wq�]���柊3s���c�I{��ƌ�CĒVE�K��o:�O��Ρ�'%��ο9���R�N�W��H��s�
>P,^̑�R��D��z�6A���͉& �9���F� {�qr�Hs���Oo\8ŋѫnw�/p��[���{BYD�����}y�[�r��Ǿ̦��z�#�}�HK�^��|�+�'�閩�yӭ��]�C�`�Ė��|5�`�xr���n���X�N�WR�]a=�
Y\m�f;�4נ��0�Λ�_��)r�{��X�H#5�~��3�tR�8�>r�̇�g��R��Ԏ�Q�YLw�I��_�kOs��!D��ť�Ɣ���'<bާ~a���sN����N�{.�S����=KJ��z|�Nr��Q��V�r2���~@�OU��erHGWol:4M��RC���`��%���*灯{ef�@h,1Op߃p=���+�,�����e8����"~�ź��X�v
��?&�F��e�=rs �n���G��HN�8��5mb8퉠e�sJ���mإ��,���'4UL=�٥��.��}��LW#�c�u+v�1^6�ߊ6Sy�{Xw�x��Wr�8��q�]O�䐽Ɂ�<S_Nz�K�p��bN�>����<�.䗐mЉ+p��i��?WY��w]�Kg�	6$6�Q9P�k�Pmu'4�%�E�����)�7Gi$��#e����X��Lij��
Oe������=��!���u��w��ˆ����~1 !7��5[�P�p�M�{
��X���LPb����bڭ�6��,�&!���W��LWI ��!�M�RyGb�u����n�N����Z�<����'"}Xg�0 �\d�K�S�Ov���,�`�� �ƕi����+Y����*ٍbM}��5m�~B6�d�l�e�+��(gD�p��$L�K�|����8��&�,����S�]�����$�e�T~93T$(1��~�m��p���B	�$���+�.��/�0ނ��0P�EGvGm��Sl�l�I��S��h ��!���6��E��jC�	�~W��N�9��i���?^�P�)��<V���k �ٸ\��!�����ɴBOG1JI#8A�5���Z�7���J�K��ʊ/|�g�b:Z�a��fcQ1���� �QOy�8Ӕ��^C�.Y�oN5F��),�X�V+���L�fg�(����*f#C��Aan�2��J-��@�é��-�'�M�f�Z���zׯ�W���6��͐��2΢�� �A�SU�0���W�W�U��B��������|��Vkʝ]�?�^&/ 	W�qN�>�������f3oR~�7wR/O�$AQ�7,_ME wӄ�GP=�#��y(��P�I����Cؖo���F���P# 6+-*�Nh�r�&L3�t�8=M����,��Y���D��@�iMwh36�J��N�@^9���ʌ���D���hmKvl-�+�-y�������#�S��4J�~�N!\�A�/�{:܃�-���h"�J�Uf=�@`�B�8�/e
�����|�-4kɢ�n�T�9�B-٣��si|M��������آ������7��m!���&N:==~B�^K�!�o4���r���E����wo;7�n=
�¡e�w��p���`j�Z�q�z�����4���P��Q�v59L��)Zֱ6��D������/B$��������w0m|m�S!����n���+�i��pKْ�������ZsPp�}����­�"���\�|�|�>kT-�Ԕ�'���n �a�vBToXAS�f�R]�}%Y��i�����u�S�zTV:ΰ��l���P]�VlF�uP�4�#.`V�vI2_q���~6疭Zb�׾a�H}�y���r�KNPT�v�V�$)��^)�݉�z6j�t��<�<�v�MX;�8�����A�*`°$�Yj�غ�-{b@�$˵j���x&�
*e��>I;�w�����rʏ s��n3R����c;��<����F��Q�v���w� j�\\rYWYݻ���@R���(ht'�^��/�4���T�n�\���t˚k��	%.J ��Q�Vz]1����ox�o�)ߍ?����>U6<�و,X��Ŷ�u]��8N?s�/����惘l@� �+�<�l��x�pktoC�f���m�p���cċ�l�|��$(��X+|���+H�}aN��4��5�3nD�M eΊ���$?���G/t�>�pJF�����D�h�F�y�"��'(��Xʟ>D'���Ff�O�7��v�=�e�>�Fq]*JX]mCU�d
�@�~���t�0��n��m��L���v��`�M�E�ȕ�������������D�on�1�qw1�C��,�'�%^X}t�h�ɥ
NW|�s�>�ΘU+�GCR�OƐ��#������L��K��&�:�U�wv� pxӖ���dK ��{�b=�DWL��gs��^���-�m�)&�{;?uvr�]���B�gjs���hBPR�#,�&�F�9����rȭ�K�@�XBJf�t�S䵓�.��iq ���5��8^ k�"c���:��ח���7�P�2��֮oX6��$���֋����կ�u��3tJB=喓��bt��v�/˃&����ޜ��:\�����_�>A%�vUlc/l����iP�E�����A��^�����|��D�L��֦e��j���ŧ�|N*�خػ��&4X_R��b~aO��I0�=`%uW��YL �� ,J��Y��E�t�@|�hbE�j�#Y���[�	>��G>i�!�K�����	H���'�!֊��{29��ŀT^��+���Ӳ�`���v�0HRTt�q����yi~�"�i�������O}�^DR�=T���9�a�qt���m�"��n������h�!��x^�X���u�0l�^�#�Z3�*70�T���ӔB�n~Nd��[G��% ['FX��H�� �UĦ�j
�xB;%�{)F��2|��f��-���&f-L�(]�~#�~��[m}��Y�[�葘���bN��Ua5��k��"˿d1�����Jla�D��\`_��:1��#W�Q6��i�H��v��+�p�,�Uz3O�e�V<5֖�yg˒���$��F�7ќF[	��%��q9r���[0CÃG�����q�f�FT��N#u�1���r���}nNbП�7���1�5�c�t�&�7Z�0=���"á��M�ڂ#�zr/C>K�	��m޺�	l�xGa��u�R�ԪR����K]KJ�[�P��<���"�}k�x�]-հ�Il=��2�8���iOF�NOts�A�;Y銰֝NN6L�Ce�����a�8r�IfVk�+]�'����Ξh,G[��i>Z��'��1�� ���S���i@}�W-x(K�f=�Ā[iّ6v������)�،��$�8��r��q�v  L�G�]��	�.N遊�;�w�� ދ�WA'����e�5����Ix7�S�B�}��"�U�!k�tb�r��ُ���Ҫ��70'R�^}^��^ [A�'F�� �v�i�jܼ��p?v��:ɨ�!n6��q�2���>�;��Wh�r����=����K����^i�>.V����Չ��Ŕ�v{ڟkǙ8�u�Q�3�ز�NW�uO��і�fL���T�;�}1��L�̧j�*6/N^QD]X�zeS�C8�2�"�_@$=���}�:��l�b��E?��(v8�&g
qae��Q�������&�l}�V[���|����m`GY`	ZT�M/2�ʲ��Ҷ�Lf�H�����=JR����x�r��U��0��dS@_L��
�}�<S_�OD�u�X-�y!�,Y]�K����'�U���F� GF���om#s�}��fF����_*����:.!����_;B��lY�*��/R��+q��u���t(�!d`�(�'rA��V�)u����+���2����ѪgU>���Ck����%�}�5=^cB/�@.��u�-DTh�����
c�SD�d_�.E��]W��u�t-*�J��{`��[���zx�4��f^$�����E`�Jp$��\��#���iX�7J��r�'��U�~ZT����p��b�@$R��.?���;>�Y�\�"��O��f��ĕ�����Ă��#BM�'�9�M�\k����o�!��U�q}������E?eW��0v'P��m���ӈ�D��?������~�.Z��0x��,�wй�&5�1P4���CD��/�6��%�2�P����.����J+���������4���Y�	!>���� ���h�`��Ŧ]�ÆJ�4X��� k���[��t�3jBAMn{���\��X�?b��7����#<b& �F~����#�����O��B�S�'��LCnp�&����9�����N�涫q
�p�
ѿ8.���)-I(�%!fo�|&KC��Y���f��|L��n�tޘ�A<�,���J���ǲ J�@���9�>����������d��tG%	eݨ�Z�,��u)ߎO��|#��v_�!��ZTB���1�bC:����~9��/cP����1��l8���MMU��q���(G��mzƞLO���s�ǦH�� ��S*-���S�h�dd	_��v����(vZ�1��%̭�G�n`��]1g�}D���{�Z����� a(}t���j�����X�d�A_	��9\pz�%�-#ˌ����9{iE�(�H/N�5�/�Eߓ] ,��$yʩ��	E����-}cL�(u��Ԟ2�бM
���A���l��7�xN�9���h7��/f�FƱ�@�83塢��V�b��_pPt_c�Q]�h�3iG��j�b�Y}��k\
��Q�2����{,8�r0�(�+����ca�x�U�K���1���3��y�	͹��@s�=/c8y��z���TSƔ�:o��x �}k~�@����!Z�T{f���e%P^�&	�Z��&� D#�"@!@�җ�ZR���� �і"n�oL
?{�6>��t��0[�����g��%����@��Py0*�\��t����)����!�'p-�iqm�H��~��2Ep�Q���zI����FW�|Rt��-n�Í%��U����n��"P/4���i&)��}��i��K�O�L��)E�b�X�8���"��IF�ب��$�9<��65M�W�\ ��9�3�����ʑY��)�+��<��?�@tN�g�zrm&:���u�`��%�)����n�nH�p�z�יf̋^�.��{�\b_��t���!$,N�`�ccT�m�!�]���0.��)����!0�͵����	���S!7��B4�I��qs�[y#��q�ga�^&��)�o�Pg�"[���#j�˵��9������'���c3͢(�::����g:̷��Sz�����[Ƀs1�&�Dl=�~�R��5e�yI�v�=K����c�?�b'm��TL��9�芕XE���k��b�j*J�-$��f���e������mᣁ������g�O��8o�Vp+z��_i^.��;۰�\|����0��ʽ��=oA�욇�V�Qy���C3a~�9��f2	�erH�cȑ?��M��F�Y9���:�rf4��".
Y?.~Yj��ȑ�{��FJ�)b0������.3�2Dt�g24c�r@�� �d�p��S����;��
^_��,���t���*�$��\���ǆ5�wYc#bF��.�������q�ъ�_��pݵ�����SP�F�ا�1l(�G���mmA'��:����,�8��:pF�z���-��������gt)�cU��"��\���`WJ*�n�1�����Tѱ�����>��� ��~w�"���>2�x�4���A~4)6�͵�˦�! Cta�[F��G��X���S[��*�%l��;�?��1uF��A��N��{�p]Ґ��K�*EB����[�ب������UA��uR�4't���3�,�fDѝ���p*�Q�����v����f�'��I
#���pAN�NE�����$䍜��5�X������9�דnU���I�p@%l3WȰ�|+�R�R�e�"w)v�%���SM0f]�Q�A������̑����G��'VL.�M��M"+_W?h2����dOJ�8Բ��w��&,��壕��:���ǖ���n�Tr�kh$(8| �{e�)�$	GVd>k�P'��m�%<�0PR�e1!�圑b�"4Z�R%����F���t�=x�z�s�pR)�}5���F%�i���ϝa�5�+4��<� �6�f{���+ft4�� ���X�	&�,΋���Qt��[�`	JЪ#롡sx�WhZ"񆙆Qo��$$ķA� ٞ�0�.-��S�������KZ2$����U��9���xhEFg�����
.c�Mk��64cm�4�n�j��R`�,m�*J���U�:���$��a�Sl�hk0��'�
޹�+��C��=��k.���ue=���qo汊�Js�cS0�dՀi�.���A|]�ϗ�+�<r��\���լ%&�-�-�d9�OWr��&��*:n�Aw��F�{E!m���II�G�u���/j#~)	^�mQo�oH����-H�Q��1�~������t����2���M=-X�7�4s�=��S��`�
�[�KC7�o�k8���u!�M��4������v0��]y
�a-�割��'EZ�8�l�DH�����&��*��+�E�rʜ�M���7F>+K~F����A\r'r��&aFц�/`m��Զ����O��8�K��M,�f
�G� �.7A�~�uT�#��Yli�:m�J\/�E��Wa#�G��!�N�k�5% P Q�R��:r���K�����^��V6�膉��ԑ�gu��锎d�B}N �-�F�i뽛��+�'`o� �%#H�&hf�NZ1����.�pc��Q�F�"w�s7'BYX�y�7�)�N0��DО��r\2��A�e���qcP�%�aC��3ԑ���>�M+�}2�q&ū��Cz�^:M���鯛4�PeM��弶��f�*.%��:A�W'<���U9�i��p�f�D�dx��x�t=�������ܔ���JŪ��7��?��ⴵ�W���3Gc3$�EvL��M.
�W����"q�u�\�������g�t&Gv��%�t�4��8��);�+L`^�,��F䮬�X�O}��KUZaʎ)�xZxlK^�$���Z�ӧ�j��N%�0F�8lS�����w̧��	Մ;�K��[�?��r8)��_(�����4Xƌ(`��^:	����ܕ����Ç�#�۪�d�L��Xރ��u�_�6�����f>Iˈ��Q���Nc���E��`�n�M�<�%-��j��R+����ǹ�A����HS�"x�٭8G�g[t^�����G���ғ{��;%~ ����x�܎��h��b��G �:��K����Gk`ԊYEQ����{zuY�Bu@6vh>���Z��k�CW�(B�JZћ�
]aA�;{����%;��"�4>8�eJѩ�&�
΍9-1��:!���؉��R1F{�,l&��Kh��\6t����Qa�H����������2��Ȇ��"���Ǡ�[����]Q#����6���cZ���)��V�!�e�2j�@��럥�7�4�4��� ���;�N��)fjJ(�G|��L����^�tlD�x�^���D�ӕ}L3����-���N�C����ۃ�_��e����}V�*��;�p��*�hv�c1���K��H8�5��N3�[����W{ v��"�~�銉��'��~�발��yƓI��ga3��ʹ�39(�s��CU/�Ll�H��b�B����]���tޅ�s��C���r9���`I,Ij��6Ef�9�����M�T�Ӊj��P9�S3�erY�0�jBcr�sz89
�{$O���`�/�x-K��X3kBS�w �[f����qj�X�Na�T��b�*Hw"}��|*���|����q�h���] ���,m�J�PR,�A8�$��(a��/@J8ݕ������qe���;��|�,��e,K��jǎ����u�4>��l��膑��4	�8|"�1��D.��9&.���}��{�~W��'�e�tal��g��A�*��F����9�2�����O���.~ ����Le��r�4�����	v�1>�ױ����IX�"W�f��u1^�����}�]��q�j���b��ˎH�Rd�n�T��/�K�ORG�	�!�C(�VX��j:F��4��[OO7��x��}�h����Ƌ�>�yQ3_#��d����(�u~�cȚ���ۨ����x���q	Z�p��Z�L�)I������b�"������r��A��=G.��c����d�Y�E/^�1$@pR�LiJOߠ���N��6�&���h�@)�G"y�6+?�{�+`'�/�C��-�l�L�8���M`�gxۑ\��49�n�徊��H4h�����ۗ����,g���G��dB)�W�p��2\ �8�����;� �5ݛA����E!U�����L�^��.��;�kӷ{��.�v ��*��_@��Y�u����{`kX)84C2��z�5$�Q�`��z��Jd�9}�ʡ��I�Y3/W��*l@RJ{$5�E����k���׃e #L�^��Coέ�"�C����&v>�yq��)1�b�ɂGW��܊���83��K;'V���b��sxy����r_�$arE�'�S�"=�f*Q���@����,�m���H���J�"�uv����K45�0�r֓י������y`p�Q�=[`kp�L�p�]� �+�QM��<VӼ�F���_&kg�ܯ�.�me��v�=;j�e�	ђ�So�GN�>H#:fv�_�H���P(���qh>P�yϧ���|�ꉎ���R��N���%?`5'������`��(ϴ$ܾ<�8(i�R�zwW�l���g	��KJ1����$<3 �iĎ��ZE�
L�(��MYq��E���b��)���E�X2�V�(����A:Kc	��4X� ���������wsH���ƊH��@�FwWy
���"�Vh[��_�:�O��7q�M�
B��B98�֥�Et�F�2^3]П>�4�3�z�M�S��D��g< �%
?2���o��k��c�ڢ��\��i�8�y��v����
��`��G�<	F�͸��m�p�Z�8V*�!E6���x-գ6���o�A���WA��*��a\S�Z�L*�8x� ��M5�D]&�$!VJ���~�~z����Ժ������G�_P�γ�F�e⢀DJ�w/�_?<�Nj�fX����;8���9;~g���oZ�T��-��	 ?�y��iN�j0�i�x�<P}[<���7z�NGH���(����)��$��8/��ޠ����9��
�����k��#@���4՗M�a�N��Q�Z�|UEjKR{��w�-�"�F��}���Rvg	 �
	2)�?z���$����UN��!�"����g�퓻��1��V�X�dC�;��0G2�+��X��J�̓v�p������D���[5�W��;�~��Յ�b�phH��Sd��C��~��B8sF9�Xm��&Wr�H�L��5\רL4���^�W�.�~ �3Tǒ�7I�^�Vͭr�s!�a]�� ^�.�:�$crI�9}o�)��%�;m��?w������b4&�㿃�S��P;c -~~;*
��<�?(�-�]��\Y|������N~���`�?T=�Q�2�|@�=`���S	+�}�t)+�Nj\���|T�y������E��	�c��݊�xy�N���t6��eG�}�#I1���6�p5�!�����tnU��P�q�2�ZhP�G��bN�IB�C`�Tn�gr�c٤lqf�����;��aʲofoH���]�a5�k_�{Q� d�\xS���觛޼;�U4~���YK�Ue�q(�z�} �������ˤR1WN�/�����^Ѡ��zHjGH�oW���66���鸽�8�IN�f[#�*#KEig$�^�����P0���6�4��񆵳Q�J�s�� �2ֽ͹����XQWk� 1����աbF�3��	�@�\�N+J�@k��W6��n��дV�a�u���r6�؍�1���⮷g�$�L#��b�tp�x$h#r8paq���Q�*�v��
FL>5\u�Q�`��Jy�0 O�luH�ȥA4�g�B���[�U��}�(gK�(��/R�� X9�ye�jv��>�K��ĥ[���0�I�L��dڰڑԤΚRś�8\�����z����w~n݈ş񛆣S�8�N�5�Jh�� ���w�đ.I�9~�
-��iZ'�	���$&xn���s*��d��=V5_�:�j�&.\o�o���O<E[,i�~7޿ܶ������K�0\ּ)a2�L���Їx����^ F��z��v�1`XT�]���L�s��?����(P���	�OI/[oL��\�W߷*�ꌑ��%�&�42T�aJ�:�o[�sX�[ibU��3�/�oťdQ���ѝ����G�Gt��۬:cק*d*w̴t�Qu�!����Iۜ�[���L���[PX��%�*$5��M����$�}׭(�� �f�����D�oK��0aN�
q��H�sf�na���i�_�M�	��`� ��h�]w���b��QjQ	�Q�{�64�F8�h���������Ӆ}���_�Ӱ&�]�t��������O霅�j���/�-\��xlO��fs�J5�a(���F
r5*�����Ӻh��7I��n뉣��.5�������iI�}��Cto)�qɏ�LOPz:i!�N:H4�ڱ4��k��L�[4ҏ�߀f��
ZU#�M���d@BE���� ?=
�䩟(QS q�Ϧ���W���p$ʤ�-LlR�N�2Q�U�-���:� i���`����%����8�DͪT�r�'Z�!�[���H�r�H�5�/k#
��E�6��~�t�u�%e!�x�y	OT,���L�;EЏ��vs�Z�7���R'�N0M5]B8�>�>��s����v�.0J)����� >�p��,s�n*��|L���/,q�b�\�׹�I�6���rwe��A�s�x

qL�W�U�L��f6�����<���@<	O6�� R �ې�S���_g��D!�T�����aڮl�$��U�s `3��s#5�VtB�����l�4���H�_�r���{�Ct�nmj���<�~zd�����r�k�,�Qr� r�ܿĩ��^ �*"9�-���"|��궟��Kr���`=�ܙ~�%=��,��M ��k1Dl91�l4����iQ�/S��� ׃&�s�g�?�)�M>}�H�D����Sϳ�����y%׻}��Y�L��]hs���D��x�A
ӆ£��S����G��-?�uj�6�8���<���H�S���s~XG��b$ o�o�E?;�k�����)�%�	谎j����=#�S�h�|���g(��\O9w���p�c������h�&4�$����_}ſIHu��C��������b^�¨�8��5Upxw�[�q�w�Ǉy<�������T��o�߂���'��+��6�'d��3���(����!I�P7y;j���T���Ȩ]=!Q�m����ޭh��Jd���.��pX?g;P�Ǹ�������&Q�b�6����r�M���B3�X����J�..vט������k���YG�=��ԬeI��r��v@d]�@��N�g�'���{r�K�_+IS�_��(c�#3"�={a��K�D�����#���'i�kA�۶�o�5kI���1�i�+Ɠȓ�%ى��I�9�R���*+��G���|�\ݐ��N4B.������n-�3.F�����
E��=���Խ`��~���ͦ�ů��dWgda�<O��>���_����m (- w{���Z�A�I�m�MvIP�U���4.Z6��wky�3�"(V�DuS��1���s�R4�jzҏKq�������V5{̞������/س���AS�������,%%�6����R�&nGu��V�zD����"����߉Y��i)�9�ʣ�4��q�#T��l��ˁ��q׹Q����A���hW��A��cn֔�ϔ�.X����T��P�74h��\��}Q�y9Q�?-b��)ܾ��IS���yJj�wK;�k�T��	�]+��7�~�z,�ͤ�CE���w��\e���	�qh���MQ�"��wڒF�Qz�������=�>~��"��،_�� s2�k�i��ח(�ջ�����BgӸ�\FbP2��4����"��F�v �;�a���ERš]�f���"�ȍX��	B?/��XA(�#�-&���\J�l��`��Z.-�i�k�*����__�ӏ1E4�r���5$V�` 6k�.����:F�����g�=�����پ�����t��fЄn�kh�h��[j�ا�0��9�[�N�Q��u�@|��z^���Qc�8ˡ�+i��P��b&Z�s�H�@��Ne<3J��ABj�Y�H~�{�a޽a�e˒Ç82��N7���B}�uGЮr8=�1�����;��%�)��V#QK���~��՛���WCe�n� N�u&��=�ƈ�pP�;��A�;h��te�Ł���Nd��ǽX&����Y*�Ǣ%�s|e�(bK�+ ަ2H��bx�3�F�n����(�j_X5:��v��RP�O��j��:N+l��{�3/��-U ��%38i�7���~7����E��A�T�'NE��WY�:������O^~� �$$�M�R�p��%1��x�M|��8�����L=�j�7���kB��pgٷ�yU��9dm�؟��f�R�(^��ԸC�s�΀  ���`��5<oc��D���0ȂO�p�!vC�w>��l&( I�Hy�XZ�EPfN��(]ְ2Ll�1�ʎU;��r��ɝ��x��#�Ĵ��)�m�����cN^��H���#mZ�N��/��W�Ö(^;���*")}��m* ��2�M�(a�g��&�a{0�4pW'���=sW}�x�����n�Q���Hlm;(<���v��ϳ����C.x�ۋ���pOE�UP+r�_ċ��
i����@��U�!�#T'@���hx.e\� ��gR➅Պ� ���/��-������҅�Q�"�c�������	����,q�t�^j΄��V���a�$u��EL,oft�!Cu��N�K���J~��z��v����0B��yR^)J�j�-�L��ʼ�Rr<��>A+O���v�A!u�� i����V{�X,��o��e���5NZЯ}�}���p�������PŨs[y+��t�����Ic{��y���|����V�:`��U��u��oae�/s^�\�Q`��7�:�H�jػaf�
�Z�ej�;hO�fВ���Ⱥ�`�?��~�>�3�]Jz9N{�\^)J��Շ���dũ�{=�/��ŧ�5��.�A��`���9,����]�?Z��26��隧F�e�ДĿ^��ua�������Ј�C�G �܄������"x���ة�dH.(Jo9j��j{�`�6��x�Z-t-��+��	D1��D��I+8bG�Ǻ�L�B�[�Yی�v��W|)L���O=?(��(p�ew<�9�^I��$�Bz��;L�j�Ȥ�?,J���,�QX-��~���g�'��f� B�$�K��m:h����K�֏7�{ox^�!3���j��k�D��?w��4�"P�(JYT��5`�Z��ɐz��Yy��E�>���V�����X��q4H���q.��� >�8�¾Գ�ڸ>"R�,�>��?O,@诅J��{��܂V������`s���s�ۼ�C푑���>�,$G��9 ��{��;���jw��gy�)��x��f��jt2ġ?1s�{�K3���Z�X�E�o��q����hc�,9��&�;,>HYy����<f�LT��ԫX�U�or?t	d�)k�0rp�Y�Q�'�$f�7��f�����V��YE!O���i�w�p�Pr��*��4��Tl.5�R������h��� �M�o���G��Ӎp8-�wj֐dR�F��_�Ji�>�~Z�Y�S0	v�eZ�e��ʼ!�5,��2Q��}֠��^�r7��Z���W��8���,`Z���X#��0�B�)osØ�t�aI��V2m��%~$�+� 8%�����[T�s��@��]�-�B���w�%߻�9�r,f�dcj�j�F����RK�v�����2�4�6��K�D/�j���&���ɣ�J}���T�m��:���m�q��Fߙ$�����B����8��S>W�g.x����/d��bh�6���s��#�nEyԻ��E5�Tnf�~)O�""���uA7D7�l6^��Lz\�M��]1+����KB�ӑ���`u4�w`t�������}��q@b]t��K'e��О;Hs�y��?��쀬/��bl�
B�` (��k�0�=��XT�!rR�$����k*S��$XP�q��/�ѯ5�~> 故�E(��������b��39z�DO܋���͒����8��R*�X��"uF�Y����[�9o��E�*��Z�Y��ת�G�g�Jsl�cK<������M}�E_����m=�.����!v�`W{�����y��KE�w���D�;(m��ٮ���N�L&���m/3�v/,<6����|��J��[I��o�	c;;?j�h
w*b��"Ա��C��:����$����&/!x�Q�%L�5kp�&���q������w	}�3�t+�{��?r��F���>���f��jΆ��G2N	� �%���83�G!��	M.{�W����~��ω�UW�9�i2_9����\� ���.	ӄB��#�j�ի��Y�KlIb��*���yf��A9;�$9�R�gD.I.����cO�f�����d�HV`��*Q|��*��'
j��Qi6�*��6�����g"Y��`kqw 9<�S&�=��9�h%����M���f��*m�D/��.��H�-i�U��u��f�ʣ�o�IU w;vDҊt�f�~�Y%"�0�D���&��1����}��s�s�{`���6F��T.�@m=t�m�7Q��L��kN��ʴn%��LAG@k�Du��z?b�o;�	#r����y�n3=�s9r`�[�V���ѡ�Nj���V��xgC�T���q��J����r�7��k?��#��yR��K�b�7e��7�\���!�<��Q��m���
��S�f�4�ݹ`�����^Fm u���|O�8G�(��_��:
�`�U�l��us9A�RE�O�f�lA��n{|�=ڎ+Sv��_%��!����w5K^n��I�y0���Uڣ��X�\6�g��Ҝ]���7�m�8vՖa�sD9�7��������h�r�KRCfj�H�������cb�Ҫ3
��0�S�	߆����{ nR8Y���lEh1F̪�"5E�X�F{�n�J�ԭ��M"��w�F.��7"=*�����|c'��dEC!�L�'����?�R䒼��z��5Q�o�4�(p� �[��K�sŮ_W�e$�p�q4�[8��|�d��ǜ�M`��'��`��4CMh`�3Y?�ML����{�H�({ұ��'W�[���:������Q�E���+�s�]�f��׽&��&	
j�\�tTJ�����𝑣�a�B>p+Q�VrK�<C�O��B\3���J���� ǘ�>77 r��Aj�r�q|�D��I��/��G{�)�KĘu��ؖ�d��`�&u�NM� �$�T��Ш��!��~I|��x��2�DB�������)����oee��\�E�g�\ b�Ue{��pB��VP���5NXqk��H֕��}��C�Uь���QH �:�r�]�|�r8X��hk^�8��Α��؃ ר�e���=ҭ��Ǘ���f��?��+<&]pzMzYO밂}�9�\%�q>��;���F�A��y�3�R���ГE�ȱ$"�{b%�:��u�L��ɟb�o�w�e������"&��@�0�e~Y�t�6l5����<ϼP@$v�.�M.v�N�N��c�橴ˇ1�_�%xc����/�F��W㠮���"T�F,����h��lˡ�L���>���;��8�P��[7da����5m�L��m����:�n� �|�I�Ѕ�i�~�[v�X���k����[�)u j�~��z�d�����c�F�����,�<	?��ɢ@���!�w�/��O�B�w�i�?�ͨ�|hu�;i�0��Vè�y!Sx<R���)�7W���E��� ��sQ~n������gZQ���q��U��@��#�PȰ����O�ǌ��
�&a��o8�5��5y˩��X���8
g���0ա�E�����;���Y6x�I��1�Wb���fqSM���i 8�f���R�+����� Q�LE��!/#�է^K�hvLc~/�w#�� 怩�U�i�N�T�6��1xaN�6[k�L:@��ѯS�Ώ�����/��!����83�
�����>;X��('x�2�}7⋲ي��c62糢5�u�k����κ�3�~���MDQ��j�1�l���Ł�����'��'��휳���=]����=`z9񣥊��S�u�;�ȪSǚ��g��K��*F���ȋ7nR5������@�)��d��mD\��L��@ဉ<c�ݖ0�~ ���d�M:�U|˜�q��#���� ,�-me�=a	+������V0��*N*b�Q�Hv����8�0CY��ŏ%��N�I��<JPi��ǃ^M{*��t�^��ƙ��KH,�bm'O �ׯ����5�M�k��=>��hL��!�/��l<]΢�f�B������[}���Vb�ѵ6n+�R:̊�����B�<(�?o�9���,` uQ=T����=��������>�_��P:�Q�|�)E��$aX��>�ڪ��w��c�C6�Wav�$���\g@��S��p�U�d�1�*��!A�,q�M���
�� �1V�"� �v,(!�sAȎ�� �ua��x'�*ZE~\�����m26?N7�/��{�w�qb��E,TcaM)h` "
I�4O�א�w`~E�K:W�
�kR�J��W�E�z�������x��sk���_8��&���М`2���<VV��N� W18����LG�����Ҟ>׵�'����L�,V�R�r�)�۲��D����'�]騯'�����N,��@�?åWY�[|1��,8qhv�h٧�r �Ȳn� WC�DK�|��JF&���迕�Q�	R�kN���Y���ЀLB���ʱ�;�I�nm\|��\�Ax�j,y��N\��6-�7����ʕrsh�r�aeX��Hc��S�:��(��[���E	i ��V�������Tc�� ^|c��ئ�$ LR	z�sQ63������GiI��WO�/��k�u!4�I�R�Wj�M��SZ���7��OY����X�)�����S܄����CM�k����R������"��p���1�g`L��s󖃮u��5��dk���d�nE�l@��w��#�{%�$^�񃍑ٻ59.q����IFH�f��~�@N^9R-x�y5��%�q5|��._L�6x�	�v�ۮ������`��{bG6��j,怉���0.J:>[� $�k'܁U�����N���@�+xeǝ	���'Cy����nޯ��Ǵ+S��fL���b�[�+��R�j �eC��΢Ϙ2�z/����ݚ�I���G�q~�3>sƎz���'�/�	�SCFd�"���2�q����7�^�4�V�F��`�IZja�Xv�*=�Q�� n���QL]2��[���F.&O�T��h	e��bA�� ϻ]�2Ws��R_(;6�˼|~�5�,�oVޥg�+���`���mp��d�W�!>��0��G�Y-�s�
��8�Qc��ܰl���/��L'��)f8z��4Z���<×_@������o)�58�%Էz;�y]�����b�q�Q�V%
����`�5�I�:�bH^����=�@��D��~0���;�O���C�Ԯa�Xƚh��6�a|���ե��q�WhP�*~�`�S4(h��}S�t��%mDg�_����U�F�	N��?�3����t���2V����#���M�wۓ��c<њ)E�g0�t�f"_3�ꃭO͞�e��?
�L�j�3V��qǖ�-QG�����I���U�;��8XYJk�O�Hk���z�T(����U�XX�c�h{�So��(J��iB�U�4����d��'���reyi闺ުeH���6�϶�qs|}��ٓ��L����#d�Dq���-[�s��[ha�d�W˹d*�g� +��q�|���$�[�<�+�� F�yq�o���*M��:�{E�����1t�嗟-��K� ��8z�e����W����R�T��9�W,/Ox�z�nxտuԪ����� �^eFZN_I�'F��i�U��H�Uu'�m0d���Xu�j1�+{���ѼhSi%�'��MC+ֵ���B�F`8�S�I��]�{�jj��9�W^"y��!�^����"�f��߆�
����{���F`g�s
�:�9�1g#��&Z:��O��~q��UQv��6`��/��]L�|�� ��U���II8g��ql���J�����k��-R0q�4Ia�đ�Z�S$C�^���a�/ogyI$���j�!��u��uxj��$��A�f�Hg�Wq �&����O`��;[v�P�l1����a�_%~g���R�K�9��z.?�f&��V�{���]���E�A��dMe�7&��>_x�g8O�[�
Py�>?�a�y\H����X�I�͖� �����'����6Яo���~��"X�m�B1�
�.��Ʒ��W״�\u�9���#���,?f(z'�!NX]��c�Uڀ����j�U&� "��}�p�>cii0��ȯ���Q�����Y�B#mS�8z'a[�1�Mk��O�x:t��;v=`�,۱��l��h�`���*������	&��Y'0i� >�A�q픥�:U�2`�;�����"Rg� @��:Qa�ܡ�Ƚ�$��讴������9���{��zF�0j��O
�A2�<�?��u:�ig*:���I�E��x����oȪ��J\���(��aw=��i%i@)��T��6�Ѿ�Me��6 ��2hpP����o�9#hN�r"�8p�?��y@����D���5�m��P�(�h��+��̦���$�Va���;��P�3'E;�<��w�}��O�G�
���h���PJ�P�l͚K{[oY��������ȕ�9s��}Y�\�nŨ���,c��u����:��c\�{����J�2������7���{�l�_���=�Ƃ�B��\�l���� Uo�X-RԸ�H��[�,�� O�}o�h�a�J<O�;��\�^�f��￨����H �QS0�Q�w� �>sdKL�t�3�G�>`��v�c0̋�!A�	.�9c"g$B���2����Won����X�7o\���OƁ�e�,��r���!]�m���"�h �f���'�Á��kL�>�Z��Ou���J�B~��W�ڶ ;�;����	��G}�O��E5 )P�<}��L{Y���Ioa�0��7�A���U]�mA\���J�}�X}�����!ME�{���'��+Y
�w�բ`�)��%|�*Y�#q���}�6M�MT�7�k1�	����~[�g6��]�JR�S��1�4 y�,��z���3�g�7Is=B��p2�i�}�+2�;ɳ�����$��	"��SC�B���y���0��&�X�km��Y_`ȿl�M���;�a����p=�4���~6��Z������I�	V�i�4e�I�$�J����'��:=���ۢ���X�3��5��u�f5���nl���M�h��styD���=.x�����ЗZ<jt��=�;W�����2�j<��,^�������@n�!Za.N��+������Nf�냒<����=���E�)?L�Ƥ��������P�W9V�g̼ e�+
�L-B/|�"llF_m��
�;#% ���������;1�cP��Xԉk�Z'��
����ȵ�7jS@�bqs�����C$��~dIg�j+�-�8`!x��~V��ݏ#�S�u#	Dp<G^�l���:�
��\�
eC�ڽ@Ĭ_�z&w���!��B6XR��A�^kB��rsǲ0;�#�ޙ� ��Z��&�E��GL�i�97��\�o�޶C����~O8�"�ҳ,d�T�����݌-Et5�X�3�XDr���#:���_��E�i1�^��6BF��aX��Ќr��u!JąK9�9�ͭZ1T�6�i���JlR�E��$��pRpA��RmX6�^��˟�V4�yd�WjX�>mΜ����q�®�v�9�������~;]KYlfe��s�4?������]�qˠ�x�d���F�3��0e`�q	��W�v�k�����J��k�I
$��0�|i�
�;o|tY����������nX��4T�о(#֜�f�<�>��X�nb��G¥*����[��?Jt��P,�to� `t� ��po-u}|J��=�/�b��Jy��iGA?��Ѣ"�?V�9F��G��7�W�3�JદR����=up�v�6h��y1U&'�۠�blL�i��7��[��Ӆ#�u��V�4tG�
�_�bu��KGH�3@�<��ai1�7,�a�TYv!j_�H1d�ì�x����z��n=��!�E� ֺ�K�5l~�J��F�S�HJ���D����.	iտ,��+�B]ؕ�����'\ 	'�]��q�{݊-CW�a�4�3pm|@W�M]��Ƅ+�c���&��V�2�)8���[5ч���H}[V�!�e7�[��vV��F7��h-<�q�B�f�9u͏���p��ڭ�n����l�����?,��^��Ru��Ӌf,M8����T��yA-lՃ3�w��7��JƟ:E��s+9�o��|��*g���{�ЂZrON�Ux#�O ��\���z���_G���!��e�ٓ� ��s_p�I8=�����7-�*��g�eV���΍U
���i�ʄ$��/+�2��K�z�;w˦��xꈄ\�<3a�?Bʍ�|%�0�<3��o0L�2��Tܰ�,w���Dxm���L���Q~<&n\Z�6�{����y���h�L�%䔫��]F��R~=в�wc�!a�c���>Ac��5 �X��&l�L�8�@*鼘�{��&���
͘�k�	�U:�Q�aG/��w��V��R��g)70Kjc@�}�yJgf�$,j��j�P�W<���>�HS�y�o��ĩ4�2Q���:�N!�ש%9�Z{����[����5����ص���^����m�9b]�Gz"�$Z]�,8���Y�4<�ܰ�GS#�_�J|�0�h�d�~�ʩ$xr<��.�B��t�s�U��Q�y�+�|Gm�}w��K��M/V)�u�Ȁ�v	ʂ���B��W$L'��z��/�	�_�f~��"�L�����*�X6-�����9~ǣi�n��Y�t�f�tg�����:��O�$��q�L�����+�	d)v:���[���d�>�hbxs}�а����:�[��g�&�q�c� 1�9>��Μi�ڐUCt�M����Z�����w�0��g��Q���p֍h��AȂQt��#�wqR��&���w��ɴB[F�J��~{E��
����SCB�rB�Q�ç
+:#ʿO���qQ���y���j/!h��v�tP�G4M�uB�u�n�0|i�R���0]۞�:����r }�r��Y��`���1^pt�yD��)_
,�(�5j�����ϵz����B�Z~R[� /&�����7V�VA�p����>&��f�^M�g�?������N2��#ӏ�4�?SX����^�$C;9{���z��M1��/?x�z��}���4'�8`,��q�'�5w]��v�v����sX���3徐��K�*�h)	L�M"������kQQ9�ѿ��_TX����3�H|�d�tKV�otz���4[�gv���9�M�ހr�x�K�na���=�C������y�KW:�
�<��v�Q���n_����@�j���&-�r��������(S/i���%�X��{��ϰ(��ɜ$����_ǒ�b;�Y��Z�^_�D}� ��/W�L�i���M�	ڔzu5�>z[6%�1� ķ6sͲ�-�v�B���N�?e�?�,����kYA�T�@K�<�y��o=KU�֤F�UYԍP��q�i�5�}�4��G�d�&'���<E�T���L<Y{��dV_^�nϡ���ņ��ж[& �31~z~���ߠ�^AC���h�t9|+�|dt63����A�pu�ǝc��Yy5�'�-F�i�i����g��BV�J�Mz'�cL UnxJr�׬%x"��2{�G�Ģ&L�{vc���@��b�ۘ��)��Ps,L;&d/�f������|��a��k���DW��%c��K.a�ߝ�{:�%��ɺz0z6�3(^��Ǫ�=�a���e��7a_C��J�B�ʏ�i�n��8�^A&�Q8�d�J_��B�(} �7�����j~�'I{�V=R��6�г��P��}��c�/���2Ѳ���D��	t5�t7��������R�
*��.���P[�����-�k{�ڗ4$����)�u6��'<u1�چ�l=c݂h�A���jȘ0�s�������J����K+d7<�A	���wo�b�y!p�;��u��\��J*\���^�x�\P���oNN��� �;�_7!��� �
@�lD�aAW@+�܊�i5-:�\��^ȎX�wn����Ib�!�%=�ہX
�����c�� w���Ř4����U{X�v���.�"�W���Za�<z8��X��p�*��0�����.A�)�/�L8s �W�-�V�Q�{��J�x�(C�-M�}1�ĩ�z�`S�(�M��f����K3o��#�#W&��B�K���b��[����XUK�q�|���&�Od��)
_�ȯB�WV�}uy��h'I�y3�#Ў���sf9חG]�;ྤ��K��]/i������Α�X�~�D�%V�{������o%R�XS�}�''���>�m�b�N������lo���#����9�#@@�k77+i��+lCI���.f^q�������� i���h��k��XXn%��N�\8�&������܅�%y���f,�{���LA�ͥ�X)p��HkDw���a�Y5p��ws��f6��pY�|]�����qطc¡NJ� "�B�T�{m��5���G�'����<�o�-{�+��"���`8ݴ}��%��Ql��<�hD^�\�ta��{O�`���&���	1R0�d�P�(t��c��;��'v"�`�M3�,t}Dú�ZĤ�Q��tW�&Kj����MjE��62��I�J��T���^ 4��b,�"�����=����r�}"Ź�g)
ZN��Ho-��b�D}Я�������9k������/��d�����Z|�'�Z�-�^$��kݧ��ef��Jh��5�2�8Ҷ]9���,�3&ݮa��VD�1��~��Q)X)cPٷ5~~.��1�cϦ�"o	����i*�'=S*������+���׺��4w�mY� �����D�K&�Q��[8��@��F��K��"�G��ãG�'�>��HDt���@�^��R���h���k�<�'ġձ�J�,���A�&`ʌRi�˜���DSf?mqQ���2��}�ڦ�`'�3�#�s(Z��$r�A#��&��d4�jA-b�)��%�k�o+��EK����"�kW�c�k��S�������G/�"۵��NϷ��q���	�ي��^r� .�G�����X�y���_`�j�B���[�tn�|�,`[;R��G1�+F��i�G�.��)�Y����̢s�S��o��=�e�X�Z��g��t�
��%什�$�#ǒ��J��-p���q��(\�1Պ��I鳘V`�>�Ö.�Rl���  �+��̃o�;	@�MG�Y���W3��4B'�vIA P����B&�(H���j	��E9�uMR��ez̜���$�;}��{=��$m8�9�P׏_"1ᐮ���`�>܊$�^%�|�_óMI2I�n<���T"��{ƹ��*��\I�P�kN�o�(����ȴ�\�Ԛ�Lhk��}��#A�jG.]�� `�	>�Ў�L�l������W�,w�(��>����b��U�1��Az��b�=������TF�P�o���k�g��YɖH�i��k�1��|Y%�|'>�&�]3�¶����J��!MN�.X%���%p׼�M��s��k�h�j��AX�f���A��{ka�$�[��> �=E�H-���K7�U�&�~&�Aф�'$�tJ����ne�^�8��B�C%��:�����8SG�|�燥�﹚�sz�3�-+��ο4��-jw���SR���[G���tެ�y[�Τ{������RF	��@O�w0T���0fd��6EQ�\����2ʀ't)�fB�h��"8,0���6i�p�-��B�_d�f<��l�-b��5O�}K]Z��č�Ě�_Ǳ[o"�Y�uye>:��6�+ϥ�}����1�e�]gǸ�'R��׺��_���}�Cج��:��y��iꐵ�q��7P/���:�����r���C!�w;�x��6��<�H����n]>
Q�l{58TN3���^0|ڿ�<z�$�-ya��U��XF�O�3$^���b�����X
�N�IŹ���r+1���AKu��Q�l��uթ�e7�Oq\y���va��a猨�|O�g�������(�����J���ћ%�5�G&��1c�k�d�R^Yu��W�Ť���̚�j�h	����,��u���a�NJ�a�n	\�;�����߿�7:HƷrv�tƾ_�����j�Ŝ�� ̍��P�c�t���q6��l@�j*$FC�1DJOzz�J��t[�iT�&FĂ��κ�%y��Y���8.���[�d>I�Mh:K��b]��l@m��x�乄짷��<�%��v�!~ ���vb	���]�ۮn��rZ6v(?��M�|6� �0O�,�1��|��"/��m���dL�'QO8>�2��m.!�N������U܏��,f�]5�C)�6�!3��Z�:a'�JC�=��X^�|�ICv�^�f�A2��=9:�~ٺ�ӥ�P~d�r�����M+<JJ�E'C�����k���'q��:�@�����?�ۺ���+�(�������9n%����Aox	Ks=y�Ъ?SHz�� ^l0�����Y����+LD��=&z�SI��a&q���f�#L)[�5��|M�Ě���H�| Ĳ"I��?8� ���-Ԃ��]�뜂w��h��A���k]܈��!��vX:YBf�M����iIÉ]��I�7��6�RmP*��ҩ����\�/J����7���¢*��1Zﰕ�~��`��U��\W��B+�{#/��}��͏
��PWo%M}O�?�y�����'��.���Sٰ���y�N�~'5��h�'�O� �A�Ԟl��Z� ��}���d� �������r.���AU�jE�2�e�~&F5-o|��qńqAXG�KWUN8Ob�G�WN_�7���My��ӃN�m}�=jD9{�#*��,㔣���ki����F\?hL�;���2y�v	�-�a���O�w�V~@���+�K��5���;9X�G1�G���];�j�{�rKh�=��$*l��\�{i9�2s�w3�i��1�-�H?�gT��T\%Z?Rm��l�)*���r���e��F��B��U¾UY��#2�M����Й���s�Y]�u���H�v99���%����+>�9�����ܹL�Rj
��sMQ���5�౬F�>�&LFݪ�g��G���-qT��h��Y�z�����l�9JR�5K�o/Q_[�q���v�w��}�Bi�&����Ax�!s�\w��*4��*��Pքڽ���Z��Rѩ+�D��U�B��vK��	�{-n�Q���T��l&�j	�;��"d��+2�%ԱB�(~qec.܉��I�ǃOX/c�
��k�lq ��o��_1���}�Q�ů���Y᛼�Lv�S����܄��2���&7ξ�B?֕!gȁ2�2�[�K�Yz�pٷq8�q�2bW�����;�`"n�śx��A*�%�K���$���!�ۋn�+/譻R>��񨥽�{���5��_j�l���M͹���P�}F[��E�h�����W=���O&c���!t��l����S�E�Y|]&�j���2)�&�ogE�p$Ї�WM�ۮ؜��W8�?���J���c���0<�f�xp�$p�������y��$�5�o+���삋�pT?�Ä́��W�K:�
a���n�hY�sŵ�	��\��yͬFd��eg�,y��$��/���9Ԏ{�o��1�D�_&yr-$�h�*�%l�����9&L1��; :��'�a�jg�
u]��EW������'���������c����SG��BB����y��h��c��#v�WL(����&e��@DM�t�>�(����*�	u�n���I��BܦP�\�g�F��eBQ��D+�]|����J��x&k*���.��4h�P.-�Vr�[��gp:��e�l���(=[_s�Ǿ�c
 ������Y�&�s5���vj,R��Ӹ�L��l��v�0�2�p�9��c:|�EǄ^h��A�Q��� kdA�j��f�PXe��P�N��:��`N^1v%�n��\��H|%��� ��#�ﯡ��e���ny�o�wĀ�ly;W[�� }N��'���m�!�N��^��Q�Z�Y��?��u\z�Z]-z|Z�ϊ[�m����.��O�)]������\P�4���aliSR^>�[���zķ�QH E���Q�� i~56+�,�A�+�!�;���+�]ٓ#��_�����vKO7���i�P�����k�<�����,6�o�¥����B�Ög��~�qab7�/�9��-�F%���[��F��@�fF���7)/�ڧ�~W��R�e��&� ��U��b3�b����v�)_T3�g>�������L%`����2�$r��:.E���cs�m��OA�ȿE6z}0�Fm�qqpL\<R�`���f���ĕ;��!�u({�9Q�gD*�"������<�z��g�D�]Os�=�*s��;��c����]D���؈�u�Ӡ쓡ؕ
+m�����:0�ٷ��:���%C�����[�a�A���Դ���G�LMڙc�{��=%J������4����_N}�M(y"�-�d׳՛|~&r�P2������' q��^JMH�e2� ��|�Z��gov�HM��2�^#k\�xZ�������hY$�2vă4�O��+܌>n�E���g�����>�,��'����P�$D�K&�1���?s2�eV"}�Hk\n���'�v��0��k�t��?�'��yt��Z��ҙq�!in~��Q�e-��2�I9^�-���{iR�X�S��6{��^�+���9�8�2y�Pi�E����0Y��k��s�Z/��<�����^%�`xҷ���
��5u�`".B<&���h�o���,�8�xϻ" �� K<"n��/P��Z�e�.��۽���X����~٪�@�F��$eGˈ�2j���0��}����������A6�[�9�kB#|�R�����\n���ASJ�UQ�u<D'�.����|�)=�d�K7�V��>���ڥ��L}Yw|��(��@H}�'<wۖ� �F(����e+G'���ϸ˨h�ZEO��������`"��7�,�W��,ު@8w�>E��ϐKj���	H�<��9$净?%����؍�Ds��SpI4i� vE���؉!�Uj2C�JSB��m{���ȸ�[o��v4Y���?V��{�ڑ�x���Bt���(��E��*:�+�R�.I�=��G�s�&�7V���r���J�� @�<[f�'Ƞ�E�{q�~�?��a��G��DF�W��6�{�Q�����ϿS�H�d�,g���i�G������^��Dny<j~����q���$�kn��Y�O�OC��N���S�e8�ִ�����u���{T��ip-�����;�����b��yAi]��L�~��@����{�I�����%��7��aa�͍'�7��YG����#��	��WC�N_�x�w$���R��m'��:�_���[����f�+�Q?��?�b��%�<����j��gK4�[�4tբ��+���}O��X����4�u���	��SM'E�Nrv�5��#��"�e�Ё�qM�-�؋�^+�K��R:�	��aj�歨T~y�`@��C���{L��0,�3�	���e�4tKm���x����32���C�I���.DV����*B�J��*N�&H%��t���7)}ٖ��?�;9IJV7kG���j"��""�MC|pGnŮ.��_QFG?NLѨ���cU6�R�(�ϳ˺?���\t��՝q�'�.���&��$1#h�_z��I:�k��Y���U�|1��\��c4P�|��ǯµ�ɪ�����H���}������M��1v6��ֲ�·��/9�f�錥a�:S���b���{�����*�T��_��>I��㽻 wo ��⍍�P��45������g#]��
Z�y��S�� .��.:��I�o�_@�&Y뿝����s�E?֌��?�����7�@��4
.1��#��?���'�p�𘆿U9������W�฿�kl'�q���r?l\�.88;�i�����X(L&Nđs���#i��5��$5|3�b��~���tãp�K�|Cu�q�5%M!�O�Q- =�At�/��؊�M0u�P���gЉ8����:�>{g�fP�yΗ9��ܦ</����ړ!�Yf$�(/x��-����Pl�M�,ɨ���8�o���*[�b����A��G��w��ǌ\�9^Ye�~�ߧ<��4��p� �!�q�pI[f��[�����qF�N�oֵ3�C�iv�Q�If���}��_x��H���!<�ł?2qԢv��Z\2gzhC-�щ�`HE�4\N�6	�g�b�-0�dEo�?��%�������	Y�x�¢[v�24�i`]��"�Zޣ�)��B�Ud�Mu�E�����ɤk=���7v|Ջ�*j�!))z5dv���9ă��,k��Ial�)I��n���ǰ��]̚�&�x1$HS��$�P$����.���#=���SCTQC3M;D�b�Q_�1i\rȮ�*���8i�hH� �ɞ��Z����q[�A�l��@b�V���Thj/��̪��De��Y8>��Fz,3WVY#w=��	�8$j�.���8�UA7̭�u�s����^���Ħ�4�����[}"�栢������Tă�s�ߢ��A�e\�HP`�d�W��S�b�Պ	�ZG��2���#�3_$��m�)�����?-7è蛲���o<�2�}�� 1-dmU�����M�g�ce�����[\�i���lB�yM�H���K3��)��{7yز�t^Θ�Y t�*�s��0�wr1�p^ULp�/H c��[ۍ!��"���p^2�#wv�=�������֒J|�����:��g��SO�&�j�uy��zSp��A����uǐ��ʍ&�.�>qP��)Ni���>'����U�ݯu�YY(eGV�Ӏ{�tu��p�"Δ~�Y�jK�Ȫ�EI�l#st+�R�5�'.<�(mT����4~�@��-��z͐�ؑ+�o-��Ϻ �)�8LE�KV��v�ʦN��1Ո�3���𵁚�$��cw U��L�;�Ǚ&5�Y���V'� ��Y�]r��^|ϓ��]$�mq��}1�㮦�9��/#���"N�#?>_�=b��L|��H~��w6�S�vf&}i�Mtq�P��+�;�l��d!����	X�a��/
Ֆ��V����Xq���s;~�����z�&���W���P���P f�픢��DV[]U�;���$�0�+SV�[��T5_��_�F<��ep���Rο�Y�I��+�ٓh�!�mdQ9i��[&�oc���* F&���!�P���5�� WP����m-���J����%������+�²�H��%:��m����f�9g��"�.�0���G���CZ.έg���&�*�v��:3��b���w���zn�>�ӷc"G��p��m㹔����]����H�Td�IN��n�Baܫ��ȏB$מ�P`��]� Ձ��x��V�5Xym�M�	�eT�������������o������d&��FA����� ���T����/��Mhl+ѵ:�T?uյ��]�%���~�LoðF��aYj�\b�൅�p�Oy!a��_�[���K �غb?�����S_V[�g����y՛�P8�{W�V����"@ l���a�ȓ\ ��tm��}����<�TH�<��������U6��A�D�2��r���P�FRE���5Fu%�z�f5M�>��eLi"������X�չ�EUi}/C�Bר��Ⱍ�(�D�(�j�U�Im�t?ݒ�y����h����d��M���w�o�Ce�݂c|k�f���"�5z�Ik��d�r)|���$7�6s���b\�ԃ�PA*�&%��ǀ�3X`�[����܉.H���J�O��i���{�d���Xm�{����1�m���B��<��`:͊�
�T��C3�ř/p����:իυ���A&�
����wN�\�T��2���FUQ�?�),&����3�ȣK[K�y%�������#�E��=��n'fݎa0;"	���Th_CK��FA����ɲADPd�4��s{Ra�A=��fU�X{���_X��TI���=0�o(g���K�V�,���g�l�����l<_����/�>vO�M�d���L�Y��v���of`�y�"0k61�{�R�w����@��S�å�� N)���Fw��r֮g�M5dF9x����Fh���\q���( ���ދ])վ0�*B�0�� &b�`$]Q��J��t���'�-9�퍎$�Ιu�	30���߸��^#EF��ס�@_x�%(F�C:���y?<�LŮ�~aT0r�p0���8&pG�f5�<!��cv:��P��g��Q�%�J�[����Ӻ�C�48��H��|�#���б�h84�&�����EA��� �d1 ~}IJ\�\�y=�a����8��쾔��}W�-�]��P��z��T����l1��b5��r��e5D�(*4*�0'��[�8/�1ǩ׵��J<�XH��讚&�&u޵��%(�W:d�x���B������z�l�|�A"���
�*x��J��L}���7�x+{���/����0a �bC�gJ����~Ե�K�����s����W{�î�BW��a�
~n�{��y۵��m�6��靶�tPJ��l��G��s@F����j��ݵ#��R$۲�ڻE],�nO���^:aEhk���_֤��)��Z��I��2lk��-�1v5���"�������i5/�tG�1��B�Ijл�r��F`C�װ����>��*$N��aZ����=ٳ�$���zosY.���]��%������+�ONY��$9�H2bb�/�{)� (�݆�B$5g����{��^c5.�7%���D@FY��VJ�NƵ�\����jSw�ԒgU�� F�#i	3ʔ��O�+��7��-��7� ��!�KK*4V���( �x?�jT��B�IA���`�ܮcvO�VLb.� Dl��U3c���Etk	�������d��_UuEI5|b4�f����7���~o�|N/�}�� q��U[��HS	���1B6��/�ͧo�_]���R�/�dS���S�v �a6�ϻ�GQN�i&t�Y,_6�3-�<*R6z1P�9�-��k�����f�(���m��fϘ?~��Q�~��/�����;OKv�M�������@����qƓ_��FM)���oq� �k�qZ"������]��� Y:%�+�N���NG�=HeNŪXy��ѐ[0H�<��V�.(��\X(��6�Z�tBH�z��I<F�f�J[�Ce&xv�sO}�R�V�I��Z����W��ĆY���L+CLym��l$��Xjkc��^y��W�h�GH!j�^b�R3TB�������I��9pd��w�J�<fc�o��xif���xv5�-�vG�
��X�ia
Q��Uq��y�ۡ8����� �N0��
���B<���E���h����Jn��i<h�9ǟ���cTE�g�x[﷎2��u��y+��7�B�*�8��jEƥ�sk�K��+�H~���zx��'��S��)����Z	4i}�@EK�B���@��G@�0Ιba�{!�$6Q��֙�I�ݓ3��������V��Ɇ��ay�
����j�JE������N�0|���Z�b��kNZ��ff���/�p�<Hc���vq,�.�2gL� G���f��Y � �����x�)yQL�o0x�[�i�sP�;���J�-��ȯ$��\h���Q9��j���@�^uV�rY��f���Fzk�52%�a�}����WH5�(���������jzQ�'W'��Fq3~&~�7��@�(�3�q�ej� r?Y0�T�'X�=',hf0Y,<����$�z�ZN��
�ݛf�\�S�Nsp��>��@�K�U��;���V�w��rOQE��>��㺴��F�����ۡ1�ò�X��;1a���R��:Y!�2cz	��ᝳ���U�h�\��Э"K96�����Mn���~�u#�w�|�x5��LRy��pE���)f��(��b"Ζ���/�t�ߠ1:��Ђ�C˲��N1�u5r~�[EB�����1���-��1�fw|�T�yd�f��X�@a���G)ʊ�Y	ٮ�H��jAzk؈�m�L[|b٨>,��/ {�Z��\�kI�!	��D`�����	�e�?Vф{Ӷ'�o��>n���W��!���nl��I�w�Tƌn��^���R���X3uՏ-1פz�!Dkö|�-�c�A��D�z;�<'�׋r`�j	�#e�A��?�T$ܴ~ؕ�JoI��B*�	��M`O��Ǯ�\�4x��C+��S��]Tn� >�S��HP!	T�+�!	�^����m�|�r��ة����I崞=�%q��u�D�̈́���R�p�M��@��"<��v��Fh*%P��M/\�'�	D����bI�Z�
��Ta�w���>���cx�� H? ��G��s�uk/��C`�!�j1z�!���x^M�D�q$�'���ԕĺ��ܷFZm���xR��?+NO8�}jTT��v<�*��@
6D�?Jt�B�cvb�!Gi<l�.����7��z�^����9QWeA�!���b �Y�l�MI����īV�5Q(�a���C��Tsi����ܷ��$�!�!tv�:![)OC�b�@Fox3��]��#Ő�w�<_�'F���dm_J�����s_��**{��,[=ܚ��uͬ�Y����dA��@Ƚְ
*O�P%��^�A;q��e�!�+���at��i��vEsW�L�o��Y��4i����+Qy�������(�����㟚;�x���r�W�
���ݑ�V�8x� �i(��u�Ƨ�Z�V'�-XY:aV|���TͮR���O	����JZ�4�Đ};
�3}������u���]���c���Y��e(�ʈK��	��eK�s�h~�"�B*������{9���|�'�����*�	�,��M�;gxT��%͹M�K8�i��	���s=;qq��[�@O��(Y�̺�Ь�Fh�Z�|�5��Z��D�D̨�B|�*@$	{_֐���%�ջ�<@#�� ��E��vi=�7�D1���Z�O�]u��r���gY����Z��j68	��U��!��WT����)���0�6+Tq=���LvDu@�i����k:���2PvI�]�R|�K��&��(��0h������|t�$���G;4Z�a��?�+`4w�H=V0�te(���:n5�ګH��1�%y�{��a��7�aa���3�)wD��.s̖��W���LJP����0��^��HA�H>��k�m�%�o��G���ؤs��B��=�4�cf����>i�WfC���u|{�?(ڽ���B�E콋|�Cxu���Lmc�oP�m&GT���\����1k��g�Q�n �� ��Rsnc<S�<�Cڧ��LO^���۹kã�5*H����0�Ĩ��/�x �M�L�"'9�_������!���C+J��$��S8�gY��	�J�*�6�EZ`JA���ǥ�y3}D������I>���Z���yC�RMT��@�N(�h����C$�$'�o�3yҳ1V�ǿE���
���ȶ䘾k��T�[v�%+xpoo$�}�bz�D�-�xc�����w+�t"8$1�>~F�M�|=j�ޑ�{wY�����Y���5��H�KV�w)�1�� ���R���ά)�ESh �|ND��bUs��lP1�V�ڜ�r&�	�ٹ=�y.�͐�T�*M��-&�ԙ��< 5a�⤗�j3�t�.�]� ��Yi:��K��<I�h��P�b�:���dk���G��eB�Vݰ�醶�m,	F����u��@ ���d�����J�e�@���z��>Mi׫dv����@����S��/ܷB)|arX�=z���t�T����30g�~.�W��&feO��ċ}6bf��U=�w�n��Y�@7
��w+�g�|�ĭ.�o�������;�m3�����]����V:nx3+V��ߎ�ڙ��Y�e��%�k;��O�A���-���#R�᭶�0OVĳ/ͼ1U$o�kU��&W�3������}��h�\�����!��M8�Y�<�pH�'<6=4̄�rf2Μ%p���'f
v�Gb�b��G�d����`�x��߸��p���b��%=�<�[�e����ju!��v+��g;�7�EX��
Ar��nڽ�TJ��U�hƄ[�c���0E�a�W�`�����/��IΤ���?�z���M�(=�Ƹ�p��+�`�����|ۓ�2Q��'k�K}�5�W#b9yE'<�%8�J7�0/>���vJ��qLs��Y�_������f�صĸx�qS��a�D<��_y�)f.���r�ɮpb޾��{#��;�[j{da�/:\Iq7��j�(?M�pޠ�0~;��E��k�0���	#��`�ˮS i�Ҏ(z��GY�c ����W+~�(X�Co�C^~�b�����A���Q���g/��[K�nb��G3&m8�3�'��(`X<0{�%x��.6LF����pv�C�A�q���z���߬�%�/s=$kȭ(�8�5�ڔ�?�p�^+�L}�\�����9Fgc��P�@3���7d����E{J��3����mL��s��||��8+�����iS��!��G��>|�����j��=�;u+j{�9D�4=/�t\+��z�xo<�{�o|��=�v�2p3%X�r�5E�-��#/y]�A�
�pcp @�}�P�1�;�9$*��y�t�#@�*���C(V�Ŏ]�ٟDb2��3�ѐ:�-�b��[��3l�����S�	@u	Y�Ǉ��>�n�c����u7����d*�(���Ţ��K;��aU�}��z��K�;jv�A����Y1�p������׃�`.�:�gaB�n����"NC��Ded�=�ݮ|Ʃ����w=��}+R!�������܁'�Y�g@]l����>�D��H���R�W2�\��V��]οl	�6�ҟ&$����g�φ#��+����r���(n����:���O dNe���b�_�e�����hw���R�"���)�F
b ���/��d=-��w�3�vzP�'����Q(�v#��C�o{����~��a[��0<  Zc�i�z���zV�2���Z���=�=�bum�s�jQk�<�7``��PS#}?����r[����\q�t���@gL-�o��M�w�ee�ac�Ym���[��l�RC�N�nY �T�V�;�dA����$�� ���E���3C�2�s�38CHZ�Z�!����� ���p���ƽ�w�M4�w�^���k`2w]J�����k�����Z0A�~	�GF��{hM!�F6v#�-"ǭz�0���uB|����=Cc�Ēn�Isk���r,���9��$nfk�ՅN���1�>Ǹ��M ~&�s��~�Imv�tXgj���oeG�[M!
z�r+L���^�mz/��ǌnV����3a�>%���_�Nx,������ܵ�#K��K����J�U6)w>�|�K�h�X��t46�ab�n�0��QޛW���]:��BCi�$I.þ/�Y���<�
��F�@�oI�*M6\�����0a�$�C�W�ʆI���.�^�fs����c�w��
҉�c��(^��M�����
�#rlm�!�C�c�ʪƳҮ]�P+���鶷.�1,��l���]��3۠����YdH����:�G��� �0y��G�O�qڟ_]�Q��6�w�K�lQ7�I�f��>�7�BW�1�G�Qd��4���,F�*
j�)�R�f#Y2��7k�^8[�y�&N%RvBEt�i9QX��D!)��=���e@hq�)̝�N+:�|PEk+g�[Mhe�T��w�F�俍��eu1���s�;cs�"q��K�I$��I���[�&{E�aS!^$�"�K_ ��R�T�ݹ������Y}f��Ŕ��B�O-N�ԕ��3@�k��ug���#�c�P��|�U�.D*��#o�݄�IA�/Y��4��n��+�(=wC����ԑ���Y�^�T�:$O��R驤�n�i�!�U[��M�/���Kɪ7�� �P��c+��ڈ�-N�,�MB��؝�ﴴ\h��0)��凨� "�'n1'���FG��et��D	�ŋ�����6*�MR�2��毨4wi�K���?pND�R�7��>;��hu]˱�踜�|}Vϻ���y*��ku.�vŎ�0ǻa��������P�Q�����aPFj�`���_94��g�к�g��d> �7b�����$��I��Ŀ�h�=�w'�0|�KkPQ@o7��)D%��T/%"�jV�=\���X���yjbc�Kq�n���*����Ξ�l�^���w��V:*�}3�W��쁪���y��հ���`9؞x����ޥtB i�O$&(��G�v:X�:+�.�=\��3x�C��-�e��H�oοhgYe�)z���ґ\|�I!��ab����S�xK�>L9( �PV4�(џ�/��d�Q�-�&��~���#?�
h-���+��I
�Qdj��
�\�&ɔ5�%^�)X� �4���f�4wN�[Ρ00�&�けi���<|�F4�� �"���r����D�F������3�L�S^Qi�����G�/Cd��R4�T[����+v���|81��=�3���8���>���/��|F�5�{MM3��2��R���Tq#.����D�cިl��Q�g,�U�L�we��A�8�HB�B�֘<�>�B�´��)��7"�w�S�VmG[��P㕣ӐoO�7�X��jd"�p�,Y�$.}�j}��HR��mk8J���8�&�84ٮb"�lk|MI�������������_��*�Ѹ�P��6�~�.㗀]{ҕ�ll�O���/�63�sǲ�-��[hAr�\5"3��Kn��E. 2�7Yl��F��9H�{�=Q!J��ԸQ�m�b��{������(s�43�|���.�;�Fa��O
c�
�e�v�!���R�t�����k��0��<1�1-�S�?���f�n:,6k֔\χC���w=�;�2�T��p8�K��>�.@�����K�Mj�{ ��Pdl�6�m"�%��9*�:/Cqyq��w��#�ѯ.o7w�Jt��vڮk�S�V�A
&
uB��t.b��ū
��m�f
������E�M^l� �|I��N@魇�l�+w�_Uj<I͎nR���{k���ޥ1�ɮ) ��X��]�V�Lyϫ_1��EZVZ��W�@z�S��IDGR���m(%��(b���� ��x$gc�S�:Kb[�����v�+Sl��ݎ�������7��tܾ��+�����W���lMz�ʥҢ��BOLV_E�ŕ�y.����4R���]l��D�Ug��O���,�rt'���O^�7r��j3�J�����'I�I�e@̉�v���˛���&͊&��T��M�T��N.�a�xy:�����	Z�m%U(`�ɐ�gf�Yy�Hp.!�O"��ǀK;��B����W�kIk�He	����Pg7he���o��m���h����p����m�h5� ��~,����B��?ifb�v�3�ɡi$���iZdɜ�2�A_7�h�S�^�oV���}B&}-R��5��B����c�'���ra�5%-���]S�w38Oiᄏ�VK� ��Y	x�#A�ZND	k���(t8B�d��HT����E��R�2�=�u+��~~�w�yBB/{2�N��p |'��z�c���^�7��X�I�s�f�܅LE�O���ɮ�'Xpe9d�������	^��]&�T�ů	ٴ(>P�L��V�w�Fᴏ���x�Tªp�R�q^M�G�i���U����������Z]8F���y��yN�#+�	w�ɶ���yQ�i7F�*�T�����$�lL�X�����$�I�W���2D���g7�:�o{g�$M:Fx4�K	��.��A��3,�����cTm�R39.�	B�l��.��-It}��v�X�S�0<�[�5��AzK�Y�s����&���qd��U5��y6S��i��`�GE�D��k��aK�&e�)ke��&A��%Kap��4��&�)�cs[O�]=�1U�Ɠ<Q[���e�=�B�k����?���̆e��l;N>X �w�!:$�4�Ȭ��-!d� ����aH�L���%�׈j����p$Np�z��ﾕ|2�7�S��4�����:��Up��{<���.�D+��d�=����GF�,��`��4��#"<����k�ջ�`�!�"�η�qJ!r����o���9�6���E��d�;G'aGAT�qs��⭗aˊ2� ��!T3gS�$g�G*����)m��!��8"\����;Q��`�Aq�cj�s_�W����x	���$�����5�V�T�Yp�;r��~�߮'�4��j�X���gyq��Joa>%�(x5�R�p��~ Rn�<�4D]� 4���K��q����a�(K�,��;�&'����~��Ң�)�	��F;�9�(��D����KZAZ���"7��;Xs�㕐�@HV�Y��(��|�/]I���6�� ��Rf{C1���Q���v�U�!'Ѷ��+���N�F�a�Z�W9+�F�H��h��xq�>
-���q
�"��p3'�P[���#Jpi�d_�@>�l[J�u��V���!��s�?��+��j9:�} �����Z�RS��cS�@L�7:�c1^�a֚%.��w��*�9��@:�$�K�i�p������M�}�|��P���
�$2w�ٸi����3�H(	[��X
��nk8MJ-e p̻Qa�J�y�kge'�?H�y�l�����(]�]ڷ����M'u�y��K�C���o�)�^y1�;�A��nb�3�.�^�[��%c��䋞K�S��3�"�0�<۫��gS�
��L����=s�������.A���XU���;_6��������{�&���s0�YIy����QP��G!�&yuݓ�"��s���
�^��6%̀(�qЕbӃ������' �bHS[J|�m�� 7S�9���9!f��is��d%��׊�?���I��t�-8=���dxc!VbK�
��pd���X�|u�u�tG�u��4Z�u�o�t���O/M29���B��/�Kn�6��1h_��~��sr���޹����ď���9�j�Z����B��^.$ L_��]S"Ӌ�0Q���7�?.ي,(G��ώ'����2Xx���<cϼ�NFu@�1a=��0Ƃ�)�V$�8�7h�P:]iͧǐH�~�uZ)�U�}�w�N)��F�}�0�c���n��
� �Lٷl���xHQ���xx��=��_�K~�;�k5>�xt���Z��}ui�r�S�P.��&Z:g*�) r#�r�,f
Z��jW�[ɚ�l�Y��I�k.X�~�-�z+x�ܸ y��M�͵a��bD/qX�5�R���%�"wc�Th�	�}�%/��L.(1w��� �� B��>�Ӑ�A�w�y)����^�H�Zhy�:��� ����CT�A��K��u����+���Ҟݩ�L����Y[��=]�Ԓ�!�ǜ����n�
���G�=r��mD���i�.� ��ɭf������.	̆F[���ﺅ3�@p?�z}�R���H�k����+�\�(�>�֪m��؄n�٠� z�@������vt�Zͺ���J�`O�Gr6�I�Cb�/u��������N���7|xg�,i�!��k��P\<��U9ʷ�l�P/	��-��%�9�C�ja���*3�vxP���x�z�qh�z4&a���N �=�E�\�m�w��L(���2��������@�b�`��l�D`#��m�?i���]��>T@�(ꌊ��N�gw1���Ƌ��(�+�K@F��B���L�/5n�BM�H��l�������j�\�9h�To���@ӌ�[
�Z��7�:[R�o7�FrB��h�Ǳ��Q��c�����ƚ$!��Xj=�r4�_s 7�/��z���p���%!_�xc��c݃�N�_l"#=X�PR�_-�u�Y���FFs��ѧ���F�>?���l1�{��^�w��;�ä(NG��þnh�P�n��v�b�,H�l������&-V���&������)�C�N�"�hR6q!a~h�v����ˉ�J�ѥּ��3����W���*mf<����Q�,:]>��gN*]��k��%@��q4�v��%���W�i���sb�p�(�	@=H��DD8�/��M
�r�k��T8�*��H���c#*�m;#� ,�I�H�xsn'yup����wS�&�1x_c��sO�����\ߞQ��|��yx�V{NS%�
�y\�[=v�Ó��yW�2���pB�O��jB���Kjp.�zf����|P��J���z�%*�J�Cn7�yo���#�1�2���TY�66D �/�x��kf;%�W,�a˜�?=U��J��欉H�1����h�囂��?�I�h�z�z�h��;m}�3�(��� 8���Y���<]o
��I�C����q�5.X'������t/а�ɒͮn��+�$E�K/�x�-!��9�f|e�`,�aU꼜��FZ�2Q���Hv�U9��&��3ٳ�C~ݨ�k\]2����8��X�����Y�
�#�R�HQ4ìReگ�O�('@��rh���#˗f�.�(V�jCL@�Ok\,��]�w&��"�c}��8�G��dE�p�-c��p*��������-�׺z�9��w���]�[w�����C���I \P�+���iʹs�T3Bu��4��<�NO_!)���و���+��%��X�ŕ�8P�x�Iۍ�̈́���#b?��������?&�F����^Q���_E��m�pç��P�qT/�C�[MPL���b��e�M6��O�G�C��2�A��L9{��*�JƝ�_���$2�L0��E��"&p��a�R	�SOd�j�	�A�"�*;�!������?��6�����w�Z
�� �$<<j�̺�K��;|��Nm�w�}-��܄b>����Q��JI�����@x���ʔWE�� iLǾb�f�����tI�4$��Sm����<M�ab^�5��8��>���ݪ�ܧ��ݯp/L��:@�ڼ�y�pX󷧸�f�?��q��*��;LS�	Fx2��a�����q�r�s����ECǎ�?e��gźqƷ���& o�}�}39��L���{5��v ������ڙ`��:���[(�e]�>U7�'�r���W3m�Wڐ���P��s�"3�*iO|�����sĲ=/P���~��\]�9�[9�S6���T�	nI�)y ̘��<W���W�c^�J���T-]�5^4��g5@ǣ�)
;g�؝�DBO�h��h;�f���<<�5���&O+��!�!}[�5y�6d���U�)���2(��@�A7�)0N����]����U҈6�{�1c)*j�Drx����f���;f@��?����6�$�"��$��8�{tXB����.�BW�']%���@������N��]�uA24�b�4����2/��[�?�׍��$f��d)M�!#~�q�����C�H]I�'��ކ�=����73��9���B���ֱڦ.�=�%r=�Go�k/���j�F Җ��1#���,UT�����E�^~r �6 �B�t5���z
�;4����2�sצ����JG'��Ě����3Ϸ��d�D���?�D�BH���("���K個|+���	�똚@Q�b���q([�Ж'������6�/�K���`�0δ+T��|
�0V
t��D��gG�9�,�˶�d7�ݎ���޶�T#I� �h%_;}#/JoK�����v�^\�іC����9����N�U���6Z��^�}j���s�#І�ч ��ZR:�ȝ����&�D�4�,m���D�J�e���a9i�����3><���ʆÆ��K�SK]�2��S�HOr]����2\�Tɂ�`L�ѵ.���+7�DnԞM�o�J��ccMif�L�}E��hQz�+�mLV�J69�ID��<��R5f��7�\J�o�FF|���J��5���f�\�˄B�Sv+�
�P����$�*�AU,���lT�}��OxG�W7e��uj3Ұ�2T�k�.�cv�	�[�!�3�)�G���ӐѠU�d�&N�/�3�,MS(ট�
C�F�-��nad�FI�:e$�M�v�e��"?�[n�޽t�\�X�'�C��w�q�O�oIƢ�V�c>�����'95\��g^������7d���$����/%�����r��͗ ԩg�N��Z�������x�K�����6�&F����ߋ���h�	��]~O9�K�97�J�p��f�;3��^���A�)��ޡSƣ���o�B?�{R�M�T�z��XN��M(���0*m�9|�8U�v��H��|B"e5�����o�ђ~^����庮�6�`���e-�o��ɍO���v~O��[�l�N��N&I��,b%Ӑdۓ������g?�8nQ�x�e	���4��ϺfQv��L:1�i���l��&��t��l�W���#e��% >�4Ȯ@��ʫA]��#�F,�ϧ�d�d���vj5��ᆾ�@1�j��1���As31b�c�Sٓ�D-���¶����-�U<=L�x!�{M=j�&�+�0,��c`y�k�hXt�ZX���1h�u�%��MD�.40�L�7X���B�䪖Gq��=���.�i�M�{D�_��güi�v���x#V�ǘ���ս `�,<ҭ��صԇt-�����9!����1�;�gK��Uա����Q� Z��Q(�Z��7�}����뾏�0H>l����&e���*dyB���F�C�5p�YKMB�;�#�h�
�fQ	jr��4-8VN|�3w$C���;�w�SJ��V��Q� C&�����D�fh!�p����6��$b�B���>�i&Ϥ���[ĭ��t��@�[/ņ>�<D�_�͈��5^:�a��0��^���;���gh�83����r3-q/Y�s�g{��+ 8&Cx���ٷ�u��H�.�LW�_�y3��ꖧL�����d>ſ8��.�S�TfN�,O�%����®�i������\Ԋr��2ׅ�X��T���rl�&�D�C���9{�R{7�J�ȡ�����{��#n]�Mi�ꕶ�l(8�WU	5Uc�D娥����U��1�z�f��K��@�چS�_I���&S��S���f=��`N���K��z�Tn�߰G_�K4�g��>���`�;e�0U�Cf�'	vƛ�>rd	I�"�V8�5R�xV�c���l6})'���J��ސ6x�$Aa��
�u��F%mq%@1�[rC@��e�am���<�\[Q�7��U)�}"�j;���$�K�����k�򼈻�����JX�ڔ1��(��K�fs��_�Ш�ˡ�a�϶�M(-%Cu����
��x���ܬ2��WG�����F���_`���Y�4�	r�Q/��bDm፦�E��C��VHԧ����d0�DR�k�}�`F�*� �W34���Kt%�h��o�q3�8C�(�tyc_#魇�&9�П�n����x�4��Jmv��E�O�\��:�G����I�w�I������dU�/��Tt"�`�g�P��C���\BE���<�s�A�똥:���޺��(u����/_�g��u�=���m��y�_�U�HE8{ A��_<�F���ÿˊV8Vo����SN��($��5��پE�\��	eo2�}�侬Q�;��R��a�g,�Az?���{K�G?�'w_�XG�jk��>5���e����p��F��Yr"����#�.ٙp�n_5��FR2���j�(���>.��5�zAAI�⦤Т�\q�A��tYM�{Ӿt�?Y�\<A\a;�o7�Ǥ����{��� "|sI'�8�l���>�jAG\��*����z�z���s��h�	�3z���ؐ�y{��}��|�mϱ�[����S?-MN0 �Y����8E�+r�;�4T]��5G��u�< ��,�i��5�u�IU��c��*�f����@�0�ЫUp$G/L
����0����CO8~`��W#�(}�dȏ7{�Ǒ$�L�h	�ir~����V�!��
k��W�������v��0q({�׆�Fї"�=۬o,�c��v^@���O06�&WA�jLP�} BY�+�A�Q�%�}Z�w�:5*b��e���r��*��]�����|���L��U�!�E/�%
�}D�Q�qu��=������,%�\�P#�	��jxëE;�� �y��BK޾�8gKT�µ&}K��ɿ�����؆���ݲ�{��.�nhQL*:���M؎���c6E�2O�R*��nNB�bY����f�����W��#�o+Ж��פţp�֗���Ag �l�m�FJAY��W��K�?����5�@�����Q
�����l�P<1��(Ѧ�k�E����A�8�D�>�Ui�F�Xv8b���C�5��s�)YH���Ŧ��| �E��������j����v�_�	×m�.Qh$��W��WL�z��-��IYaJ���c3n�r>�7�2����Bvn˒�l~���kԧ����G6�$�������(��{��� 0�_!*c���vn^�,��_:�4Mv�pE�f�RWs!"���OEY�0�������[������8-J�:g�×��e�jq�A��j��.��:�q��Q|gZ��X����)[`��so��i�bF��#滀w���MLHKr����zm��~�/��`.i/���tU3x2�eB�`ؒ�;!9f^k�:��_d� ��,��'cQr��K�\<��I�d+�Y����ڛu�t���cH�=�ؠe����@'��.0x���|�_��~	m ��2��n����:���B��H8-�[���JgX���=�0��'՝"��*O�8�"c�����K�"S	���Z^���FkZ�{��w{�A*�_D%�DY'�1b��4��4^W<�.��ݟ��hZ�ȋp4^y�>�2ƆS���̆�i�sB`L�����pA.Z��*\1�?���֟�
Y�-C	4$�