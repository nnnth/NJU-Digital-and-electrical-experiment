��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�E3�hoA�zFҿT毅���M�"�w�g��޷Q_��E��.N�^��� �Oz�=>Yj�-�({_@n�� O|y2��9���/��a�o@�l��{���X"�������G-�Z�VI��#��Sy�_b����hwŉ�8���\���bR}t��a\I�l���

�(I��(�O�C���w�ߋ�7�1#��,K�ʲ ԩ!��~��ܢ�?鍤���I�SՊ]� �x� _�,��0�u����G�n��H�����v�i�N�gm�{h2��h��޴C��T|��;k�Xj��_OEvƬ�Q2Nπ�q����6����@IC�@oŋj3#N+�$���S3u|�y�"%�	��Z���B��|Of�úli���76��2$�j��8艣�Wz#'a�Y��{"�)&}����F￿�V9�|��4�q���&P%`�:x �9�?g�y��`;R��H��t�e .%�e�@�2Y� N��+�U��b������Pc�'%/a�蔛�)]@;&xn&@�����(#9�@�7�$ 	(P�k{
�2L�$��AI��	F�AZTG��*jMb�5N��^e_1�����h���X�'��Ηk2��
���j�D,p��"�p�^���B�"��!�����?uu71�fZwD֓З�a(o��},;�6��T^�C�<_��~��y��_={��N,�l��~5�f�8w�����7��},�H���$�M2������ȗ1
9.oq�d��#ns��������(;�d&f��H]S�1V��ַ6�!�$��,�l�B2�Ss��]|�n�)�:{��3c����J	��	n�-4z�1���N@�X�W�/:����)���t�E�L/5>D����%�بͷ\u��o6�"[��-ʉ����IaD��]�c��E��I�c�Z�g� IN�r�G�MG�6�@�����*u��z�!sM�V�`l)Z�����z��?�)���Az%z���k�Bp<�۟%� �'�+���Zo� �A?p�JN���m�ո��J`J-���T;�2���?հ��3��.^�Ht�<��&G�9���Լ������yw+�eU�i�[M�����C��9^d&~��٬�_g��O]�ee�뀂~k�ǅ��u6Nc:S�]Ш��	a͖���fI�ڂF���d%uf��Ko��d���|�j'ӽ f����<O���S{�N�'#~ֲ���� ���!څy%�e~�I����ɹ=�J
�H5E69d�Cv�{��������r|{b��Q���}Y��ݔ۔O�����E�x�V�a�T�3��.
�9�u����Ðo-7�M�|���<"�XfT�^� ���Pٮ����$�IҌ��ζ �3���?�/�d7���L�S$�3;��b�=��1Dt�!�6b㸐.1rd��_��t�LP�m��*���c���0AN0}5[�_��d���TB�b�-���G�ݩ^�:�1����Ľ�amL;y_N�B�0౽�%���h7�������匘����O͛R�&/��1U|5L�-H�vS�ceJ���`�l�ɴ#�<�ibm�<i��ʸ�<9��beI/	�AF6��lW�5k��:���tQOmf"o`�7Ns�� ��dk��j�~�?�Qi%Y�]�����V 惉�Z7lu��ي!w?����@�Գ�dr4��s��R��d:	+PLu�������}�;����!κ{��[_��≮��Ti-W�b��o �T��.q�0��*�r�B~�r�#��u����Q�^�!\�ֹA�[sҿ*�(��e��z"�FB�.��F�{62ҪJ�'_���GTݣdU��/w.u��xH/~�0����$�j�0Zl{2���
�/6�ꕯ�y�����m���}���tv8l�gz�1�������0�&�K�L�Ų��Aa�Uuݚ��*��n�F�E!�����  �ᇙM1;B�f"3�7�'�,�g�ں�f$�?g��G��/
%W����f�?#����p�<g�ס�Cy�LBϫ�u�� �/Ӊ=Q���?Xyvߘo}�d��Ӗ�	ez��g��dj�,eB���A�%]����:����oeJ�)r2��*�0���q���Ǐ!�ˤVd��3��ԩvl M�= �l�C	��ʹ�9;��<��8�(�X�!yb�N��=��C����А{���׼�G�Z��M{�O�W`�y������������&�R20��=��K���򢼗��Z=�Ʒ�>�kG�鈑_��\�D����y����|1K~��"��x�ϲ�tl�îpH�L�l�)h�L	O�b1�$v��Np�I�$�G�M�\)���F�����@d�� �j��R�5�Dy�\n��s��Tc���J���a��8-�Z�ѫX��&	�z�?,��׵t�k���'��R��{�T��2�4��2�zz[�3�1e��Rs�QB�Z�bR�0z�?_�����<��r#�.?L��.��v�����%m��19�F}���,����Z�7�#-�
��ϾD.(�4�N2�1���:�
p�05���:~JD���U��UXf��w�A4h���D�̗k?4�T���u��NOu~0	\��1m!�;��%nt����J�zOs�q��T�^�7B�*��E�|�h�'���[�+T�~�f���\�;�"��wi��.^]ΕX��^���F�%\�-��ڣ�	S�!�X�_ڬ/r�}���P@����2���G�f� J��FF#�P3��<��{�DZ�?��ʌ�p$	[T����nU?���=���]���w�
z�3d̹�ܭ��>H�,d�s~SL���k���e�i�t���;_0�}�Q��O�����52����X��Q�kZ{"�o�Ӱc�v��� ���4q<ƾE��2K��<�u,÷�\­��+��MV2ʘ���[����E��Q�>fX8[&��^0���Bpn��0��L^xGw�}�R{xi�Uu���g�CL��<F�7Y����.�A0Mjw��0���b�`���S��r�s0�-���Z�ў$�G� w&5�*h��a�׌@�I6���i�VpI�!���z�V�2��.Ă�W��/���(��9��!�C*"��i?��`�H
��%��/��.E��}�>�鴪�+~��'�^4�g�O������A�0��[��Kkp�M�{菤8�<F���Cw�-�p.�8�S�ςEY�.�g���
p�)u9d�}��L���RF���q���i����f�_.��`��-�ˈ޵��k���d�
����ƀ�D8s{�X��U�3��y�ܼ丑�E}�n���Ǐ,�V��ʬL	*�V;(|q#���z�?�����I^���T�� Z����b2������C���%�$���8/���#��$�a�ե�?:�i�r�|�@\@��B�$U����DVV�?������h�.��i_�Z�)�ڗ;n?yc������zeo>�z_ؽ�,_�ٵ`�}�7�8�d��d0�N��9�b�8�A�)��P��&�O5=�R�7Y���|{���ڋ槰�r�*0=��3��G\���&���*ޞ"�Mj��G/8T�������.�%�L,��/�z$6r����� �$�"�Nj��;}���(�����J�Ϥ۶{tC���#�_*wd�[�^�#o!Sm�21v�-%:m^P�Wi�>�b/ON�5�=�T�0�=g5�*_�������(�a�w�r�C� ��S��c�9��K#�*~�R��u�Eu.�6�sЁ'+�4���t��A�U�7=b/�~#�Q�K��` �e�z!�n,�C[�əb�z�J"�����KY?#	盖و�V��Z�c�Ps�X��^y�2	���^�*�k8����PCC�l6
�	�s�|z��F
-Lxeg����W��Q�7I���hҷ�*v�xV3�P�\`5�sI�&�T�D9�rŒ5������� [Kn',��+JY�E��GΩC[Ϗ��=M����3O��jc�WN�/�[�X?�����j�(����B!�;r��{mZ�zx&,K<�y� ڝ�����z~�,���#Tizρ���>�0c��4�vb���z�?� �7M��^=�>R��`���FQp������i�m��W^�	�M�6�ꌤ�>�>��-�ZŢ�j� ��bmZ��:~K�8'��A̻Y]������U�?K�Ȓb�~;��m����"{��`M����n"86G���PDQ��ޗ��egN��>L�����r�J�A����D�x ��p��I�z�&�J�e����^��$߶ִ~��bC I\��W#}�n�w<�Kx"v5���N[�����xYLY$*��Kd,+�IP���5��9k�j��� 2�3x(&uc�'��'W�;�[,I�=�����;��n6�1l9�:%�}��}�r����a:ݟ�$l�~�Y�h���S�+ͩ
2D{ԝ����`$��mjڌx �Ǔ/w[��V���M��T/�q�'M���&���i���y�2���o?`����[�z���aC@ ��1��x�s}z�����E��,{��.�(��8ګ�=]��bK8��aN���,�_�� }Z;�]eI���]&ccf��tp�@u5�$C�OΝt�6�C��**(�!�c�mH_�1۝�XV�Sԅ�U�ۋ	H�>\��Y<�t�7I_([Mj۷	���	���}\e	L�`F�M�yQR���fܤ��#���
��}�tW���X�Ԃ$W�#w�٠a�8� ^_��9��K��t)9�R�������Žr�Eg"�D��M�[_J��M�T	��Ge {�ʝ�BgC��j��M1�q]#"aC7H1 �%���ୋqU�2���koނ�#�r��\�{�[�==�ǻ�c,�@�XI��rK�r�g�hй���a��77��<�6/�(�A�#�1
eY��d�j|շ�	;�D�rX�H۽ۈ���_�("����;���WI����K�������`39����>Ot
y�9Eݵ�G:�������i��Y!UW�!-jt��̇����Y�)qߚ�&>�WzQ�\�6�hX�U'�BF��g�z��B�W�����']"�����\�	����<ek$S�R�cO���e�������m�)��qjl �M���-�'�!�(�4�?0:IUEt<��^N��֗ݠ(jL/�F%���s%�Q�g�����\~��0}�v��L�����/���XH�tѓ�����<�����ܝ)l���P�Fk5���c5A'��f<i����d^zw�Kw��U��@�u�r\7�TԹ��Ԫ�9��4�c�|^i�ӕ�5��yػ@ёϢ�2vmR�Wg�D�䞰
����L���P���������~�r��*�`��_Jgr�8� �<�������UٓգU�`��ܶ�Bч���m�X�A��R'�I�潑��I�Xw��'��b1�dm���J#�<WK"j8�M�/���Խ6��pD~��Η��;)�|���^��v������͠3�<����_��r�۸ت�\Y��ϑ�n!ϵ��dD��^�*�~�c�n�!7�kb����?��2�V�T�⻇t`��7��v����]��'����E�DL_�O`1p�q�1��:�)��8cQ�w�2�4�l]�!=c|&\��)�IH'g��D�y�oE�:��6��������h�fTh��Ɛ`
�lQ8PK8��N[g��d�{{dϺ[3Ԓƍ�j�PF���y���	���� �[����r����c�kc�%��ix^#�R[��6y��d_�K�{������8�g>�����'T8� ��l,/�(Vǉ��uL�JjEYq���&��{�.�m��KM�t�V=��:oz�>���$�9Q�8�-+z�YD��q�g5��M�s�����\t0�����s�(�9���c4��vM:�2�Vg�0�;8�P'�X�p��eC���Ш⌠�%�w֦R@E�k�ӱ��s�^���ȹ��,��h��9D���Mj��� �]-�1x��ed��̌�Fˀ�"9��Y�70��kZj��F44��	f����n�ǰ]�5�Mf��(�"Vҡ6�(�d�5� R�>Kn�eM�ǎ2��[ի�����։�:�c���5y~\$/�	��\��b6Ҭ����L�`�ء���H�~a��_o��=��}��n����6�0����㓗o�g"��GS)(� `+�}4��KAJ���_��s��ۛ�|���a��FE���En�\�P*+<�fO��(���HA�	��nפ2.g�������=ؚ%))5v7�)��H�d
�ў5h��c���b�ᣢІu������-I�ʥ�}�s��\���ir �5ɋ "�9���*#ks3T�o4�qW�1�!T��u��5�do�v�:m�Ke�z�a�(H�H�'����큵L:���UrzI�H�g��?ĘO���	Y[�S���a�c��#��Q�y8�n@�o���nP)V�a�����^�O.v��A۝=�/a	�sމm��CvS�I����~j����F��5x�
˦�tD���r�F�^kҞ�>��Xy1L�)`�8JR�k'��v�s$q��]��.$"�S�h��S�9�2T�z�0$<��ׯ�4�!��0�"������D�%n�,��J�֢�羴C�W�x,��o�I �! �X��_y�&\V�~v�X��t\%C&>��W�m�㘂�g5N#�9����VG8�B� �teY�:���tٞ�A��g����,<��a+�/=����ݼ��R����$hHcUb�o��a̖��]�C���l��EΡv-�sڲ���3D4�AJ_�78�J3&-U%|5��#�i��$yw�H L6���!�oV�$L��!՟4�\B ���}h����u�f]��8g�!A�{��qfΚ1*փsC�k|
J��w�&5}��c�h��/�擞�B(�>�`0��84G^��/m���*̴Ś?d�0�7�W;� � R��m%��u0�O⢌�����/V���?oޤh�����IE&<tީ�@\>��:i-	�As~��?��]��K�qw�z$a�����D��N�.ﶴw��V~�2ŕ�X+!�����a ��{�B'���]�r��"����Tyt �2>V��z�M������)[��2}�=%"�ATI���t:{9ͭ�w6�d Q���I�����b1�j�JOrr6L42��J\TTv.\�ǹΙY�
����5\���P����zq���	$�w�p��}<H&��<��>&�{�JN�A��w�GD"�HeN|�+)�x.߫���:�"C�X��ш?tPA�ک}��5PHEd�S+M�h1$M�W liŢ�^����T��J��vE��CW��ٳ���f�=���?�ز�2#ӱ�����/:�=X���>vdd�O��ʡ7Q��I�R8���a��,�u-n� n���Z��(yc�M{)��]�P'����͂ƾ�|T�5�J�I`F��ȸԿ	�T"�0�FZ������"��0���}��uȳ`�0�ޕm�\��&�����@BJ/���ӏ�,����d�`��~m���JT��x0N#]]��Qj��,,-u�R�-x�f&�w:��H苿�<Gs��R��7�Pڠ�]��2��~i`���?�aT������o�c�i'yE���O ���+5�V��Ukk^	�Q:��n �i�HI*��w?�E���m�k��SCէب�q��n�)�����{�t;���}kބ\u�.YUh<�/�
�C� A�5�)4J������Ф�N���s&NCz��(&D_�8��/R���QO�
Dl�������*l��:�uw7�a�V!U���䂌8�h��*����dy��d�E{�x ���^�=� <P`I�|���
�����gh�i�^-�,�AIz��s�)w.c8E)�(�!N���N��P�ph��`���?���m���2��i;\�'5���ݵ����~g.��2�,K/�G�Ci� 
�j�U0)#q�W�V�f��;�tG��8�5ظ��U`��l0ޱ�N��eɻ\����J�g��Ǜ��`m��=����z���j&���k�� ����}�4Di��cU�5 �'�\eS[6�Q�Go�	.�}����#�����bY�\�m�ٓ�ˤ�:�ou�P���݌MM.��H��é{Ijb�%EA�t�$�csF�"2��'�����C�f�,�b�0o���^d|6�/e?��d��"{&��F�\C_Q���#��u9���w�j1��8�C���F����&8}�P���l��~u��f<K��M
v�tmn��n���D�-}��g%D���oK��,#�ޭZ�
9^;�SM.Ι^�e��sK�"^����Y��~��y�Y�+ �� ָ�4x|��K�'���w�)uj@�Q����9w���vx�0x���W��mZ#��S;承�����]�9go�1
z�+�U�[W,���_*"	��ξH���5����BQ9heҽ���aU{~���F�_�ð#K�����bB��
c��>������(?��L�����R}{�FS^v�Y��������ӎk�8��t��Is@�_l���Z��@�����ސ�^�� ho><�������\�Ĉ+Lz�Y���q��16N-�;Kԧ����I����[H��M&N������IU1�8��[Kr-���Em�?��)�}n�k�uB�Q~����A0U�}-T,V.�1�ߘ|��[٫�q�i֙�t���,S(�F}.�)$efY��#N<ɔ�m��7�W�����f���h,��b$��>�)ڄwo�䡗�B���?w3!�(��]�a�r�6�@m6�Jx�����L��,"��Zl.������װi�A�F��F�����:�l�[?taC����/69/#G�5cä���`�ćZJ��T\�v�}+��l�T�|!aG�)
gPX���l��<�I�Ӥ�鍝z}c���|�|G���EDn�mD3��L�}V�W- �v]����h��
����Frꂮ���i쪽�|�B"
X����b���~�[�bJy�9�Ѹ�LN��A��\�|7Ԏ��+�*%��oI|�o�%[֣ul\��a�˞�H��֗x��hg�K�>yI����ӣ���~H�c���n��5f۴�g�ӧ�?[}�E@���T��N����CԽ¡a499p�"��Q�c�Z	�#r d? �c�����Ę���:�yΙ�T�-��|-�l�q���^�g�0�.����u�L���E�����2\Ww��ny�4	u�|����"�x8I?�xo�xu�.c�Yջ�U��.<���C��ݾ�2KB.���F�g"�R:"=lC��LF㜿�wϢ:�c���ޜ�6�\��Ho����=ML����t�uw�V�a0ϗ�~Y�<��J�,�r˜�\�z��Y��[��⣤V�w��:[c
��T� ʷ���{�ٿ�X$azW?��p�	�U" Ⱥ�#D�)�,#�ִA$�ƽ8��|m��F����f���W��4�-쳅��Sp��f���2}Y�r��L�|I���e��_	���y����g��
�$T�3s��G^_}>='��9��K�a3åM ��ՠHvH(U�X|�7���5�>���mfq���iuRM����+��*��c�[o˙��q#n���+����9\�!	|�h�է��v��J����,&|�/GA�Q4�O`�W�����]ʜ�Rw�Z9�lX�S6S�����/wg!�#X�����GG��@]����|=0%���^�`�u>�wA՝���u@����Z(�BM7��ͤ
x�f�k��6^��E�C`�|Ƹ �sf��u��$Rk|������YcpAO]FZ̫�.����[z��'�qa�&���)>�Oo��Ӣ&���袋ɩ�N��,&���d�@Z�����2������"S�'��k�&O=Ɔ��sϣ��p,d�a�D���jk��D"����f;A�k*�C��ts��v0���r��Oy��z\(]�r���6S���A6��1����ɔb�fMy�ܮT:�y�*{\/����>=W��
6w��aJ>�vP��*I_�)��oA
aèBL�I!��z�p����i
���e��䈋S��s߻�b� -���5�[+���ǻB���f&ME��gh\{�Y"�#� �6d��@K�jxv���4FF�GXc�1S�_�1P"� �� $�<9�P�����zs�'�X��Ǥ�xc��[��QKq�����Z��z`Ƽ�W+@3��wR?�^�t�"7��f��
	J��t��<L�/�'Fiw�l�r"H�|�.f��+��q���Xc��e�E����c��c�T�E�s�s��C8�9BzN�ڐ >�W�[2�&��/��鄩�.?���ҤI;z�g`�C���*�\V����mē��OH��X��b-hH��n`�:�o��H��aN^�=f&PeR޼�aQb2��b6�,��,G�FY�֗�8*�V�V�h����~�I{A�������ym�EB&d+K���4/ՠC��5>� HV���'���*��m��o�cӞ�| �B5�(���Yy��C��!е��%���1��"��G���Q���M��D��wR`J�°+��h��6]h�;p��XnU��1�'PGyR�<����
I!:1 d�
Uռ/��8d��L\|��Ȧe��^��&��_ڈbsh���f��,�^�i*��J���5�� `���g{�Lx�����Yvf?�{sOV|�%%jX�J���3���_c���}�ts)����1Q�c���Μ�&| y_��Ib�E&���I����=�����k���w�e�%0�Q���|Dp��q"�h*ОS������L_��폜����k���D%�#֙`�@NG��ƹ(�ɬ7��8�p��u!@f]�uL������:ݻ!^����0���A�x��gǝ�r��~2�\��?��`�TAgk�~��&�¹D�����e�2.����3��5��h1�rA�I�S�Y3aQ#�Yu|�M6�k��g0�%��f��1q�������:�v�x��m�v+�r�\�05��U�zJy'�t��F0��+7�l*�J-�	�H���t�e_4��+���^���c�r�9�k��:��UI�Ekbؓw�Y�T��<Gi?b�m�����MDΧ����X]$��׍�.8,�d�����L՞&m#���@c��q�� `�P���l��-�uc�x���E[�WOr`Zvh��bK0�|)gx
#Ӵh�{�ٞ�\3���c������!�I|>�G��TCs��I�s�%��J��^0iо���,�C�o�Ӓe�j {�����'��M��d���EK���hq-�|3M�b��T��(�_iA�	���[c�����?�����Ό4\&S�i�6�غ ��n��T:7��9M�N��%��s�/v�I�
���Kf� oԚ���*d�;�R��t:#�c{�R׿G�u��� ���`}�!�i*ovS�0��Y��y�<Q�J���Q����4���S����u�zE�k�:�B_��fa�O���La)>�&�e�`M�ZΧ��@#�������fN�>`� 0�U�yp+m���C�e�J���Gm쾒�vC����"pF�HAq�Z���zxP�;/e֍�ԑ�e��b����j>]�q��=0%�n��8����h�1� ڏX�Vh넝�B�E��U{�����J���H+�����j<x�`9U�y�35DP�Z�7�����˲Wo��0�&��(b�����{�u$we`�Q�Em���p�~�E4|A
E&��3���p�B&^�J:�o�+<�C4���i�����1%�V��<�'�����
���,<���L�X��FX��8��wfh����ɪ�(R�Sv�d�����Y�l�K�I.��3c}���3�����k�z��ѯw$�����cw�1�#A�(�#!�W4��%���ԟ�I�� ���o���DYL��}��3f ��i~֐�N�즣����6����f0�A�ʤ�9��әI��±�ޮ�N@��,�՘U���r�h�A��lJ�)���R��W�N�=� ��Om&����Jf�f�azW��T��?�ŵ?H�X�:�xÂ�V�8B�ܦv-d�~	T0C�'�ڒ�>�P z%U8q�l-Uq�/C�\p(u}+��L�� ���ؾ�\��	�i�r�� ��zU��=�!^�B�$�����[d��a�[�8P:�]`	�}�(�Ii�X��v�B�c�]@�vS �0iؖ��D��C_#�-zn%��*F�[��so��GF�<��F���3�����<�+��h!t�|�>jʆ���12�S���!+��Hq����<��*K��5f?�ޜWߴͦm�f��8��f稪U��U���Yl'�Nᗟ��� �������}3�a�U��C�;��8������@�-/Q��xQ:�B��&b_v� XL{��#�5Iۯ�U�I���:�L��$vP�MJ���n�RC��&���y?�
��<�v��.�B�<ZK
�O��:O�M�=b;ñ�V{��6&��Ӂ-��7��vU�()h{p)����y���W�|g,��ˑX3C�������%��lV�;\��{����a�[���Y�`�*������(�3fcI��j٢0����{tӏ�&���|nK�f��U(|��^��� ��qI��.�t'⌷.>���p�0��;����Oe%�RƢ�iJ=��m�c������<��ь�<�#���B�@��k���ۈŖX���s*�Z�J�1�l���Sg^p��Ƽ�Bï���ܓ��2�ⲗЀ�
d��* pVB��0C*�A�2�_I�7�7rx����R;�x"��'}K?iyKl�{�ۺ����@��$<`�]���
BG�Q�ԳE8��������z/�WW�@Ng��7��$�� ��  �H:��u��$�(	�#-���8��l�O�[�X:a�$냥7bdV�����]+�{����]��^���7�i��f��I�g`���a��~'���o�Pl�L<gW����`����R�D�4�|�	��	�lJ2�&���#o:�n����+�L.
��cRv� ��+���{�,5x��`M2�nXL=��N��G����L<�
"(y�W���)x
��5�����VW7E�n���D#�����iU�W�dk
E@<��eƝ�� �v�$�L�]Av�a�Aj�&f~��T�����XB�/�t]+��� 	��  �)��ª�wor�o>A��B����8�-�������z�f8���C�3�p�
��/����ڨ��x]ET'aW���	�Q>�������~���)�4PA���Q���EF���^��;;��N�h��,���xlu��wT�
V��q gށb䳐ie����P�v�M�;�-	��U��"r|]�k9fO4�N�A���ƃ0��5gܿ8�Y�so�>:�mmO�
!��V�}�1?�sk�y�T�6]���1z���_k�8�{�B�Z])�.(���D�,�̊P3[�,�s�9ےo�ꋖI�D�|Ԥy�����?r���)���b��r0��ħ��~X�K~�mgb$Y�ޞ��87��N��*����e�trl}v��yu�v۪e�mfv��m0Qf�n�
�pڢ^ ���Ѣr���2��(�C�<֡�.̝6�����y:|���C��;P<C��jݓ���E��W�ӄ���a4"�X��Qa��E�����l7�Y��K���݃���g��!m|�
�	�����,B_�t�/h�@�����SJ�������]U��dP��[��Z8;�F+A媼�+Z{�-X���X������I:5�쏞e�(��0��)��r�k��0[����;�d�E�D��طGW���D��L��Z�^���߹z���˒k]B���a~��sOP6e���K<�R�\S�ݧ�\W^�'�Z��0:�R��6�@G�J5�RLQ��I8�M5'�9�����m`�����&��qe���d6��wP1���	��\��]p�Wf؏�m��sJ����� 9,�+tz6U�����;:C_�_��EM�v[~j
��t��� %˙F^����g/�V�x��_���^�9X�M�#=`��E�,��YF]����Ό��'K[�;D�W�4!�ua�������d�O��t��I(�Lk�Q���=e�b(���%�K��pQ!������n"�r�?O�j�m�WT����(W���E^��h1�Z�u��7��׿�vMC'�������|�F�
JO !��7��$8s[�sI��QV��ȱ�Ȉ�3l� �K@<�bLxgGG(I���J?����_�mx4Ԙ����+a���#��*�9j9-�L��>���/	+���|�p��>Sja����
Z$��:i^�sc��3�>o0����J�\���P��|z;}��?��q�Ӂ�����e���84 &}�h\��i��p�����#��"����Q���Y1�wY�'ؚ�@�8��\5��?�h�!
u��"�v��~�s'��eh�4�G��$���2�s��]�^�m�����C�gk����h��N��0[�X�K��c��ڀ��M�(|VoA�;����J$w$ݓ��[{����Y�%u�V��Eƕ����(hhQ��Ʊ�0խo.��=@�����_r(;w��;��2�J'x�`ó���R��-ͦ`�Ǩ�)4j%5;X0�p
�K�y[Aj}��PY���3��(�C�[",O�����#&�A�������.��~p���rN��4�'W�c�*�����H��O ��<%DK�{���#ɅA��Y��Q����d&�����$�5���Ų�[,�	�Tz>@.���t�����W�;u��'m��o�ZDF[����z\�"�xOy�.J�m�,�����C�ZZ#�r��o;۞�����:����r�N!!�p�K�;7x�lw0���]����4��ϯ��{?�p��8tY�������?�� ����b0W|��P��8��M���Xۙ��S�x�I���Ú��C_���.���!Wڴ�8#C�s��4�~��-���-��Cw�v)��9D<�Є^A�U�'��'"��w)ԐJ�a��-�b��6�D��\���8{Aڀ>�O
RpNlþ����|˴�TA��|�57Y�*�
J�fyS��(6c�áSx������#�Y��֠J�h�&f,��ϋ��bR�}5J�n��M��;�����(h�� �E��Ƈ�7�ل=n�Q��!��k�R"t��s�l����Y٦�F�vu�6�Wx5�5"���E��S�7���s���pvm��T�2��� ���mt�B��Ps�Yi��f^����*��95d�����I�R���(%	�������
~u���']�tw2�$UQ%uy� =,�ج�B+�<�"]��uA݂-����A�c�y�G�~u
Z"�\-�y��ZW"1��'t��ކ6��O��k�����'��傖8�E#[����p9�A��|�����z&Nc�/rVk[��K͞Z�`�}�91�F���T�}��)Y��j�Ʊ�zU'�N���PQ,dX?�oF�0�T�5�R�`�Z�a����@�&��Ry����8���:��'O?�x\U�O��֯,[؈h�%��6�heU��f<��SЃ�#���ֹ������AY�a"�E�Z7o6"�ZV�^5k�d�^���5�*�)�]�/"T�h1���n�Hq ȐX�tר�/���_Ui�eq�$�����6���&�g�7A�6����#�!�%R�O���7�����^���Y���#�����0��-�1	� ?��_2zz�Z�����'&}�	���E2���G�����
�k��WqV��CC^��s��*�_��"ߔ�4�^J�v@�I��{	.���U*�* ��5�N�:}��
);�(/��xm3��cR�Ax�>�b�!�"�j�8����fi�|q>� �8B����ۼ�B
?���D���<�[�ԮNo���`������)ݗ�����"�fp�jk�,���ۨoYb|o�}Hh�dY�����,��L��C>g��bC5�}�,R�D�sFT;�P���&1��n�ۙ�9�Y�5�sj�!H]%��6�&'�;o��W�w����)Hr����帧#���-�|��.i�^����gډ����"���-��h�l=��eq�^��S���1�Y&t�WV��Q��C xj�ǎR1��:�;s'�����4�b���.֬pL��5�۷3�����6KR�?`v�(�7�GZ��η�Z���Ee�6;h�F�g�rڞ�c�w{S���PRv`���i,<��t�+{��������<�
&Vٚ����#dCw��'j��i���҅�%Q����t,ll������r:�b��ȬpA�k�3�2� 8���Q$@� z�xN��߰���T(pk�vah'�����h��4(���|�g8�Nd�ͻzN�ͷ�˷� ~�{}��&��m ގu��� ��%0>��;�>Z=*i��Y�̱m���m�8����#.���{vY�f`T�2�ԣ��*ɤء޼�j|�%u.�6���xAM�� ��p/oS�}8x�7���ە��]�΀bP�� z Ja_����K<��2��g�Gnn�:!qԃGo�d�/�Á/J�IvL����d�����_��u��=W8�������S�-���k�#���f����A�&g+WD�.��"�H$��\p�����h���{��4�\�S� �z���I`h�pCx��`�����N�+����2v��E8]�I�|X��3r�[]�|y�����^8t������H�K�?>���V~'{Eqi�֒�	��V��h������Ǣ�Oѓ��\�gQ�-����&��D$��J^yĸ\L�T�~�9{��	�;�&��^1w��,a���e�UV,ӡ��u'H_<�������p�L0H֏�d��t4�S���e���)���ҟaDH[S:��r�8�A і0ʦe�Z��}�ߍ�h�:1:��ϼ���O��� �?�&����Gf�&LP��PT��*CR��tP��Q[��	�am!����@i��m���	��7��{bG+u�ȝL&	�B8���S�zݮ9Q�9�˛�y�Ͷ�(�]�4Sꦼ�j�)9n���gI�=�U4_} �I�l�r$	��r^����֧(��a����}��-��{�[��*�_�=0Փ���a��#Ս�w���!�������F�0k�� 9~Сdc��0
u�z�!�<��d:��VD�͕��u^��b��p����TNY��F��b8��0)$c�.r�	_<{aL��:,B�E�+.!�A�ku`c�����>����)(̗(��ui�n��?h��VZ��C�22^k'ɼ����8G���j��B��ݷ��Z���g�%���hR?͉�",<����^;���9�n�"v�=`�؟�_��М7�Q�>%�@˪I���S&�5}��V���L��l��%2�zR>
#��]��4f4�[���M.8|�%Qa��X2q�K���zu,j����ȱ�[7sZ��3��Ǡ�ְ}i�k��,Ҟ0F$�|��C��&��|��}Bm`����	A��8�Áܴ�(�+	[�sz�u0sCQ�u0q{#���?����>N����\5�����G�ld�n�T���u�F'������hf�/OxL�S��S&)NZ%Gw�rs������~錄*�i�g�9����ف��)8E��a\�{�۶�� �`��A��ƙ\�j2��������7��t0�� ����~=7�0���Xۻ7�����������^�~D����h&`�'qY"�?�2MP�<A���h�r�?�4����M��E����X8W$�������~d���	�����b�kO�p~s���H��z4�wX&NlY�k�,*s��&��b�n�~�W��c���$���/��Y��j���*$Ԩ<���8�1���#V����Ã�Y��D�L��m�߈��;7(ū*��)����o?1"��j7۞�qO:�g�� D��b�D�ݝ����7� dC�����Я�����]�;y�J�g3�ql�o��"�d����B�C��o)����|+��ao4}��kn����ۤ�[��0]�4�bȁl���|a���6��,ļL5����D�_�B6��v�_G�[�wu�P+����Ɣ��l�dN�sP��U�o���A�#��x�b�[����-PX���_�J!��t�7���� ��O�H����Sa:��-�
|�,y����B/Y��+�����eP�2gH)�.fu7fS����]	��x�~&�
*P;�����_=5����E-j������#K��Z�l�d�p�'��@������m����=Z��Q~�S���NKOM���HvN�sܳ�6UV;~�G(�eK�I���u��J�����S=I�"�눹Ϻ�G����.z�'DiUFl�L��luv�6��Wpl���ip�nkE*Q/�=f;G����S�B5��Me�hOJ�uC�Z�� L�/�.��|����w�_> z͝\>7��c(�Į[눑=@�-�^C`�wGt�2�~�On�p �O���	�M?��a���QxL�G���36���3�9bSK�	_@�GXG1kF��4�:��σ�ѥ�o�;��( ��\��{�*��$S��ɨ�r�0 ���@'�=W9w��Z3����5�쎧��moo��B��y�uN��T����2�.(�ϞK�D��G�0K�ĚT�<����j	�o���oP5�bOS+#���L��1�
m�j�*��<q���b��|<7 ��B�C�b�vS.m�o��.��[�)h��B��D)��B��c�Ɣ�ݏT=����?:��Ve��"�H��C�7��H�[��yӡ� �e�l����z_sH:����:�]=�ot��EB�,�A��*1�55F�V�"NЪ�
�ܚ4��Ӓi����Wm&eڅ�2k�����+_`�գU7�լk�a����bn�/ �mh��1g�`\<���L����@Q�!��~�R{��_8m�?Iy��)wOu��*@Nՙ�VHL-�?�8�!>����κ3�+v�j�pj�+�F �8�\2A��W�QIE��t����x�� }��?0��+��/�*P�}��f��;�
�x9PBWic8�d�,c��sM8�Y���BCt��Z�lA�Kf��k2�[���3Ԡ�0�v~��kJ��p~u33�c�!�acߝ��	(�1ubm�J:%{a�0���F��Q�t�7d)���i��=�R���bf"���*�.�Xm��]k{�t�����'I���ݾ���ƅ���`M �;��ݻ����Y�~�T<���O�9x#�7�<
zR9�`�����㈙�M��ں&�M��6�)�������>��P8���1�>��K� J��T�я�R'� ���P!�؀[�e�ؾ�,0�i��L[_Ȏ�e%e����s�_-�S!���n/m���'OR*�ޛ��uI�CyY;�-��{|��1	�03f�z�V}�x+���9�ew3�jp0���n�o75:��Gp1/�7�
}?�d �⭟Ї�&>���+�d�O�Ha�tFĖ~$�t�v�F�2��G�5�g�Gz��w��+[J*�����ـiQ,�M7<�����=?-�D�۲�H��"t���0M�>N����(߽����TAEb�Ğ���Z�]�_b&����ݎ�`p!Ƌwr�K���{~�>"���w)7�p�������c���XC��S�C��}W��fCm`Sx� ��Na� ������RE֭&��uܪ��ΓQq�+t�j�C*��i�ht\<����i]�{ ��2�3�{����w_yQ����K�A���L=�V���>ѱ���Q�Ei5�og�����(=&�`�I�KG.,ו�Q��j��I��{t)�-YZ��s>)��b&���x�۲�p+�������h�F!��(��x��@v	�C��|Zx��5�my��~�	���"L_75m�l��u��p�)��fTx��@��p��0q�4��'����j	�?�"��I�O\rY�q	kj�u�C�m
h	k"�]/!ӐO*X�\EP�	�+����ϣXXc�B�,�C�.v-�4���y~�R��f���ăm�M4²]�3Q F��6$z��Ō�J��DT7~if����ѿhm��;f3����\����� �nʏ�uf�n�ʵr@�?��������4,7P��x�9��Wn��X�16�8�
�D��>&���a�9��H��N�\hS��f3�AQne���:}$"y�+>�Mӹz����d��G�,c*��e��!~�
a��H2��vo�J��y����	����.�`´o"0m�,�z����1��
^b�,��vH�H3����M(�ٞƸ|��U�z���w��`d{����(�K��/��:�`�C�H'A?1��i�"�w�`qX��7�4��t�#��M��{淥���$���g��*�@Q����M"oc��}6j<̨����P��D��?p�`ړN^-�7�<Sq��v�ZNn�9_/E]�n�����'�XQ�tJ�9�~K~jmS��t�ކr������4�����7�3��G
���t���UYߔ̐3�"�ؗ�z���ڪ�ˠ���)D��p5RT���?�	�Ź�6C�!ZX(�[���*FR~����7uc��k��HK�8�|/�B��S�huXi����}���<f&5-ښs���W5%~3d�Sr�Q�g2t0\ƙ����>H�\�^�g媍�7�â�_q�2�W���J=\��g��8gޞ�o� f�M��y���/� o��_ע��󯗆�����]�a��l+&]�� FU�Q�?�|��]��FP�A��5
�W]7�5nC!�6!�T�s�D4�t\ h��\�P�Ɩݑd���5 ��7:ā-ЌL&�fz�����2p�Y���9�54&���[ [���ѩ&~��'Խ�W&�B�Ui�M�Aπ�-+�>o34�jJN��<�A��S�n�^�X�`dv�{��A�B���~��vC�F���2��4S�}l]dtL"7�9m�0�� Sf��F	�<�w;�awԆ��ԋ�N	,	a 8�a}BoG�e_��k��G���:Y�lT�F7��'&V@���ᫎ�e)��Ċh~�>.����O)q7����V�4 .��������G+En�����Orr�y��I#g��G��� r���q�X�|�M�L�W�Z֏Ү�}a��֏�6QK����a_:hk��/��M7�=� �J�3p�[��C��3�S�҄EoѮ�Pކ������_��m\��G���U��J�3�I:	���b^�_�H�$�_Ԛ]pht3�������ؤ����y�������%�2�;����6p� Q����Vٻܢ�XJt�ͱ"XY�-k7MC��+�-�f���MI&���\�L8�Ln	���bk��E�UL����۝��H���4�I�;8���[x�15^���ZߵcqA3H�д|�C��6{Z\�&�Pww��i�D
��Ur��-̨g�V�8�[ݢ�Be��j�K�"JA�([X����X¦��a#�6%ǅ?��-��T)��0�Ԗ��Y�gs.���zZQ�Df�c�=��5`c�����ԁ�V��ym�K�����5��>����3��x�y��ZT��/lSV_}4�Q����{<؟�Iߎ:[�� 6�NI�f������������C���ʿ�d�z� RK3�]>���S�i��4��{�i�I�����t�6��r��i��� 9��\uhQ4D�{�u���:kf�R��q����[�˳<�[U�f��x����%�3��i��t�u(@t��,�;�}�G�e��)�moZCI�q�ݼ8f�;����|�3�8�Ё����8�%U� &��!�����,�	�,�K�)����,?�����*��VK]�i�o�.�o�i_L��O����qî}Y^�Ok)Io:��}8u�Z!���E�8��*��@�F�&/����8�� <��� y�b����ۧ�QL�\ u)�U�֟D#m߿J�����c�Ճ��n��� ��}��-[�9่avy�p	�1�
��L�֝ԝ�wj��
c�Vw�"�Q$\Cq a��� ����n��;��A����1�50m}ڪǔ����<v���;�޶�K] �X<�Y_e��`��'i�DS,�0�0���wSI[�p�g�	�ρd�j2������#ip��]����THЌ,�ͮF �L2�#�V�n�*ף��>��ܣ�����Dz��+n�
�A�����x��is�4�?3��,-�tßH����s��G�؏ �!���������"T��,E@���f�,�,$��
��lT~s���'����"1�р�X�l!x>2?�U;ϯ�� \��P��הq�*\��U+��[z���h�.�{�˾1Y�6@4�a-���%Bg�`	�L�%�|���
�dc	���o~�x��~9�9PZV��L�B�Q��-���=����.�b�" ����EB�~����%����=�%�&$�sW�q7�O{kdҌ/�F�?1V-{�P-�B�� 
6ٍ�N����0��.*U�X1Iy�oLj*�m\f��/���8W050!���y8"�")�����z�R8H��ѧ��U��K��"��ϕ��JC�Mp�9��U�iȪ�H�GȠo}�zs���%\�ld�.��4oyho;)Ѭ�:�ȉ�Gm���,x���%Z_$�=Um������;Hu�<���C��hc��7����]�����qn)�7�%��g<˸�[�G�mD�v0�X7�#3�ֺ��$vЈa��/}���r�<�	C�����Q� }A ���gt�xݨ'�!܍����X��K�Ӵ�3sN��L���.��R�#�0�
*�~��D*ۿ���kn (�%ȨO���r�����`I,��J�VV^�PRy(�㊃��[�4UN��.H����<J��}D<'���b¿,�3��V���k!�D�)��;�C���2�׭#�Q��W���2(�;�@'��[��WH�蚚H��;�ku���\]���'���1�)���������&\5!�u�H(�!�d �L �J� ���50������X�c�T�0P��;��:HZ��9$%��k��%
փl�h�C���XI+�_�&��I�� �=2�.�u9Z��?s�\��-1�I�6�K[��bDsx����[4�zM��[$�@�?i�R�g�	 A6��D, �P�N�ql�3��%��ꡓZ��!�y�
�$�;'�����&!)7���8��×:ﲈ��\Gf6�FL�z�et4�l��*��Qh���:�z�[;ڧ��=e�[�gH#`���ی�%�ay�tN%a����P��
��8b�[�IC�d��ci4I�kﳰ^tX�iF�IZ��oq��	qt�/a�@簬�ͣ��-4$@Fso0���HT��5x)iL�	�`�v�3I��E�c[�������W ���g�H7k}W�=�w@mp	�.J@^F�0�I@��V^αh\�/�F>[����ݨ?/�=�W<�p�1r<���{�}ǒC�eOzD}/�*Z�(S��q��q�r����