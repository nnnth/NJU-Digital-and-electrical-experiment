��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���:����~׳�jB%�h�cdBf�}�(���}��I�̜g���I]WUS���M�V���`��y�l���깋�m�� w��7�N��~[Kd�]�.:j�`H��j�|*$Hb�ZB�օ�
����[�U�ٺc�1��L�`a6}h>�`��ˣ�������=@��?�e��슺&+�6�z*��el�!��GF
#����#K�})a�Z�Ֆ.�2QG�-����h҆x�m�j?��yָ�6� �gJ�[B��;�E������mDz3(#�R�Ib�	6�7���޻��W�eHY��s+Q�y6��T�\�,�͉I3�����Ҍ���h��:���ִ�勞&�e5"��&��y��\/�^��lp���x��0�v����S��zW���	�).扽^I�r�<����a>. �����A�5*��)���-H��n���F���+P%�~X|�!x=�����>�;x����s�l��`�U�3&�@_�Y��ws��퉴��o���u�� #�W�mR�u?�iص[���p���$��G��O�\D�l.d��ﶬV���s�O�d��D7�|:��i3��H���`�\�K��{�D�� H NN�!^hk���-�0�����{��%^�[q}���G��	l�7���F,=�G=�\�D���ل2�����g6��Z�r�{�P���w$�v@(�m�5��NXƩ~��Κ��f��9��#7H��(
�	1�;��A2���f�M|q�B6�U�s)),� +/���p��x(1������#��F��]GX��+��}��H����c���g��biJ[�����0�sSGT�\��s�\��U%�q*�J?�qO[�á��Z�^"�A�O .�=�$
�������/�1�|��{g+����z��"N�>�EG���-�wD��^pU�Y��4�Cc+�-z2�n�=�5�_�����+0*S�E6�]�����Hz���{�P��a�����&��J������vѳdOm�a>$Nׯ�;>����a1����g���ѢD~����J��&�����6�3��諗��d�S2|�����&��4+�ǧ�d������ �f񲟇1&��o3dKK@U�&³��=KcG����|���@��UZ�æ�3Tu���Di�L�T�rӛ�l :/�
������2�	���Dfl6{��jwA���_��p]�2%��@g�	�ؑQ��)S}��0�נ@��2���,^�^�х�-��ţ.*l?���[�����_���/$��s�s�Ke(Ԑ�b�w��U7�zĭz�wB_��0!n��x��o�eC��*mBt��RL&,�E\���,u�V����Pn����w�$�-�~HPc�U鸦�e;�k�ߏ&�|���yKOi-���2{t,��'2���l�oWi��f\���+t��c�rf��+�m�;��b�u�(�ԩpl�Mk�����c	�%����#��`:di��E�K�Qr$�8��@yO�"9���/;��X@�"1xϥ���痸2�Di0�ؖ8�}s��y�K���Y*T�o�����(������6$K����&gU�o0�ݩSl������h��}v�!2���Z.���E(����J��AE#T�z��T�c`�Q�����)i�H����(�x�!��u����(o�7��L�2C�x��ϡ�,Jl��a�����w���4H�c��N�Bpg\�c��zrn�n@��Y�[�Ε����ҹ��]��%ۙK��¡�K$�G�Xd̂g �	*���fX�sH�è��Zf��e-Y����lH)��D�4sIFҔ�xL7܍��Ln���jx�d�1���ɱң1
�~�s	�����(�yݟ�h(<~V+�1ε�QD�2�$�<�Gܸ
t���y������͙���@#��*5P-HeFǦ"T��P�V���=gb��c*�!�υn�	1�Q(�z��qm3KR�!�K2ᔠ�������\�3\p�:�F~p��`[��Q��D�.D�I���b�zσ���e�Z��F��Vٱr����A�M��~���b��5s�	x2<;6v孡ˀ�w�����h�J���U��]�y����R�)�X/��l�H��b|P�*�L��D%O�hs���Xp�5ت|1�>s_$�d�[����`��������'X�݉[�Hf{�T'YEs|ܥ瀯��u��
��+�����C�Y�,��:���x�7�Iƅt��ʬ�/X�B��?��0-��Tj.�		��ksB�{�I��u	����(J7�bz���Zu��γ���W�"NE�L�����Q�e��%�Vh[�k���;In�|v���E�SL�����2/|L];`_1蹢�ZX��T��X ii�'^d1�2�[�9�2򩔈2$嬒;Ga��;��5�4+U�+�Tarr�ID�rZu�[�y�>� T�C�~��fjtV;<�Q��	M��a��O9\,���>5�����%>Ԑ�t�L�+^�o�^<��]�'��7�n��b�ꄋOrr^�H�Y��f�ة͜��ncӋX��n�e��l[�0�*�������!��/�*����W�TvC���Y����`	F���=p۝��8�sT���o��'��E�*��we�L�o*�CKKl�78�#�zp����<7�������7q�z�ޛ����w�	���ɑ�N,o�ù�6hT9vB{�):��>+�cO;�NfBT�2;�Ӌ�AbY5�(�:�O��J�P��FsƸ�`���2l�{w�!Yp_t��k�-ӂ]1�ɳ �ϺI,��[�dk+�R?8��Ɉ��d͂<zn��g��u��H��,w�b��e?(ox^���k��������}�H��D�(���$r˟K���F�*�������Rà�����4�T�N���@6��/3_�2�\��3@��
����yjz��INO��X Z�ů����a=��xu�=a��8�e�N)�p����DcR�Q�GU�&�/\�G�&_LY"�XJ���GQ%�Hp�8�,KD][���D����ͻS�lH�9
,��\A 1��<7O��޴i2c���hГ�ݴ�бҡ5�hӳ�����dՁ���p"��SKc�����d(���O�Ux���V��Gǟ�[ȗ�ݵ�:��[:N�#�X�܋щ�C�)���\tv��������̍Eu+�{��+k����83�-[i5F�n4|�,��J͘�vߠ,Y]�ƻ�R��W�������>���V�٣���� rY{�����������D5�F��c�˙|��'�S�����W�%⬆Ln���l]��w�p�p���A�+7r�r.�`LR�F{��~�	E��.�0N56wVf}��q"�"n'[+W��V�g���\/��n�F�P����|4��K��=!���� ����*��o�(}�9{Q(6�Eo������d�LS�P�o��xHG�A�cw�O�zt��"��Q>���l��m��˓��՚i ms?���W���d���y�/.�5_�(C��vh�X��g���*�$xA�7��fψ�s���$TU���+�X���ϓ���X�����h�cVZ�K.�w����8*ɱ�*���'x���mB?M8��9����n10���A���I�_ﶰQT����I~r'���@�=T:��&q�4)b���nLU�:�Q���%^@�m�{�7f[~����#鮷
'M'@�Q����/?[��+�,p����Y�")gg�.��ԯO���e����2ay��mp~p��>��u�X5����>���Ǥ�KK�b��:�`�d���>m�d���Bc���p"��M�Mm�=c��S��>2T�>��W'�f��L_Sd"ۓ�N��-��P�<��
qԶ���q�H"%��F��0n�w�6���{f4N6������~\'h	����wv�A��]���ܟ�7�/��lm����֒r�/�C���a��b,h�̌��4��h�?:�m�7i:��\�<�D�{p�]C���=�rN}�b��s,��t �cP��d�	Fd�9W��B <1���t��a�Nfg�����  z�����i����xD��7�k?ʶ�Xج��&Q��]��zSX*�
���M�Z�s^Q�\��2�6,a�4�v`���1�*G�B�~���:x +��z+����0)�I)v�Hڸ6��%������瘢٢����Bk�0<�JF�DDE��%�US��'N�kk'�.�ۢb�CM;vzkC}�S�m�e�z�Ү��&`�s%F3H'�$�yy��Cw�A���_����ϭ�)W�W�r���^��z�[?�u?��yi��j�+�B~��,C�v�n7�o�+&���3ל���r81���F0�+�L�崖��	�Ă�?��V��,�<����^�T�M���;��xQ�Q��O=����焉�3]�Efh˯�|/�CA�%)KC��a�5Vڞ�csX���eep�G��q��Z���L*��E4]�~A��>�bi��� ��	�x��;���Z�;{\@�TvNFTw�8v`�x��=�DbF�Q�p�p�!�Íι$E)L�T!��J8���4���Օ<��o�z�("/_sO��o����� EmZ��8�H7���E�iu�#%~.��|���Ȼ�~�<�/��s!��~7����5#�<Y4ԫ��FL���i����k��=��b�f�����o��i&el�PFpY~N�9,����@\*�%���8g7��@��F��3H��̠d�{�+��]s��:��3�+�2]�5-[��IL����D_#~�Y�w�E����S�[=L�I�.f;���0pb� ��9K#�3n�*6a=�x���U��x��&%oH�0���݅��4�(��B���F�ze�	}����4NR�Ν�[Kr~�b~l�Y6^�F0h]j�m	G����'�<�-�}���Љ��)����53�/c7�ӷC@.F\&�%D1	���.� J^=��@2JF�#CAɺ��x�jx}��A��w�[��C\�K��fy8<MR�@*�F ]n4G(52 ���C$�V�&x<=��Gb>C�3V�����2.L���f�<,�q���&\�a��8��#�~(T�!�>o6�Pr�;�J!�(;,��O��q0��㍁5\Gg鈖O�Kp�໯��X�^/-9}h���z��@�E��H��`u��w���*�Q�Rq�ԕY覊%R(U��7�2���/�o����|�z�����?�Ԩ�Y�5�V(C������q>���������ֳ�JJK���h������=oiҏX���G��/(�e��.��jL�U��;�����]k~�Å�?�J	7z�O|���4�Ffj	���M�k��0p��A�*��n�-���%	�gh���#&��g�O��U�2��Z&s�C���[{��0��Ƭ����ʨ�^����y0��^���V �R��[ \�����k�'��N��u��3~���B�m�%	�v��u`������U��O�g��|l�-���J���{�TX���U`/!������G�O���i�d`-�����7�P^{��T�7��zſ}��>���Q4�V ��C���c��;���S�'���3�Ǵ�|���H���_�����ę�s�@�NkX�2զ�>�/ߡ��{�Nr{�" A�#k�����QDŦM���ѧl#��c_�ʭ���rW��K!�Ͱ����k�(ZK��<ؽ@LM�PK�^�ې�;��TeO;���1'��~'�m�tʔ�V^珡>���8�~�⠙(��5r�_�%��b��ޖm��rD`�V]�� C��h?��l�1p��;xe8���HR��@�3�x�+�C�b�e��痮���my1n�SO:��(p�yD_�������k�S�2Oɺ���`�(�����'���%���~P�s�7ac�ݜ�Yi!k~�'��y��0���?۾7w��i�����;϶S�*iHIo#qr���}ʟA��ã\9�2�f�A��Ɋ&�u!$����N�fo?x$Xj�	nS�i�rr�B>�!u@��9[7%���j,/R8cV�5���!�O����1����
�R�sF#�/�����xQ6+���글W��A�q�.|�+呒z.�bq�����M��i�=9cע2�Z�W�_Vt��Ό��Tb���c*�N'W�	EF37�#�52oBog|/B��u��D������M��z�/�� �6�Td�����/�XW �"��"��;��̃�l\w�Īz����7:O���M�MF�]MF_�Q��1�)�
���*
���߻���v���i���_w齠Hۏ��Ir��������J9|x�6O�X��E�Ӹ��i��_mgC�T�D�l��d㏡���H��7�@�/Y�]�0~ŏ�
�|fN���-@�5���Ϊz5q,�/^'�o�AW϶�F����X�:�d>���<tBF�l�d�^ǩ�wvk=|��� ����(k2/�

������B�P��7�Z�V�{�.�i��%F��S�=I7+S�V�<8n�iV���~���|��kM�+���:n�G�{�m�{7��=<#0�G�,��y�A+#!,2�`=�k�R����4��Q.Ի��y�F�K����R65�?��_���~;��(��G_]�ˉ_��>�2N�����4�ϊ�<�M��[U�'�&պCV�!�i�-G(��_�m�4̥��#}�^/H��F�8PqU���  �U
�\�m�ê��~�r�n ܋6s-!�Cr���1ɧ;z/! [��=�2��Z�c�C���b��x@8��t_2/(���$��-�slŮVC,Ш��(�M)�Pt, �~�W�Nc|I�*����Jk����#L�ߛT��[�'3�L�j��2�2��������� �4����^�lMi�wX���Ԍ�byΖ�m�I�`�a��<M�`���"�`h������Kn˺{��x��Z���uc�{΅�.�+��w���m܅���R�u�,��v�����_E���>���#�z�ysr^<���&�E���� w�����0������~I3/��*��x#
��|ZL���#V}_���??�T�0,��Of��Pe��/�F�F\�^�8C&�=�Dsg��t�LT ��������Oie�^-���"����QK�O�w+ym`��zT7������]4��d'[�/�"�?O�k��D��i�Q�T��0���k�Lӟ	�ŋ�������/>�J;��r���a��\���6b�Դ]��u�;����{��D�aF���8锌�b��y=��ɕ%}e�)�+�rW+j8l�+���f	.�HM�B7P��cD�)X��p4��g��	`��!�d��:&��ᡳ��`� ||_a���v�!%t�;����Pp�,˲����q��'�-̒\Bq��3%sD �3Š!
�b���n��{�� *	�p:�Lrb[���!�M��t=u!*���zH�m|D\���U�>0�:~�&�#�C=�7�*=�-������`�<
O�%l	�@�J�yǹ&+�A��r����J�L�Pn�[�Y���*W���</�+��o5�9&;�0���
8A�ū���d�/�R�ڲ��ĵ�a�|2��z�p
��=`���1�4����s����59Lą?j�K��|�u�C����[H�yg���G�sBy*�Ml�W��$Ip,�#�ju4f??�`�>�(�Z���ԇ%F?_���7q>l@�)}�Z%�Z�B�Q�@2����k{��O�8uEc��<џG::w�6�
r�W ��ΕH���d�A����P@Ix�ZZ�+m6�<�B��G ������LbR�|��#n"y��w����I{���c��K�l�z,����O��d����5�@J�{퇭ᆕ���W���v7)a��:A�w>sJX*��؂@�����y�J#�h����]_�����(U��eV�?u���6��͔�s�e��[�U��5����F��������JW"�hS��H%�m�X�rN���Հ�P!ܿ���&���T��B��~~��O9���u�f���6�b���x�|�B�$Gb����;��_�u�4RG@	ˣ��=�!�	�-��z�l}���0�ٯ�+����(�]r'�<���Pޠ��WU���ʢ[ߘ�ИM<ml:�o��З?���U�p�u ]�XpD���F��`
�����P$"��t���Q��\OU���ӱ-$�;"3��|a�0f{�wL�B�<��W�y��\�jG��r�WD�J~�D)T&������k�ǰ���2_k�v+}�������"œ/#��!{RꕵW|r�x��t���sj��z��VП���w�}�J�*ܱ1��f�������[�DGka�?WKg�?bg�Yi@r>M�>.O�g"{��2: �2��?�o�� I�ޓ�	J~aR��C�9��(ʁ�п��+��Y �&�YpPÏr���Ԭը�銩YS�������k�*:��4}����=�K_���Ü}�����l�d�@/e�����RQ�?ʋ S��[e�l��c���&gn��V��n���~Jc�I�ž�&�B�iE��vV�rz���8R�Mf��敺s)���Q�����y����p�6j��$]��r���ܭ�,"���$�kʐ����m�:���QKΩ5FU[V�U���B�޺�N���?�����2j��cܶwq,��k��#�aײ�D�:�c�4�=5���#�;��&����;nՀ��ilI��E�Uq|ZT�@�l[��R�[-��bR��s��3��%���ᇊa��+�5^�t�i�%:��v�C��|���l�׉ԗ����������s�xb���x�;"���֝R�[.���=���в���	����#r1']��MJ1#�Ȱu�p�#�7�߂Y����<E�r�p&B0:%�.�[�]�!��	��Sm%�!sI��?E;�gʹ0��P��CPr���4���=����cQ0$Q����J��oL�:Z��&v�uSq�bH�x��h�6m m��qs/����� �p<[d�f��Y1Y&r��:8| ���)�r~Fƙ�/�%-��)��}9�d˝���ض:S���\>3_�L��,<�",`��^�r��oτ�Ӯ֋�Yh����p'8T+����=Ͱ%ގ�ɃW��N