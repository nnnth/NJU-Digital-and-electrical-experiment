��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t����}���e�%$�oA�jv>V�j�����MD�*ܧ)w�!������+И��`Sp�$��/�=_�pC��Ԕ���w�6��@;�2��#���t5�N�O]�?�� U���b��LǗ_��0l���,�<,�t��Tb!�#�f�F�������F��&lv��)����Wq�sȨ����.;<�c�K�	�Q3��e����nJB�a����n�PX0h���<GI�o�X���)�~�Ř�l ����������!tO'�B��]Tc�Y߯i��H�G��ie��*�.�
D���g����+N��i��L�-'�o( �/n�Qi�y
I�9@�jJW��=hߧ�nzg*.���5K7bݞ��-��/����u��:讍�d��cLyp�9����KE�ɔ����n �`��	���7��"�Ƚq�����=��5�-�VG9��9n���D�k*v�����z~+9��Q���̔'���vBi�>�ژ���WYS[�9��اS*ܟe���Z��6s��f�X����@�bJ��
�	�v�JYR9�N��쬕`��v���ʦ���v�7�x5!�:�������g~��d� �Z��q���	p�. 6�>i����?�ҁ�1�_��
��:���3�6>�!%'.�]�n�w5XPC�Mu/(2��o�5B9�������͈Ql~(E䕮�5�u��m��/��,@�w���o�-��n�ľYg2�z��%���6J��B����ɑ.K!�$\��6��c��N��K`[AH�i�7�6e�C�gP�m�^W5Ҽ��Ku]Ü��9�l�땞Ҡ���|�c��$T�Oq��3Ttb=D9q�"N�:�}9L�;'yuÍԳNu�qc���$.uS���9w� n�oԔ���\xk?U h#qQ��=�A$�F��s3]�(�n
 7;���Hǥ�nhM�^x$^+�]`�I��}ӈP� Z,�-�L[�E�YP �D̹�ʖ��J��풹t�yc�<��^*�.�A�H�[]U�A+*��u�V
Ɛ���ծ�^�u����X:��Uwo���Ig�`M鶭�!㒇�P���4Be�����cf���� ����STG��th�zY�&7��/�*����簣0ƶR��?����a:e#G���-��ܫ����A `H�E웺�舘�r�~:Q��}�wJc�9�(s���Yc7,>K��,��Adw�[E^�Z���4��'���2|�٧���<����OC�t�����>8�t�L�m9\8B�z�7�8#yP�>��o����K_������wH=`F�%�0̳\�Afd=n��j�g�h!q�}�Hq��J����s�
���8�5��l(5ʂ�ܓ���Щ`-&B����{嶆��u >���5^"��s^�|�i����'� Z݋�������=L<��b`�}����֫ �{R&|e�aٗ^�y��j��㜩�o�qY��9w�!�z��'9��6$/�FKL��ԖR'Z�R<g�5;�!��9Mh/�����. ��dZ�:��3ޫ z����s˕�����V���,��l�$j�&C�_��w�~�����"?�#�DCA�<��}�)���Pڔޅn!ֿ�Ev�B�1��`��+��6%�ƛRG�)��Bm������d��L;M&����X.9����tI\�|W=����iN�^<��{���o�s�gɧi�e/0���� �yȖ�<���0߬4�� BK~EGpt�.��3I#|�e�i�:�r��Ģ���!�*r I
˄��_��H�w	�6��a��X���Wq��q2*b��7�.��n#p�Y<j�ݐ1i0�M�U@=��o#��L��\�YXR����;�*~��V�(I���uY)1x�0�L�9P+�Y�ON�8��?�	�(�dKt��G��P�3��[rc�X�~*���݆��:��㄃�"Nw��u%�T�#�[��0%%�h��+؜,,��X�N�j	�6Do�{v��Jaɚ�}�)~�i��'}/J!|��[�4ރǑ&���kD����sop��Aޒ,���q��i�aഏK��_�q�e�6��1;�(;�8���xr���p�I�%��,���ev�ܙQ� B��U 9�B�Ý�P�`�w�=)#\��vB@��/n�#8(��i��a�s�~��
�q(��w/N(3��:�ܥ� ��QZ3��LamZ�t)ֽ��}8���p�R%��Ӌ˫�����	���^���"��E{�LP��HA��-���������EC�W۝.�Ar	,�+�Ge�I����c/)R���Uh�y��0a*d�X���?��L䒼u\л��6�V:��J w얭�{dd�Q��;��L�����cMg
-"_�"Ԏ~�����.g�i˯����ӧk9�ԭ�l�c����5T�{�8b�G�k�c�a���0�>�s�䆍��5N�rg��Ƃ�Sk 1k�����b�Q�{{֔g�Ґ�Ʒ15�d��D��]nJC��/g�5����U�rEYh���]�����%O_���	�#��*i�whQt��SF�,��������>ߦ���� �&�|aL�L�`Y��֞�J&��Mlޥ-���8�KZ��B���E�0|:�m|�u3���'Q5S���=YK���[���h�y;��߿���-3@�b/�-��zz�au�=Ұd2:����0S
�6)��rd�N�f��A�Cw�jC��n���l�������=�C'p�R>[TZ�I@Ƚ�U��Qj�	�k�-@�uPP���Z<����΢�\�'.�+%�]�*倁U99o�=r��<��;d��,W�@�~���="g/���t}n-/��}(5#��z��L�ƥcx%"��+���-����}���*�m�d���;�K��M/DN !
�����כ_ĈP�)Ϥ�tI��l��r2�T\���^�Fq�xk'�BYt�w�fa��	��F���6�	�]�/l��U�G<MuN� ¯�7��Wl���y�ta��{Z?i�(L���-Υ$cׯ �)�8l���o�0��^���&g��m^%���ep\&
sT2s��0!�wN+}g��{NK�|��I�f�r̢ Q�c�o�e�/�W/G�u<�zH}�1��&����O��Ih�=Ɵ$�ڼ�GT{A�O`��P8q0��$c�
��v�l�;3�7ר&g�qU��$�̡�)!��y�0xXYǒ�ER�ثD�gkf�J�"�(_�W\��a^��)��O�2�W	���7�I��'������	Y�Z�����0���b������"�Χ5�mӃ]B���3X���C���&�����;��	ӓ�)ed�森� Xz Ծ4d�cE�@:�7]t���m;�V}��^�Ҋ�9b�q}�8$��^�?��i~�\���|�z�w&�ٶՌ���jn��k�o�&D��a��$�0V�@��w3z��9)��>������kzw5
L*d���u�6-����szj�J����YI]���G2WP������8|}��X߱6�PpT����Q�6���jYp��.^捖v�U�h u}��P���@uk��@���6��>Y4!X:=0Y8@��Q�UX+�"܋UȊ�o���i�i�������65ǤG��"��Y�����l3S�t|*2�>�G���v�2��	�O��-������[hVݓ��\j!��y�)!?�6A�.���L�?s���,Uq�h{��Ec��������1P�n�n��d̏�ϡm�W-JS��Ny��,�*����J��U�z~�����-�b�&��� ���p6%X��}�P�4�Ɗ��<���������`�LP7��׊��V��5�p��P��l�3�����,��H��x��� 6r��L/}���t�E��/���S��9+x�QM�Vݗr����*Cm�s�����v�]mYO�lT!aE(O�BV���"���a�3�8�2��n.���A�@�A�ƕ�߇�F��*g�d��f��vXuf��-e9`ORO�V��VT7����f�`���hQ�2G�ܻ	��O�}��wJ�U�L4I>�ř5���2���	W���A�$�����(`�n��Ha�a�!�����̊�h�a��qBJWz�j`��и�j��&>۟���"��=5K�ג�
���]������nU��c�?_�f)H����Q��ƞ ˰XA?�0�N�\��@������G�5�%���ܺJ=��8X'�$Y��*9���v�A��X��<�g)=�3=k��q��[��4Ҟ�8��؎<+G����QQ�4���՝��7��G�qqrD�.�4��;��_4a�@������k9qi)d�PК"�o�x*�Q�;�3��؅�M�ȯB�ķL�cZ�/:�sKB'ȤH��+dE�����hg�p��򴳷2��/Q)��?�z!�`�F��{V��2�/
�c�,�b5�\�Зkȑ�����٪A�4����D�~�4d����a���q߄�F��K3��̪����v3z��v�u�|?��?}�%ʡ���g`@p�5���B����v ���j����-XAZ>> ��HFOP�]����FYKï	û��&~��y���
q�����+�Ѝ�¹���M(`� ��ݾs���(������t�6��A���{��"n&�Y���Yk�;&�f{q��j�r�4����/���d���Ҭ�kj�B2���m�cD���Ŕ�$u�	��M.�7��8���CB^���(B��@b�����4~{l��/*�������31��vE����c�WZ8��X��8'��F�}PC����&�g�0����TY�w��_n���bꘌ�+u�h����$l����F�)7ng�r"��N�yҕ�d���l҉s�$]L�I����p�g�Tn��o�ц��Qq�t������LW�
��(:�q��x������4�FHj8T��Zω�R�9�}�8�����e����[F�̅�n�I���E]cL�Y�l�LY���3% U)p�s��FWO��-X0Z�AoY�g�0�(��_�V�����ͩ�0����v�����ib�`��#����/CڑGX��b9lL`���M$X2��m��z��Y���{�P�
vt�^��R��y�!��H�^�8�Zh�}��Lo`w��Ji
H�8��a�X��H��u߾X�,G�ދ�����{e��¥����R�m��|�/��#�uΞb��� >9R�����o��Ж���G�rP�Hܤ~����&i$l�c����8{T�Ƃ!/��H;}�`�×N��d	�iq=��m.GNV����tv/וѴ�����Y����9�ڙ%\�I�i%X1��ⅶk�| .m�ʿ�Lp3W�Ҋjg��#��n�ǌ �;�������`V� �3�5eЛ�+��R��B^fv�GӌL��8���ƙ���m�W��챉�y���~Q{�f$�@"<�����njM잃n1'�x��-`�;i�
��Q�4���Kci���'8⼣��4(�
s74E]LPmW�x_d{<�*pQ,5z���c��\rk��~m��Y$}ɼ�Arn`�$r	M�� �L�=�ݵm$�#6o�ڭ$] }Ӆ �)Q�U'����u����l��m�aKPb��Cw1��	4f�۷���2;hX��7֪�Z��|���r���*��� ����Um6v3���V�dO��)�H�x1S�4���7�	�)/����7�x �J��"���ƘM@�N��]z7v�z �C��4���9�u9fk�r�W��-N����xg|�pV�BscVm	�n��vv�~���yl&0`��ԁ*�{��ps���-}P����	snq�U�]�{�uĖL�����Q�·�)l���e�� 	Ųb�gZ�F\U�-x�2d<eQ@��d �o��p�z
IC�z7�9,�Eda�	���p���=O�t��h�w}�.����l�3jW�1}�@V�������A.�h̎��&����
ހ~�q�'$��<H(�E)5"���ůX�!;>�j�aC[Zy���(��ܕ�3��T�Z�wĭ�9$��@g�X�[ �.�?�䝇�y�S�-�
�E����/�ԣW#Xr�*v��S�K�d09�k��DUç�<'3��ڔjh�6t�u ��Yn�ER����b�Ҏ7)�� �E�T�kS�w��we˔�ǿ��-�je�T�$�/�$���r�xn��1Ь�ҵfG[[b0��j ��jŷ!e��0@����.͔�EY��$)&�;B�|))� �6Q�4�4D}���Jύ&u4�(F�A���ڀ�:�X��)k�� /��߹P���x�m>�*t@�M�;�qV����)��D'X�������-��aӝdvV���Oʋ��(G�)�.�\|-A�"g]"�l�:<4�{�9����#^Gω��@���Y9�9=�z��o57k"ڕ�3J�Fi;'�_p+p���Hd�}�p�1��1��2�d�����R�N��}�c��anet�Jʒ~e�٘d"޳@w�:�N-ӓ�,H[ʄ��� j8l�3�A�7l/�KL�E��zmz�9DI��몐V{���PAF������%��+}������3;+uJ��d�e�N�gbK?�UWf�fW�H$v�1���My�F)��B˓>�����J�Dۭ��ahμ��<g�9�6E��U!jC̈́������:����#�,Q��:o�`���C���d�Ѡ&uw5�.T�B$�x���OU�[%�l<�SA�߀:�V���CD���ͷ�yЬϨ�G��Ӝc����YD��H��"[j� P茾�;�h)�7�
���xؙ��UzCA���l����fZaE
S��j�(�aB ��x#�iI�MB���SP#�9R��i �(Jk'�����T<+�ȉ�)7{0".s޹̓U_+��PX�7=k�x5���u��у�G1	���=�O=e:�	P���JEĬ����D��U5������8�e���Ϭ���N�|r�Ű�Ԁ(~�3�B���ȉ���;���r&݂0�j!��E��q��A\o%!P���%�I��;�R�[�9�V:<�
��Ш�4�'v+�o�����"E����6����Z ��?��O��6<A~�����J�/d��O���-�R������(�+�B?>azkȘ�xX$��DM+���Mls���MLO���}�����Q^4�3�Il]�?7\bK�ei�o��R���z�
NʔV ��N�A��J�������7�i��\��ޛ���!A ��U5�"-��Q���^!}��:L��A��������p�����J�|�t
�"p/��=���fܽ*���U����"��y�0��qi⓪a=}���[]u..���P ��9,@��sg�sF�� ��a5�c]Ϭ߹�_�Ykiyȍ%#�8+/�f~!�6ݻ�:*��������q'�G?
J�����F�OLc�n��./EUk<L4)��	�7C	 ����hcjA�ox��ڳē�o"q<ג��~,�ǃ#��Sc�΀E&�"gQ:��q�:7o�\GF�,RH��xh�\�]��^��,7>}��V�R�\"
$�O���N�į�Z
9aJ�\7��D~sS��� �%�a=�k�j��y?T&���$;�X��T��Ψ�����K�B��=O2J�/���������L��g��!^<Y.)�����Bޘ�,��وs�sI�)���Q���)g�jM���79��G8X�"5D�b�mο���`'��B��w�C���M%��9F�E"W��ˁ}یGIP��xm�ݔ/�%�C��.���'z1�����	�W���}�V��@@�s1z��t
0b��DSW��3��D֟5q���̺&bPE��� ��Ϋ55NEdQt
���]��0[�D��G��ga+и�%eu�%��8�������n��@����d:����"�fF���H=I�9>�������a3xl���r��ay[c[é�-�s���˩k0�z�F��߻f+�29WX�f�
������*"�$�+9v�ޱ}����V:pN�p�i��u��<ºE�Q<��5Zptxx���P'�<?�dt#��U8�@Z������)�.�f�i��f��z�E�q{�!�V-�x�ڵ��4��Vn�V���t�A�o��Ա�=������� Ŝ�3��Vl`�x�דF���jDz4{�����w�)ݙ8�ީj'��Q��C�q�>��*�И5�!���XN� �2�NfGAR�W��6JYw�@H<�f� �����1F�M���Va������2�Us�߀��*�����a��hw�ݤi}i�xOxrv�"|0*�
<�a���*]��_��9^ˊ��E�.Xe8OgLH�l��̋�B���"[��Z1=|����y�j 4JF}_�U$�w8 )��*�P[N�rN�
�N�����:U�tmA�R2���M*�2GP�,��ƈ��H�������'ܻYVN�+���ƟhJ�~4Q�.�V[B��jN��J��C�e��).ʐ����	3���dQ	��{P�q��zµ��ܓ�UT�����	�*��e+����(�����o�*���N��m�y�� �f�R��G�
������a���T��T)p*�I<Ƈ(�~J�W��Z��f�
@�tT��1�4n�g~��7��B��J3ǌG�$�l�*�A� F!g��o���KY��0�
%�G��g�E�QB�e4Z��X,d�Ku���ڠ�)����#�p�Bh�1p��� ]�	(rh�'��x���dg�h،g4kN҃ߚH��ld����K��BO�cDfu�W�/��URmv����
;�nJ�	�'�ӝ�%G��\��D	d+��k�m�"�
q�;9F�Z���!{�e �xӳ/RON�0��p�5�m�N���:X�tgW_J�6��B��U��Ҳ7|� 3C�����u���8���qs��F��`"]�4\������%{(�`.Ļ,��$7��MW�A7�,Wn7(��;0���������}�G�Rocr)&���dl+1~��Q9��V��J���vL��F��D��FQ���v����n:�+��8$����}2s��`�]dP q��%2���F�7j��T������p���s��M��S�դ��܊����?�K,���aO��`�Z&w�I��nv/�J]��8Ԋ�	��V�|��v)E����[��x���������b_��b&�i�^J��+ ԰=�d�n;H�݆=% �w�sJ��M t�A�+E�q�²�����kP��bx]�@#��o?�jKa���Wk|}kb(=2!h-�E2���a=�k�P�����@|�f2��w�����jnVu�rׯ�J=Hx��1��ڙK�z�R�R�غ_V{�^�F��3_�T�.�G���W,�Ԭ����ʻ��I�t:NV���N�_@� �gQ��w1x�]��	��S(F�vZz�HJ���g\�����h!^�SF��,��	F9��Ac�y0҆*	 ��W��^i!�qz�m�-"�c�$\;EY��#�m�(�|;���������1B�T��t��U3�k�i����ӢM�Z������S�tj�|��H1^J�h�a�3��i���kG�]�@���A�g�v�ʮ�S�[dT��c��6×f�x�	Ԫ�Y.`	x�f�(�Z"��`d��<lmb����
U�*
N�u=�.����.��;=a��k�ydpy#Ͷ�-�7��y¹`��5 �C�0o�g�GՓ���I�и���32{�3�������E?4,�/�%�m}�`�?C��F*�1�ۇ��TҸ/�rhC��7��R]C��y_\�[`- �4�h��RV�5�����P90�ݵ2�/c}a��>����?�T��YK����1�<q5H`��(��>fgV~66�합���X+SE�%|h����P4y~����X�L��q5�Dh�j�Xń�v�D�9J!�vr3��`�c2fk�~uvD�)��X�w�Ĉ܋�3�{q���A�%�H�kb���1�K��E�Qi�~^��C}��SZ:�L΋cԥ������`2��'uc%�w�OEx�*���#��9�^�O(����I�û
��v+�cu�D�΁�����RƜ���AHT�އ��{���J�X��i�������3�tقK�:�%i���8�a�x�g��C=[�"�"�B�i��ȗ��.<p5`}��ez{�������r���ՍN�����
N�Q>8@�s�ӯ�i�&�Ԧ��V����ʅX��l�~���:��`:�k�����Ѽg��e���Z���Ci��N.�$�낻}���ё���bճJ�c���dq.%�e2�ϣS���E�y������d�3�D��TG�� ŜQ8vȶ�a��@g��+�+\C�����1��8���*��ShbrZc\��gݗ�"s�#�Ǹ�bf�i����=9M�{�!=�;3\ZΓg2\�F(k��{Y�'�����;�<�Si�"@o�x�ONO�F�E�W��9��:�*�s6{��1�%��^.�HE���|ؚd�?���> #�۝�� �^A��1�P�{����%������Z	[��g��|9;�\����usܔI{�[ӌp#�RM||ɾf�5>�um&��x|d�q�|��ݟu�i�a>5����V�vQ<}wn+BV�����\,���Yy�^��ɽ��44Q��O�H�^N{Y�j�5C�&�^̥&�;!�w�����F��y�E"���G΢��w��V� 
�'e@!�Ĕj�o���%���oS�i9��[Gao�+��2,�I#��F�05�͉T������ê	(�w��pf�nxyf��dzZ�5�	y�rbt�a�4-�Ev�����퓦�s ���87���T��V����.��He=�'�Ţ��E8~�A:�r��A���H�5l�ƾ����m������J�pB$e��#q��vX�Vr磢�Am�<�=���B��Ӊ �h�P��C��=t���1=����J��[�!��R��
�(1���������؉�)1A�@��#���z�5�yM� ��q�A����U�g�+����S^aVR0������R�2;L���uW��cP֫b��k
(J���J����.� %*Ǯ��Yy|�̙��q���(��K���|���SUE��=3�o��eq��L��f&�D��$�?�@���B]�]�MT��"�%�o��c�#p�:3D;�`M��pn��mG�k�u��u�}M��נ4dQ4��'�=�g~�i�\�h��W�:K���M��"j$�6O�~�*��}/�0��((�fAw�䝣��쳽v�@甆 �{�m,C��D�`B���-��fߝ0���E����`��ӎ���䒼�S��}4�Uұ_���ml���̯=��N{TvCa��}`-،�V�B�I������F�����G����Xy�·d������M��m�����B[;�cI|�=����E�I|�o�C���;a���k����=o���WH�֝��>���X'^�M�4�B{��Ið
��`�~�!7�Q�s= ��7�5�#�b,n)����B&X�B����k��VTIv�f�y���ω� �������Sf���Ѧz�=�� �䓒	I���o�OS��2�
�` � ���Q�����\��eq����� �]�vV�w:F&=FƠ>�<T̳{l�'�H/@��,pǃ�`�q�@�p&�<$ӆ���Z�K5p6&�����r��~��g+��' ��dQ���"��ha=��>2�X��*����s�$��v2��Y����5U��a'�!a� ׁ�,78�D�	�J�{����§=M6���hu���hw���\��Ԗ��3�*n�&|��&�YI{1!�9����|�����p���b����s�cbJ
�-���8��!���~�P;�����W��(�٣��A�m��7/ۈ�6�q�;�+r���Q���h�7����S�\#9Ȭ��d���2x����nF_���U�0��j�+������H��p�F��(��cd��kDf��W�~��IU��Tf491�t��d֛N�$cg,J�.X��,�L/���P�:���ɖ^�/���z&�"���[\c������{!1�~�B�EJa�)ohg�ึҞ���+���)����Z�{���2�!�����ư3�C�q��#�Ӏ�pDd�O�|�� 4t�����}�np�t�)��Y*p��da}Q�S},ȗ��/�4x&s�ID=5~F�Ŕ���SER��Ӓ�����'�8ޤ��Fk:�`ȉ�ܲH.�G���4�)�ڊ�j�4��y�?JG3 V��^>��`����I�_��S�L��&&�YC�U�ߓ] �?G���4�����p���wӯxG#ɱ�CY����Y��9늸O{��,����֊�5�Ƒ�_�G�����6�e�c�h��A�S#���6
9�vM���I���W�	Vi��߄���������|M�	��W!�&(��`%����G�F��I�C���s��k�P��9���w�!{P��f�,s������J5yI���o�e���p��u�����p<�{�$�@8��-������EI�C�G��i�����G�ha� �1�-��� �UD���
@�Q�(;|�I���X^��*�c�3���5�V�VA3�qn�zۗ��o�>��o���Y�z TN���k\"4j�k�fW�L�V��{��RG=��ݱM�tXn� (v?�(�kk˼�UI+�n��u.û��amk�sK���3[��Ӌ>�d�<2JLͲ2����XȆ�O����Ǆ1(�v�}9.'���7�vC�C�-@d�t�m#����S��=F3q!��wc ��%�T�^���z-̶��ʒ�=p��闚ͪ=	V�U/��7+UҗH�Sr� ���G���i�t�����d!�#�Dz�D�%���IC����7c[�{������g����e`�>&S䤨@�9�g� �,i�ID��x0@��ߜW=�=3ne��1E�0y	���˚P�<�h䂁Qr�O
���=�F㮝	R��?i�qB�lY��v�	[��!3P!��^N=(��o9�Ml����J/Ώ������z��<B`Qgˇ����'���m"�c~?s�>GZ�v�D�9��|��u�@�;,��]#x� t7�����V3&j恃�Bۢ\�� ��5:wY�|��#B-ַ�h�Z� �WJ?��D�t�D%{<#rI�~���υԏ�d�=mT�ֳ���|[������}�����4S%�}�������+��,�as��;� ����U�R���?&pd��]@ApA�y'��[[������%��wC��W��p�/0��3f�i�S����X#u��)��u|m��9���PP������%7(��td���#3�P�Lu\T�>��HDet6��h���:�Ұ�q4~i'p9��X{��Ϩ֛ԱXa��0l��~��i�Gdt�xx^��q�M*nҡ����X���dӗ�R_�"�uF�G�)�� T@���=��eTJ-1�!_P�Z���1��Lf4e�f|k~quj��W�!Du-7:��4�O�x�`�fi���� X:��ms���|�<�)`�~�x��]޼^#��K}�Ζ�_��*&�֪8��d�Nm�x������"�gQ`*��S������~��1����4�pT]E��~�Q�ѧ�@��-�{1 ��*�/�����G�O-��	c��{��pk^\(_�^<T]d���Wo:?�z}��&秳uR#{���+�㊘fɲ369?�܃���D���UG6�\M��Csxl->�{9>���ܑ)�Da��R̷u�G��j@�1��p�Utk�E�3�H���16�*�/YCQ�n�Hw��"���!F��U�^��աg�J=M�{����]wz	F�R��vs�,-a�LM>MpY�C�MT���G7PP�l��&H�l]�[ǜ�"#F��i��[�v��C��1yS??e�|`V�Y�:�@��y��� {�!y�n�lv���Yx������?�ʓ �����2�h��S }�#�I�\�q���jf �]�r��|Z��Y(����e����J�P3�ሚ����o�%C��s�̧�.*U@�z7��o����z�Sz�A��
0�.պX� ı����)��{�e���	�g�@F�AF� �%<w��L�!�ec�<�b�:Ik���e?
� ��qى��tp�Y^�z^t���AǊ��Y���ZN��7V�>�<Rw�xE(�v�����s�w���
�ю�qT��HUQօ�����ϙ7?AW#6ĭ�_/Ro���PG���C(g�4ުV��e=�K��JN܍��>���n]��R���h��->\��D/*��O�U�V�l]�C+�q�^>�q��-���`��Zų�t��$���9�C�T2���ΩV��:���%Q��,9�V�O���R��k7'Yke<�=-ϣ��o��t�j��8|�0Í�"���u6�Z9�i�ǳ���y:������c2��,�68_w��@�d�����<�
4r�#3,�0+�R9W��9ޟ�)�B${L��!� ɥ���b&d�^��%P(�K�|�>�k�&`��B�pO����	~|	@H��?��%L�pj��[����z�Lɢ����J�R�}�0㗯���Ӽ���}pw�*��O��kl:�y�U�:j�&�v�߮���o�/��O�[#�Z��C!-#�%<Ѝզ�j�t*oTa ��*:I4��.U����"���c��MA�X�vٹ@���"]�(ZCL�[��;��8��I=��xfHmd��l�,A�T/Vr�˧��)A]y1��<1��Ѭ~�V��x	�B
�<�,��6�3�v5+�Ѐɛ�[�ː�u&�݆ԯ���7���Q��>��O���M7���~�������G�߇�E��qJ��O7Bdis�������|�	~��7�4�'j�|t>Ҧ��v���)%�����1z�U�փq�(�m�U��D�=O��C�����hu}*����9fC�h
^T��U{�j��`C�+�9���M��V9鹡br��=]�r>�&�=ag��uȏzn���"4Ч�N��7��ٖ�a7;��2c<�J�J��b�Ҥ{*{j6+X2�^e�4eK0s'�ִ�����U�D�/�m����6P��P��]���ϖG)�|��\�R�'��D0�<,t��?�5��_w	�԰�;`�M�cl�	]�b�ډ��.<�]l��᳔6����%���S��x �v2���z���msu�0o���4M��U5�;D+�J�Fk�D�h��u�����g����zS���$A���P��c������H�΁&�(�<�laÆZ��8h`�C���r��8*f:��!�Z���Q�|�8
��آV��sO8q+5���Ctz�+;w��ݒ�∊+z1T�ͪ5+���2�h{Tvr8ԳKz�s��X��P�ڡ'v��%��W�̈��e��k�?uQ��(i��\�8*Aly����:�zy�R۔JQ�����66P�F�4T�YB����X�kM��N��ˮ,O�]�{?���z���@S����6G:��IV�}���|�����j��=)��=0)#�_����ϕ�R�T-4��"Ӆ��c�$ݘ�A�z1�.'��$�fʱ���H c4z�"��~X+���;K���.�Lf����3Z��4͞���W�$τ2J�\�ʰs�S���G\�<�\�;X#�hi9g��O�q����/G~�V��	�74B�"�θ<]qj��51���Ch��7�./�Wvg�cȢ+F������L�+?{��I�;ցY�.&&��J[`�<��ܡ�%Y�#rf�-�Èe�ݦ���E�*�)F-�jڤSRQ�yH�k������^�tv��$�[�Ζ��Ҧ�mK�E�,��[iSg�6LD��P��o��)�?z�\�լ*N�0!x;��V���}���/�`�Q�fΔ�`�|��Y��*l����s_k��\VF����J�t��:&]x�Zk���ڲE��T
�懐���g�����P��] '>k�]�%#���y���IfNI�Wxk��Tȱ�q	ӯ��6�A9.�����kp�x�!��blŽ���_j�<��䎊J��Uu�g�K�b�� 7XZx+@�$�P֬�&me�=e�4���d�܆��db�X(2vn��,Q�馐�Z�˲���*�aOh��Į���Uvg�/Z%���䊓UO��5�~� W*ި����q
���,�&�۱}3(n�M�`��b��lM[-r�S��t�$�RV�q��6BZ	u�z��gH�a&��&"�@ץI�E ���o�+l��Mk��&F��1���J�9*���΀O��@e�H.�Ͳe(�*�
����ӧF��H2HѾ���nv�E����[�HP����/ >���xb�1U��ޏ�;�5Z����s�$��/�V ��XOr��B���S��`pC���3B!Q�j��V��	V�\B�4�H啵L��ۑO�.z:(�Z#e�=���CsdZ�q^tfԿܬ~�'`2��V*�RjX�`��w�
����=��E�r���� �z+�׺�a=y�^.�V�E:}��#�@W<��������������bWb�\�8*��K�'���7&I��o�#:kֱa6b	�/E���5��ܧ���8Ʋ��h����K �Ax"���ޣ�1y�1lWZ�}4�����0�ɩW���UP����E��ݝ��Ì�b Fix�����U`��#�������'��}mly *�1>&1O�8Cߤ������Oբ�ˌ�~̱I���+8�e�m�8�y�y�*�H�Xi��U\j3i%�p	G�+7!%��`[h��;��vo��&�x����V?��Y^N% *[!���!Tu!UV�g�$�MH�`�D6��p��>��$_�w�"��tў&/'�����=�긠S�b\��#k��k�!��@M���k�ѻ͝�����褻!�^�׉�A��w���w���B_y��鸆f_#��#�j��b����a-����;d51V<����>�*$�3@��p��|����>&9;���v�����q&LW����8dh����ʰ� 0���㴃����\�Co,Է����G��Q��d&"#Kq�I׵v����2�'�:��쨃����F�֫+i���X��\�l�CB-��ׂR�J�j��՜&��M`4BX����WCޟc�p�����+ޙx�0l~'��Ǿo0Zjxe@G����4����`&�I��5 z���Fdt���f
����|�oh�y�v\{Ĭ6�a�b�ܡ嫛()�ן=���P���.-�;t%��Ҷ��z�^c�Њ:���&�]�:@(0l���P�v��݀s��|��]Cf7��6Yv�1|������ �2O�[�YE�����*�P$}X��+p����C*K��R�C�Y)p��!�,��'��)�7O'� ���)E�n��Y5TL��(�6�#�,=�a�I�Gy�h� �A6��K�Y������V�!��_�M��.�u��n^!�m��t�S���Q�l�����I��("�R�� �p7@��["���%�x�%���~O�n9��[j��l?��j�c�aQ5�e���F3�'K�~ѕ�霘���U��iPZ!@����OۖP)5���P�M�c:(&`��RV��O�}l��i!���l�H��fΥ���LA�ߖ����f����W��W��'�t�|9�B�; <�{��:Fe��臊f���rGҁ
����[���y�ok��R�J��}��j+}�Z�[�Y�����hyе�a���A���5��be97b�8\�"��w2z=�~�S��Y�ǀ�u!+�O�]��{���O��߅s�ʝ���{�W��z�h�!���Bd��'��-я�O���5� �R���Q��MpV�܆���fu&.�坔h������n�7 U�����<��6m˦`�`R_lӻf>�U���>PkB$��]o=-�d/��$.�a����7��6��}�޾l*��*Mj�f�2��K�&8sb�� �ѕq���
&����̾�;å.��_+f&�@D�ՉF�AB@�!�AQA����X�F��p�}dL�%�K�~y]b%����3j1�^���	;
 :�P$�5)�'紎&�U�OF��h�����`��\�S�'��d���6{{&�����$��c�;ge6�BK��0�j�t�ȧ�}1J�aE}8�Ȳ���Sw�����v����8�� �!nC���ش~')��SYh�YC��W-����7��eAIIZ`!$�HI>և��a갨zji�qXu�q�ĝ��}`iZ>�u������U�}mȑ���?���C�&�L�6� kE9�˝�!�\�pt�k �9��F��
YP銼O�v)��ܥ�P��2��t<����Yo���C�m� �����zCb��X��M�o-wN��pK&Lc ����2f�u�t�W8�����/�0��
�H��JpjvIIa0(�W4*��Xv"�?�5?n�H:5f��7����A��[`c	�����2���o�4�X�ԥ[+\tr`���ʼ�00~��b��{s9,�PZ�~�2t��'�E�z�65	-�������"���|���5䌊d�֘������0��kFl+L��W�UB�c�'����	䍶�M���۠ז��G-���1!w���O���N��O�I���8�79�juGk���7-��`�l��X�f�4��,�57���xy�#~F��K���1��l�Q��a��c(lz�l
��q���^a� ��0 ��.2:�â�/U~ @�L�-�}(-� +TV���*t�`� �2���-�b��w!z��T��zQ�\5_U��L{ u��m���׻���ݾ:��m¸UD�R&�y�К�x����>�b"�0Hx�[�l�Υ^�����,AO ���@��K�Z�+��J�K��EQ��Q�]h}I!!^"��w�����Ԛ[?�yVK��sGQ,�O��J�Me�e��ҷRA�Q  p�4�:�xv:��lsHLsu����JA����U5���h���ؚ޷��ə�����:Qn4vȤ���`��滩�4�M��j62��e���ޥ�|U7#���2�3�c	�Oc"�ٴ��6۵u=pV^{��=��&(Y�HE1
�Y���fGW��ӵ�'Ԟ>,�aY �o+��4��E y�[?_�djJ��y�{W��#F���7C�ؐ��x�ӟ-!�=ԟ]�R����f*X���_�x����?��[�`�ui�%��������d���8��V�������!*�V��q0�$�U�dO��H��
}@ޥ�_�w/>l���̄A�o��3Kķ����c�t�x�}�?@J���I��0x��K1�l��i|Q�%ȍ��إ4�:�������9c(�P ��)2���̕�i�Y�z���[�^�ӂ�7�����{����\k)m&jN��^Xoڜ�G�jUjZ��rztwf-3�����~_��+dfѷ� �j��c�B�����-���B*�u�x
�}��m�0W۾|E�$#�+J�Cy�ьp���_��6*y���$��n��(�,i,w+Rq��fz�8��ɟ �y���Nu�}�#EJ��!�������U�=�/��X�~����	�-x5f}w�.,�U�{��!�����^w���3���(�B�~03;ك�[	&�s��y;��uaU�~+Ra'��f�_�9 �|��|&�v68Io,	��U�菌O6���xJ��]��˸�\]!���P�R�%g�#͌��͡l�Un$YTna���f�u�܈��f��)Q��.]8�=�{vp�!]U�GEJ��M
�S�c5'�����eL^U�:���%�)�z�c�P�N���~�'/�J������@;s��Tp��\���#���/�=��p�@�6!VD��J���u�/N&�����W.��������=b;g�zl��m�� �>p���3[�,�f�?�h[ߣ�##�x��h�B��@�9��3���:�7�>����T�{S�ۡ$�o������}����t�P铫�R��E��}��m�Y<8�m�8��;/� �6NjS��`�4�tE	mM�����o1��z��FxU��bz<4#�)�Q�~��X5��"������'��ɨ9��YS���2����`RFݰy*�R	��֥5��� Yq�l���&B$q�q���Hc��#�<0��q�p$d�T��� ����aKz������
U��ʽ�ֈFB��7����s�Ӭ�tx"}�k�f{s$Wg���� �t���Cqk��߼rv�������+S-� ������U�Hcթ���e�����a��9/�IAk_�I��sV ��y�9[f]l��	���,�6��n1~ȿ¿EF���#�M4dW��+�G�v݉8��F#�H�,��1Lp�!�*J�L�%���L���.��E�j�������4k|{�E��Ytmr�f§����4o����v����X= ����!��V�(�4m�x�������CШ�x�y���ځs)�d�������{p̮�t**߫$ʖ���G(�n<d1@tSl(�Uĩ}?�Jm�kWNn5�u�Q<�o�0d��Rۮ�V�l)��
]Y���R��:XnRB�*�I0��H�p�c?�wj��~v0�},�q�x�b�p�|���=����d�G�1T�x�P,���eՕ��$c��%�R��5ض7�j��v��oI~d�::<�`^��"������YnJs��;�*��Ho������lCDl�m��]i��� ���N�)�A-���=PD��z~*)N�� >+!(�l0}TwM ����N$�>��O[-�9�86�^��|z0�U(��(Z�&j2�f}}-di���!^���'�ƌ����"���eb�<�'�ʦcR�Ź��50��� =~�!5o�n�6���ۏAmʣ�Z��Z�R�s�݂L3p=�H�&,��+!��Qy�ڜ�M���2ҫC��ꤐ��������(Q�c��N�?c��wҝ��Sz�����'��P@u���/&���a��^��YE�_*k�A��/>��4��|����[h��#"�'�솜��Á�:�PnH֧������-K�K��X�fd;�����@���Ω�X��['�ߥ��?j�fӦ����
��8=u���--�]��~���gz�fO�1;���� ��3,D �.�`����\ap���C,��u�c$蹻W1�o���-#79�"�����_��'I�fR�)�ٲS=�x�z��bnS��>S�s4?��Y��"�fz���N��c�*_0{��D$�s��7��03�R�nQ��#�+���NZ����Adؒ��F����Qa���ע���3Ǆ��I�s�� �N��l��%�Y�&j�w����0j�.���?^�;&�,�IS���;J�Q�8���sӇ+&2j�����Q�|��S�����t�I���ԗ�ʑ�m��{]?)�R��0���	A�q�\�qEs4�i]��ja|kj�⿰b�K�m�(�u���y�0������x��7ms9����@rzF&��&�� H�&gF%W�Dd��+?%Q��W��D�E5��!}F�Q�Nc!V[�����w�'�YA����b<0����6���	Mb�^�U�}����wyA�.T����q�t�BA;b���A����H��E��/��N��MI���wX�;���Oȳ{�h�S��̉@X}�Z@k?C�J�A���\#p����Љ�eۿ�o��������*IS�%	@�\3�p���$i�ދ�BZ�]���pZ
�1z����u������%����R�+|��u��n=H�q�Bm�E���ިm��"�M��k��v��ɭ��I��	�ݛ�e��`Z���=d�H�_=�[r9�? �܌)u97J��j��A�ݠ"3���ia@9qW܀6�PW����56:Qpi�L��7���w[B�H%z�'T�[ N�؁�q��8���O'\k���s6�`��GH��