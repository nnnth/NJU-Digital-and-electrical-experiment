��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�����U�|4�}��3w���n��B�2�Y��Bر�An;|ܿM�MT�[�=��Kv^��L�`.���kS� z@����$7�.�'@y�>Cf�(t�-�<��l���|�A�!0K�_���{���%B�`�%�a4�>U��7:�ģ�-�y�zռ6��*��ܻع�QY����
~�/�����@QQ��هH=O��˷N��?�[@DtN�����s�Z��S�v���E�&�ai�{���6H�u^ҕ�p<gx�\Xv��ʁГ��걬�� �k
����: oiě��8��9���3��h����o"����Em��7]?���Τ,���\V�}w*���+�%T�¿exa�ӛ~NG���5z�3RN�'���(�RƑ�Z$t��f��=G ���gkӔN#��M�	©R٢0сT�-X�u1rZ�EF��VpW� ����S�i�QS���&Y/��
m�s�1�E�x~�c����t�=�\�		)R�vf���dV@�Ӓv"��!�*�Jӱ�Ԗ.yuܘ&#1����.���u�oj޴�綣!�0C���&�C/���~jTHN��� 3������jO�K�:%-T�$�Ո����i�Tg����!�DPX����;�.�RC �3�����c%�U�u���F�_����O{���c���~�W~䗳����"���0�`�������u���z0Y9+���bl�bӎ���}�<ބr�v��2�c�+�mJK{���i�X��~_�!du����M�Lf�۔	\��k���qA�����/�3`,��l���+��~"H>^H�	/�����I������CI�7I@����7�NI-��k�~�X?�R�VX��/8q� �|���7Ok�ݢhgL{��,r�s`��"��S���.�w:h�����?�@�P7�2�Z��q}����wS�G�g�2Z�t�=%!s5��o���]�;�"/W�1(Ӱu�n�(�����W��NO�Tym�@�Ǌ>}~�nu��x$a7#�')��Ԛ&Hf�.���"�=�Q��n[%�$��C�ȝ����q�TU�*�	��*�N�6�6�i;�cO�
V鮒�`�I��	ćj6e����YX(a� ����4�WϤu�ڦ��ƥ!�. ΰ�m���r:;�ٮ�3dh��X�h�/f��z��7%����&���L�i�7Qt�p7���i�`������9�5�/��md/�B�Y���s(П�R���s�b��b�Um6��B�'� [^���b��&�����^QF�I�G�ߡ^,�LI�7Ch�n��>&E��g��\لCtQ p��x���K����,;�${�*���BxFt^]7�@t&��a5��)��^�#�?;� �]0}��p%���D�u|����\n���ͤ�F���]��H���9s+;�>�z�]��, OXB�6�C$X���sP�v$@�c,jg���Sc��R�ޛU#�--���:W؎�?w.�)'��"��M�"'��=�r�5���[k#fW�	�}X�u,��^ɫv���],��U
��}��M�/�)�#N�4&�9�TpK:3��f��� 	�Nh$<�щ���KT�C�U�V�$�>����	D��N��[����c$����kz��]X����	�z�|�/yUDf�,�h&O��ݑ�!oH�"�py�S�Sp)��i�N��"=IGa��l��x������|azO�,]�yc=�]���{;Lzm��^nK�Јh^-]L��Nۧ?7	�|�F��ԥ"�E���y�k�5���G��.�a��;��-�}�������p�a����H��zS�aL��	�o��o^)4��Sl�������M�X��v=�kq���0E�Duw�ʺ9B�����G�>k�O�����;?�א�y2�:����D���$:`�πK�}ަ�=7>J�H�����Y��ގ���s��X��U����`�@�H��x��qV�@eՖ:	�	3k�p{��D��4�����K�F�.���7�U�#���5{�Ҿ<_z.�|�nz-�j��Ϯ[Д�c�~����G�wݤ�&�o�C�}����70c	�S_:A���X^*�",������m-Y�f�M-�$�'�T���.8NK�ݲ>'�t�K��:;�x�F1w���Z��à���~^�K��r��C�ô�q|Fhə-�5-#�������Y�Yk�;
4�>��2�wU���Y}��T��ĺR��&Z��jt�o$��T�ť�?��_��zL����k�}���~~��O���$��୨��SV-�S�e=謾����|������g;�4z._�$���j�@���	9Х[�e�\�2�HC�K����,�P���z��*{���+;{Z�Qכ��D�H(�1VS0����?�n�3W�'��iO}���� [����as��Xq�DS7�L�r�)�-d_v%���	�ܲR��eDh�W �޴Fr����[DD�$0A���.�O�ѓ��ѱ�j��#��B�v?��^:[p�dq�X��۠F��T��i�>�)��J�PZ���{�d����F�!�p�R�[�Ҹ���(9]3oح���(�+	6_�P����Iu\]��MI����FJ![�c�tw�ʣ����hm�$�2����@�T וq�K�K]�O����9$Y��i��H�0:��V���XW��F�TXkb�}���x�v��NB�Y'�~�N��$�����]�}��KJ6�̴�ˢΑq}�1�������'z�ON�-���rP�#��|S�7AymfЅ���X���̿�?��DK�X+35|��.��T*6�Z�G��5�*�����lF�Xj;v�� *�GWg�tY�:@�k@��.J�#�����W2�����/������g#(A�^��V�ل�c�㮤��<cċY1�W�M����7�3�E��a�˚2�l6�M�˺�1=�R��a��� L�;)��t�E��,M�����/
,[�����S��S�-��p�h�m�]n[ ���0(����2:�nH4#�S����>�okt����R��Y\�d^��xҶq�`<��e֡.���@����nD�����<'��Q���K	�m��q<Jt�?p��ܳ���0v�F�׍���WA����&wM���i�@`��_U���&�],,V=��0OB���E���O���q�B �a7W�0��+R�ji9۳]{�-�#]����
f]>�J]\�/t���r?n���-����\3���ځ�d��kž5���tVD�m��Hŗ&�T��w�`WYS&�k���%"c�0��	�'R7޾@N��{���bj����i�Zc�E^��W�FZ�L/��&}hP���7�'0�M?�ls��]5?��������\v�,�I�T�,-v@�|��F�H�Q�b9�	ǁ�U���	1�G(_�5�Cb��c�Z�o��W���	��e��i ���,d�9�}@�����]�B
� M�X��G!�n͡ꃣ��6� m��EWΊ5j2w�O���m��U��	�#@�����AdU:��w�+@�cN܅݉Gb*d7������տN�W�L4y�k����[(g�WA8T���7_��u��;�Ⱦ�9���R�Y]�AR���l�r�����ƋDHQV�$+�= ��F-zO��6nh�G��`so`���~�Րhv?�	
d� �r�LD�w�p�%�3�����8a���W%�JW�n�#��Q��$k��13Q�x۩tȨ�+-�����,�0�J�p3�aOO�����j��y��E�3� ���j��{ݗ�_G�5Ri���&�;������w�sҐ��	��{J�>�U(�����u	��ݭ�im�%�d=+�>'���h��w b��q��肒9���Z�nc��?�du.P�HQ�F..n��DP�K���� q�Y���0�{������m}ݶ������������UC�a.U��m{�B)oM䌘����J�� <��"H��to��7>I�:y�\�����,��;�X�X��$'�h �����!�<!d
�?a���ҧ��ۇm7�'8�A�u�k5������C��;Zm��$����>�r8Q���4c��D�q�6̄"�WF�"��	FZwV�����ĝ���dU��<�������UR�KJ��o��l�B�4� �R͔#r4�ƴlځ�����a�wEԟ�7ӳ��>L۪�-ca�|��hW-��~&ޛ�>��E-�S.�#�O��?6�FQ�n�4O�%z�^��C?��!���l��y��J��ʺS��v鸖x'�{��f�^�t��_��5�������Y8�7�-)��l��1��s�8і��U�k|
�X�g�6A��b�3\P���\����/'�KmK�Jb��i�z㆏���3��)%mf����r`o2^�=Jmpwn:�0�W�����w���}�O,F!
;A�8��J���0\�M�������?�?�W0C�$��>j^��q�)4�������&f��f���O����ѵ�	[�N�y�����S��<���q
a���2�'] o̮�7����^��;Kᨌ��!��L����^#�r���{�u�ī�[ɲ	����a�WB���56M=�m�O�B��4z���2~j&,�Q�+����"<�L������.��8�"��5�ׂtD]q�[�aQ���eD*��z�^��;"���>�t�-��%��u��̳��U#�n�a����*���k�=�Q�ޚ��N�b�?�AXN�Z-~��t��$�B���+������4eJ�S+0�����b#����'8��^���A�7A��>S�UC�� б
K	��f����sCr�2��Ηu�Q�8�ڪ�b��PG���\�q_����(uYK�FH��)"�g\�
=��u��-��Y�\�<��%�|���dѱ���l���� qoZW�-9��ڵx�[	�>��t�d����M��T�ԤrA��t\����׎�BŁ���G���#�{l�}2:�7�<�v�@���s��M�\7F��C��OA��j�qHW��ۊ�Sx�R�V��e_ћu�����v��
�ԉn� $IP�bBȃ��bB��A���6�4�]�s=�l�p��X����h:ɝ�cE&�T���d��o�	��F~�,T��d�|�C��-�� XT�T	#��� FP㎕M�Ԧ6Y�mIr3����w{��'��1,����&�����M�ﱥ�앺i�ny5�{M�w���|V#	[UJ,�yA�*�I��fK�h�3�=k��K�k�����Wp�<��C*H�"
Y���ĄTecVg{VBj�Ǥ��>����`>ҷ��d���"SƔEy�o5Ȭ�<��?�WH7��x�z�FFB�l�t��\^YI������L�Ll)�������[:�$c�v���D���{�0?7���-S��^�/��ڡ�\�=dJa<~ݞ��.�X��mx�f+޶����͏�n��.��-i��N1���ai�m�`b>��6W	���]K�����}֘m���wb,b��o�+�(T�e�y���������־uɸrk��i?�u����q-�:j��� �1)�3��(���oX�F��y��aoG�'oD X�`A���Bs��:+#t:ao�]�	��߉ꖸ�x�V*���C�\8e�_�� Dp���-�F�Z-`f�A6�U�^S�͇�JyC�G&
�x"z��+Ļdٕ�
�v�(�*��-�@ۣl���3w#���%�t���w��������d;ٌ-6�(`G����t-�C����6��hj������h��RH�{�:G�aj\e+��#�8���޶�M�����s:�8�b!�����-�V(n�b�C�nTُ�Q�6_4ށ��:���=~��r5 ��+����0L�Dɸ��OA� �Q��m�B�(��}j�A[nX:K�vg{7�N�)9��\�N�xR�p o�J��X?a�-�j
ZyW��b�ЅQ�ôrW��G�'L�X�-%.���4r��\�*T?ox���eg7�]/��L�Sޫ������!'&�DA����<�]E0Rd)���aj3:`���.*���u`���j�^GQ/��M0f��_��#mW;?����8�JKS���И���5y�H�ŕ���":��җ��%��ag
:(��=����y4���2M<��qp*��!���'��AƋP<�~��X�e-�T���]K�v��25�{;���m�ש�ﳮ��SX���@k6��
��������#�#Ű� I���4ؘ<��F��Bb�2��4��t�n�v@{"�)�t7N�?@����)�[������?g&�(Eb�lh�ı4n�M����as�F�4Ǌ�S�F`jX��OWy�$�n��L\��r���A��}��#7T����n�}�o`��s݅9ڧE���F�B�6�+҇��i�cz�U��w>S8�U"qj�z��3�Cv����1$Ȓ&z�=V������O*���/�5}֔7���\ 
kjuGZ1�,E�6�+�%+�.��I�jv����*.�U���1 /�+n��n��-���	��G�0&<Xd>^l.�t���O�GW��1��AZ
����[���R�Cw-j�����G�WԼU���Oz��q��!�<����Zd���( �M��
���t�Y_�t�2�Yk��jrEb+a�K���g����cK�(NP�؍)g�v�{Ej)�;?�Mí�߆�&H��bu �WE1K� �_�s"NW�SRu�w���4�+�B�$^��"�AE��b�ݖ7�W��\��´�c���,��X��*}n�7d�a��@&fy��n�K��@`�e���\�n�a�S��;���41[!����@��ϲ�ɫA�@U<P�D����qY��ّ�~�%:#R�a��MWZA=a{HA�R�NY�+P�f�?�V�o)$?̑��|��Z���M��
E��rh�t�eq��	���9�+c1��c�����c�8B	�W]V;0#�ڇ�nl�U8Ep��.!C��}��BL�N��@-��nC���{������*AX��+���9J<�$����t�(���&�&�}��`d�e�@�|�9#���\m�.e��gk�=�p�&���w7��)���ۼ��R7�%J<�.קq���������"��r�ª�WlPj@S��g�E���Ѹ�����=�bM�s�R#�\�Z'�����d�:|���/pm�B��ڣ<��Ru�t��j�@ՒŨ>K�+ ��Oj{�ߖ�`5� ������A��F>tv9���ǠQ|� Y��y:��!�O�ݏ�J�]�d)�÷�3)�w����!�lH�����[�t>�f#;�ّ=$wN����#��Ms/�f��kv��e����m�
� #�O�:0m%~X�f�j��S���$�\Xgq�N����tK$Y�l�@v�mw���/Z�ѶP���߃���-Q�H:����A!��H`�����ed���(ʗ=��MqT�͍�ێP# ��68��29`��xїf�_�o��j �X��w�gٻ'�'���'6���,��KZe�'	�����tS6�y��]�ə�>�Z��9��W�A���l�d��v��;��q|@�s��\Ó��S�)4��e�<Z���:� _�����к�c&3�n�zS�L:�A@�ރ�=�i��I?���@wM�칾;�"�D+{ ;"ړ@A��3��ۀ5�N.#H�>s�Ob�-ިk�YZ�GƛM�tyHn�W�Uʋt�Ų�ɫa�nH7m�v�����x��y(�ky7@D[��w2�;Jž��5�pZ �FC�b�=�VA9D�)܁m� ����+3�
nl!�S1v����A@&^m##;_�HM%��h)H���f��7�B�0��-2��L��<�l�̘���vpT���6[
.f�A��#u�>R�i͡���x�Pb���#�^�&I���ty0�ć�s�=ط)}`.����^���
������u��%�q��oRs�d�A�g��۩ɑ�n�jѯ�Ǒ�"G*��Hpp��?�"X)�$�� %�^]ʩ��I�T��«�;��-l� ���C��5:L�b0�e��;�R���Q� ��:���(&g���ӯ�_�59ɐ`������W��W���FJO���Q��ysJD�Z48 �b�$�����L�V׊jnߨ��b|��{�ྷ1�����]���v�C�"�/8
�r��Y���]\��@N8A|;�!l2�8�&8}>t���#��/�L�Ah2��=����j��ݸ'��>�q�:q��Y��(�<����6�[�OY�/�St���5 ���%�����!%�59�Q�F�1yK�"��$����}!z��aO�!���[rV�[Y����b�Vv�unMŤ9V	���{{�����U�5�V�X�,�_�9��N���猵�O|:_��8
ǅ��L��ٿ�
�&�]!Wc4�O��:x��촾d��ZhyPֵ�n ���7o��~QMǉ6��������W�vǠD�^�&m2�{0h���B���#!�#�l�5؊і����V�֤����*�X���G���|���\~ܲ�����5��&�K[��]6�3���Y�}-����mD� ����ܙ[���*8S�QG�f7ީamʬ���z�A���,d�a�#��/�<������Y�Q��^�y5�$á���p�Ų��у��$1����J>F���qk."�L� ����'{o�b[�+�E�l����	ܯO-U�?_�����g��"
6Xj����adN�
e8Iѵ�0��!����f���� T��S0�9_����:���A9��]���+�+�;,�H���k�?|#�_�Blo����I
wŹ���1f�ʜ�ݿ,G��e�H�ޔ�a*�۬�����$>@S�o�i�� C#�|P@c����%�jt~��=��|��o�荲�%'`��ӿ��Vq#�|���赇jB�,tq*Kfk�ԝ�.?ѳ��DX��󰨼a�&ءǇB��*��p����q$W6��e~�q��K>ԍՒ~�w4ƆmIz��@t�خ�k���=5��=V�
>�����/+�ވ�g0�U��v��$bB���Ǖ��r.Bҏ6橿��TA�{<�� ��7ItR]���ʨN7w��Z�a����_ �'J�y�u�EVt[�����tP�ף�p�x�bfe��F(��L]d���5-��R�e�yL��Y��nV����ʏ�όB�����=���{\�=%*��=~�>���NN`�]}xr�G�����7mg�'Ha��uީ�RV�E��@�F]�����]���Fv��k4��15��W�A�Y��XTy�����S�6N�]�e�_h�ɑ�ǀ�	!�0��+�{bkɴ�A����ք�u�{U��;��s�f����p�v8�>�v�m������Tc��{[Ҙ���F,A��F�?$]�H�4+ΧF�M�u�Rvz]Ph��y����Y�]�@�<G��Ê����qQ��}�sg�0G��eD�`#;[���O�������`����Ѫ��t�꽃a�gu;ۅ�d
t�t7�q�I���h�=M�FE�8?���c��$_����u��!�`�<�����׊�_¸2�ԧC��L���P���L���4�&!��A�4��O���R�gBe�ݫ�ASj���`�o��;��9���mBR;��0�� ĂoA���M3��u|���f��UQ�`������Y�ܟ��4�T/�������+Ծ�y�fm��~�6x�]��(+�	#U�Ny$\�G�H�S�$ƳdK����E�6tX"���_�4��#�e��fJ?����2�tz��ɣ2+$���9�6��<Ξ\fªi������{�Rᗱ������q�'4�j��e�xbq�P��' P<XЁH�����*,�Y��o�J�PrM~���3�8��xx���~�a>n�BP (��CQ��~5�Jj�1�⏖�"��KM�ԑ~��*�٠�O�g��c��@.D��D�;:M��9�c�#ĒX�8�`�ǰS�j���w���r���ZjZ�׈�PFP?�O���9d�7L}��ʍ��]+~z=Gem�.��]�8ge�T%�ƕ^�%عw{V�2�oЋ��~`��)F~�شQ�a
"�Y'o��]"�%C���Qc��
��{�K�� ů��^.GQ�- ȸ�����Y��׬[��|Ŗ焄�m^�&�JN����
�(�&�u_�	��I[ƁMD�S[���ǇP)��i�����w9$�)S(B��^����a&n8e�
w����Z+"U�&��{e�g�mwz�Q��dԚ"��ÂcI�RNo��T�LrXʞ�G����G��%�h�Y6=���g�9.�OP�7 �䎘ox��l��X�&i�O���'E_�_�������ꋗ]_{:�Y�s��<ޔR9���;?:olz3���Rm7jq\\����_���r^��D\�z���	����|.	<ċQ4� ��6��ɀ#F��ش6��<B`\r�M�Su5�$KD�&ɻ�W@�e�yIp�%؏<Kb2�(M�W��  ߓ�n���� (���~�r���;�o�:����zNƱD;�鄍N�%6m�E���RYw	![?��M(0���w���z����1«��㫄��\/�^��}����Z��<CI��/D��*3�Z?��`$
�;�����PшZN�
���\�u7��\:�jg����&��&R���^��hę0~4f^��V����V���d.�;��-�~�
b��(I��rl�6i"�̹���][��~�d�2�����N�`E��K;�9G�l���Md�����F��ԘT'�`[KJ]�H��+%��<�}��C'u��"�{����V0- ��0c��vx�O�g�*k!�^`�(̧�TV���:�V[�>�%�4D㱑������e��!��>%ñ���$�u��	��}��C� ȵ ?�(U%�w%�w" ؒK�.LAa_d-ű�]�d�HE�r������.ǾЀY;@���/�ЙX�C�a��Ht���5�q4\1]XّC��R������\	�LLjx�"���Z�5DZ��آ�Q�^V~�o�Qf� "�N��DyK-��,��T���]�	�5��)���>�>U0�u����ُ�;��Q ^�eWx��Q:z�4 #ԃ�\�OK�z�8�s#��E��7�4)#i#��ήt��
g�q��s�o(#S�-$�#�Ty��Z%�΂5et�FC
i6���421���>��	d�������&)�K�dw�|g�t����H�a����%}��@�ݏ���S7��g:wc�s�A������w�t�F�z�Q������3.�t`��@��y���"D�Ig�˗I�;�S�z�* ����ݘ����ZB��4�t��w�P��;���ɩ&ڕ�Py�]$���&�"r,P%9 �=�q�
��Ɯ�G��]/)<K��K�)�+�6����Ǫ/��J�RZ@%��슷�7J����P���5X�M.nZ�=�d������9��E���í�<P����e���ʍ���Q-���{���>D7�(���e��z�� H��.l\~8����T�a�Æ�0��璀�3�>aD���zM<�߰����噩=������>0U!C F�@3y�䨂�{W�T����
�z��wi԰�m��� ��4F��2�3b��Z�v[=�)�80� f�b2"��R��9ӷ����BQ5���JC[�+�!�eAUL�_��)S�VMJ���&,VrSt�_U�xG���Z�{�^���}ưm���&b�y�^��Y�򜅃�@�7�"fK�I]�4���f�/(+޵C��E���:C�W���z�el�Ch�&�ԍV�3��Yΐ�w k����L���C�I
l���n�ڧ�d��M�^J���suI�� i���������>�x
o��&l/	[=�[�1�oz��X�&`:���.����������5�̭_ϋ�_ySU�)߹[8,��,���.���O���{��08*b!5T���'v�*�)3b.,�^(:��t��>���9�*����\��L�����O�d��U^W��ݨ9���� 	��0T�}��#�=>�
P��FD�_=���xG����W~�r2{��S�c93,NW\����)�僝1S_�������*X�%,�ph���m�x��l8:���Pķ���Bs�%8�zΤ�+�t�1~��EBDb�d�K /=����b��ȋ�睔�B~n��Ʌ_q�Y�ي����#��I�KF��� eN��R����<?ǣjW���J��������%����)��(�	�oD�����pZ�$h,o?��esY���Eȴ7�
��,�����w} ��~��&hNA����� ��t6b؆l��D������D㟣{ [z�	�FYŊ�������_� >��d��,���P���t�z+���K���J
 F�S�CZ=h�^�r.M�������Tx/�v���C�t��ɺ�\�����]1�-�zS(�pnokW;,���E>J/��#+^�^޵�	4��b��E���@�h��V�������|$�~���tz�i7�����D"m���VXf6�'�8���e:g/�ˢ�y9��YBX�T�I����c��.���3� ���[�	�аi�f�H�$�����ڹF��/��Y�Iͦ�-��7�X��@��miZ��L��tu��]{����i����2Z���N +i~�ǡ�$N�+n�V�$��O�)Y5�')�$j���P�� � �c�LsqQhQ,����O�G�S�+ݭwIxMB���sQ]:�>��M}�]g  ���vF��ByMh䦘c�N1[�:i7�?��`[m�S�Zܮ�����Z���R����)�|q<�]��Y�����@'��u��:T��\0[��z��cC�@Q�X��'ʺ5��;�Ji�y�u�}kn*m<�ۏ ]�\�p���a�#�lh�+���ip����Ϩ�����#T�04o܍��|������&p �BH����۝�-�-�/�G�ɲv���5)��[7���zH�v����E�UϮY8m��(�����s�C2�;>��]�e>��4�'������4ܱ"z�HM]Rs������Ԅ٦�[�"=Ǭ#:QR�ں�G�����&R��u�#�%&����ڬ�t߼��!�z`���]Y��>C��d0z|Dk��At7��rtP��� h{�RV�l|�䦕F��n�ʦ8qȷ�����, Ҥ�	5w���Y���d/�����Xw��^p�S+�P%��׫������k�f�$��ָ��=���oJ�����x�R6�h�Y�� ���b�f���u��V���7���tm1���.��g�q�os��7�c����)�9���,�C,��c5!l����
�,&�q���ED��� ;o��䅵�E���lZ�,��J]}�~��N$�c�"�6�g�ύܺ�j])ԝ�CSk�鲍�1� ���"|E`�p�?�[p���G��j���H/�|Nl�ln��J��B��Y�f�%fd��Icؓ����\��Pf@���l6�p{�U=���q!Zw���u5+��S5��Og�!�L�Ƭ��%�����)<��ح������8��A�l��Z���֣X�g!5���I*�SJi��~��ݬ�S��C�(1�*�('��7'�ot�@��"
w����(�"f4ڿf�GҶ��rg�d�����zN��k��~k���Rm�����Zt��q��t<@"O��}�mwQ9�I}�nX�ÅG��n����Z�egC�����D���;�v7jf����#x���b۫���4M3������P?D��D�z��w�ʓ��ͣt�ё.�n�{/���{*JtK��w������4^T�gϖ��r ���&}3��K�k] n�	��fx�a�����&.��4��< bck�p�.�� �����u�e�=�;k���2I���sN_������R����M����m�4����Ƴ��R��A�8��U@�A	k,�A�ʙ�JÕ�� ��|�mm�ݩN�8�"��zc�d����`Cc%g+���G� ���[<u�H5Ͳ�"���z<��:����0�L�=j��b#�QC�y��Z�M��W8F"iG7ᔾ�	C�y&Һ�V���٧-!�i���utd�'QӋ�ĶwM	�@�����N"uq�x��!�v��}��h#�ݾuA}c��e�8���/+�����:+�$PnIg�껃i�����e��ȔZ������\s  ���G �JYlŬ_�?s�3�?r4q$��͞��A> �a̜ D��Y]�c�+���B�ϣ,��
m�X������������:p�g��_�n�i���t��j%��n�7}�U��\èA��U�p��硎��w8�u�Bu�bU�p�l���V�}�����ҭ%;��Hr���߼��	$����ԙ��Gz-�� �bk��~����,�&f9�R�i�����-����q|KhYD�8JQ:�B!�=�[�ͿbЯz��Oܵh�wE����RĒ�^�Sd�|Ȅ����^��Z����_'P����-�u����r.�\��K�����MGe�H ��|����3���M'���%��$��>{-D� ���7�y>`��j͋�V̹� ˉ�][#���*؛�rq�>Ek)MN��ѷ>�j�o����q�������j�`b�����h���՟9L/+C�i��tG&�)*sO���,�s�%��?hI�Sޅ�5fOV�9�)�ie�񑕐%�U�\~�g�Õ�����_s!t7�2���{J������+'�:/���!&*���n�uNS��"�6������0��}T�� !��������Ƽo�3��;K>��:�E��R�C'�Gt�4s��qR�Q�Z�ov��J�kV���Tmd�G�	�q;V4�����V��m@׮��,M�`�]Z���+�_u{˚P�l��{Q��	�DϔC]�����M�D_�Ls�
�2<�k��?�b��m�=���<�k��fI�cN�ܜz|���9�)��Uw\��;�>!p�m�D�v��~�)iu�
�1�;�	icx� �1���H��[��s�MW-p{�fƕW�J ��z)X�����D�[�:�@�)�G��`�|�,�6�lMx��~���2Ԗ�*���Ə%��"S�,<cØ�D2�X9=���̀��hC�
�>�Q�	�{;�#==�#&��6����`�.|�-|����Ww�>��%��a`NY�B����h,9o�FEƩ�vnX}�~�p/��Ed���nB{���n!ˡ��C��ظ���,�Q���C�Jޭ�S�I��~�#Y��>��wqz��>-сm`���"m�m�i��ƫJ�n�k�}��&xk�t��=���3.ϫ)����[#|X�-�yj�b�.�7F���������i�b�@���>�:��RX
�`_������q�q,S�s2��PƟ�t�R�i�h��f�w�����K�k�j���|k��I��L��E]z��Hݣ�!FC TSlIC��O^ߣXFd�I�Ha��$�q��_'}���T�.i(s2J��q��᱕:1TV�5�q��;9����N����6�`w�m�|������΅-aZ���Өy�6��ϱk�`x��J�]\�o��l�K��5Әufh����(�N�����`Ԣ� 6�o�m�yf�i�[QeK�H�.1ܳ:�n��j��z�;
'N�]}��&�+zn��!Ꮪc���6#�p�_���U��\Z>>)�lC�� 0����dmBr�T��Sb#	�[�XS+�="c��-�_�Wx}M��b������]��5R�9p#�ȾS|=�]m��%L�q=k���+�B4}V6k}f��c�da�&����B���#4�3��_4��:�����!�
D���F�,�,��R�����=�7��b.ZG�-fㅆIz-�u�n8�t��m+z���%��۽�q��S��wa:���	�&c��V$od{�0�����Q>Ft�v����s���ܖ���:c�F{��j��7�*���ES�-Y^':o�[�}\K��4	/Ҷ�FNȤC�Z�A���qa�<��>�Ĝ���A()�l���5~��vԾ�k4)1�@����BzUq�*,���V��.��C�D0-凷S�ҫ�������҈��ꍵ�@�)��>��g*����An��a����C��-���>$f���[�T&��&Z!/0ێ$���/�3��h~3�#�<��r�-����cn�پ]nq�\�aE��)�Q�p|kt'���R��F��:-)j0e��,n���S=:��٣���xU	>B9�MTqSN�\(^�4`:#�ZY7^�`�[�Lِ���`2UҰ;�p�>�N�W���� ����������FA�Gմ})Q��ǳ��Z�$�[�S���~A�ҡ���V������5���ކ��Ҕ$�*��ƙ}d��էƤP���,&g�r͉M�"`�&�`�+��oj�kwzgv�T���������n�P��%��ӾY��pU�b���HO����r1�y2c���L�@9ʠe�v�Mv�s
s�t���ʘD����.�.�'P	&-�MSf v��
�X�ˤ��,��nh���!th�zwgE?#mt�������^�L��'��7����V&��Ū{8��|ZT��١3j����#?J"u7�G �I��3]}G�>��b��m�����Si��{��=�D��&3t����r�V�9AnS�r֒K����j�4�f�_�+6�'!�J�WHT�5��J�|�m>fg�Br3��3���6�n��#��ݑ1���Y������H��%o�)c��j����^�'���|<{tգ-��A�&��^���������U�v9��)#Ro�t��(�
ǅ�3��B�w�-��t�%4�t�^�T�3��?��*=|��t+�v`Iv�4��>`�R+ʟ6m��D��uk]�),�@�ˈ��re�UE�#����QG��UC�K����Uob̩7�;��������M�.�s����`_KU��Q�E�;���ku��5��'�n��1�;\�����?=��r~/Q?g�C�(#ͧ?���)�g�ُ��
I����\�;=�gh�1f�p)�]3w��v��o?��>9 1���p!:}�a��vp��1
Z�_�m,+��8X!��%����gc�%'C>�%��'��F����D�/Gs�sţ�V�/�׎C�O�ւ_��ρk7j�yp`:��;����Z�u�QJOOs���,75���wvh!?[������X�������[���M���pR�=��F��A�?����#�(EZ���Ysi	�P�
��~{7� v7��6H�gjS+�Օ�B߷��w�Pa)[���4���|��n���v�i�nn�]�pD�󉁴�u��o�xgH��M�`A�ђ��u�r��y�R�v=%t��ir�rnx��4�MQ�Ka^��a�������|�'T��g1�1yB/���^�o74�ĝ�G��7SsO �����dU��vp�\���B_h�b� YN ��9U�X�t~��`X֔C6�ɛ�5��Vv��tŸ�T���.�QX�8�9x���$�P�`K.if<"�D�g�-6�@��i�\ˆrgh�Sj�)4¿�U���Ru)��ڣ��2= ������m!$�`P2֙a>�f�����T�O0�D���R��d���o��x��><<`�@���s9֠O5b�w2
�I�h@' ��=9�A���m��ΰ�z�8� [�����c��U��~�x��$S�.	�[�f���֯�cN�0=�A�c����j�_ؗl8J"�6�c���.=�:kڀ/wEW.��@foY����`��2&U��.��M�z@�d
���w�-]>Ŀ��7N4�x|W'�G/>S��_�t����[��:�,�5v�@���_u0aT�-4+)3��S�͙���n�W��u� �b�w�=ϱ��F��������<�؉�>GypX�Ա������]���;sTsL��,�S��+ ���fx��=p��Ix��F��@�q,�i���g�1DJ�5�[�̍��`եV�#ٲ�;x
�����R
�(�>CcrŅ�W���q˺�Y�Խ>��� �C�)��E�ΞM�"�l�H���62D�����P��Xãy`�[��U���s���Ύ,l���۝_|F�50;9�~���x�hC��:p��(!��2�PJnn�B��0�|�lQ�Yq�R~!N�v���Pۄ�<��F>�6��!�cHka}���'����@y�~����0�����G������5�۝���]oG�c��8�)W-=���9"�S=w�����HцizI�i�(�2��ҢY$�.8�g�y4��#�y�Ȣ�l�m�t��c
������#H��2i��u���$so֚H3t��nK�W���dt��)�?��Ĉ6�O�}��?\skʔ�7���b�
�7ǆ�'_����,c8�d��Ʃ�O���QT���u�Ed��M��Z��8`έ֘&��?& F��1]-��{�?�GW��X?����`ж�oc:�q#Z��ɀ�, ����7m	>W%(����S�b��0G��o��	ißnnA�e��I�B	"��"�,-���y=ƚ����*Z�#[©d^�[$�bh$��V9�Je��2�e>��2|�����y�r�޴Ș�:�xa�N��L���i01ɝ�ݩ�/ҡM���d��s@4�����:I��{�x��\�=�V�ᶑ�7^��GZ��z*���7^ ����w�?13
G�oQV����l��{���c+�_�)�!�Md��� �e���f<Pz��T�)�����R���~:5�N�V����Xכr�O$H���jO�ѣ��Э1�!6l�g���##���~�g�a���Q�u �r���)�*��/�i{Qa�1l��6KN��u�����p�-���V㜩��6��U%��c���6�4�B��RVҵR@^f��`�$��7�*�Hw���x�d'4�����)��x���i��?��EwJ��;�3�G/4v�M��@[�r���N��'�ox��_[k�k_!Y�~�w�BB3A��Og�ժz���L����zg��9p� R-��hB]�jia��t�Ϲ��HU�Ϝ���-�H�1.�o,,U�!<|d�'u��J!.����t�J��]]�0��WS��Z^��P�dxҍ,x�bt�jd%�ݥEq虓۸V-D>Ĝ�+N=5WN�q B���c@�U#�<��gk���A�f� ���6a�μa��F�\ߗ�{}Q�"$�U7�U�ΰ��7�����&���e�懍]��5чɶ,k�G�;ҧރ1�th1�F������u��W8�qUï!�+�-�!Y��V�*)�U����4&�����}��ȏ�V���P�T�Ee^!@\�@V�p���E�M�����#�nJ�dTl�SP��e��j�{��x�do�ߩ�6��8Vj��5zk�'�r�,����ƃo�xC�}2�AӲn#0R�k�^w�+�3�wM�c���!�BL���T.8�T��ӆ���U(�L��b�*J���]I'Ĳ:�m�ׄ	���g��>�^s�0�ݡg5�'��7��y�u!�A����HH��4؅~<�<���(�v����t��3���F���{�	!!+ؔ����ȗC�1��4��wMN����4�jQr���1.�x�V�w��Y�)0fb6��M�'5�e��k��ZM=?����Sӿ=tH�X���]k�����Ŏ.����2�Y��J�.���d
��8����z���->'� L���Mk�Vor�tNc��KC�)�AZ��6n�	:8�H�R�YB!��SͿ���"���Zn��HQs
�@/Y_%�{���؎Ѽp]���Ϙ�
U����@9۫l^X*��?�4k:�C��+��Z�J�T��r)��-RE[�0,�ܭ��F�
t�o*'mX7��j��{f紼 ��o� >�����U2N%)���<I��R�
�0[|�m�L6�3Y��-��X�T����u�\g�������;��$,�I��J�.�zox�6R�<%}:Ul���ú
5$������8)2�X*6����⓸�$O?@tɵ����w�q��_�r9�f$�:]��t�����`K��
/��Xή��
����Q�lwGԖZ�}[WF���%!��\�e��M�W����O%��Dq�������EF���:m�m�XP�,)1\*�ǥ����*R;^_V��@9�� #y�H�hZu���I�,(�g�=ٍ�0˳���-��'~�����k�	���cɥ ^4譏�Z�z���`�w:���� D���Eu���V4M�,!M�>��}8o��&rN{�˴�N(D���=�N����v��n�Pi��ǅ62(b������eǓ�xb�r'
**�h��+J���\Icbt����5�+H�6ki[�|�S3�[c�����IU�X7)Ӥ/��s���	6���f�����?�#u�G��P�'d��Zg-#,���/\k9����6��o�V�=W����n�iҌ�yw�[�t,"��4�`>]��LZ�8,��!{��?	�C�#&a�Xq�������	~����� ���J�aQ����n}kX�)�g8���N"��}��$(�uV�vD���yٚ䱕���M�:q_��Os��8a�,��(��2�&��ѥ����j}ê������Op�+�GiP.�ɝ�y�1��p���l�b��E���U�FKUNJ��t썽J�ϓW��Hj�J�]H`�L���^�ł���2�	��*���i�W�ڸ��ϩ���Ɔ����s�@�;cY*��,S���\�p���k�������@�H�4����1��l��\�7�4��"8
�5�c�����eZ�b�+�v�֨��F�g������)B���{D�lj��Xy<�]񌽷�b�Vl�3A�5cc���7\��9kyrP����ol#�Wm�.{#^���	��s�
]w,Uy�Ā����������;[���|H��Y�>A��5#��e
zm���F�=���ok�U%z�{ƕ����*���$ݫ��|�N��m`�W
���q#�����&����I0K:��X�,�2�0t_�[m̣4kj��I��A�f�����ϩ�R3����S��ۄ�%q6`#j�٢���j�E�l|�5������u������n.��*�Ud�|�_`e/�Di�R��7�R���j����x��?}��k㚋wty?vO�d��o�����ࠊ��K���{5���\}�0�[�Ď>5���e܃2	�W�,���y�FAϧ-)W�uZ��*�~��1�δ�	b��������?P�=��lM��v�?�bb�i��G��_ߺp���c&��B5��$���åV��F�\�I�k �t�!�l���8�K���ga�v9.<*��S�6��#��lhw�P�N�t�)�m ~4��:�4��L[.�	>��������s~�8��x�<��}\����v��~�a��~���?�2Q���2Ǧ2�q�e�zE;���?1s3�����.��3F�C�uO�JO��b�� �+lX3�~��������M��0�RZl�˴��X���[z՜��/ȣ��֘�{�G���� �ʑݧ*����[�۠R�u��aԁ��#�cA��<&�W��>ȴ���Qȝ3�ב������ ���y4�a}�$/�ğ�k6��>R]�i��3~H1�{X���&�1���sx��T�$�h�a4H��J��+u2��+���@�2�Hq�~X�ܚf|������3� ְޔ"~��P�55���� hv�`21���o;pr�d�PT���� �`����V�祳��c�T/8��qMFb~p�d�����0����>�'���n�#�5<.�ʤ@k�P�LpLl�[�}K���d���MJ��#�x��0��H�[�kT�~hj�@4\dc���Sډ���K�Nݑ��\������K/Z	Trvs��ь�ĵ�i���u{_f�
ٳ[O��b���ɬ ��oz��Y|�l�8�I���hDR�璧j� q��U�����V���iY�ZuN�.�q��31$�8��<�!0�i��*d�	��e�D�я?o�ڐ�3V| Z	s3�n~�V�)�5��z>��W�\�q��@�c<c�P9�f� p�� >h'ѱOfP�.s/P��a�N�� pg]K�W�N��6g9��w���k�$���nn��:�z��~8-y����V-,����! jO��+k��d�Jģ�GD��n[
X�;�}5��I-#D��I��o<w�d���2�k���e�&$�|��\cE	�K�ȿ� ��7\�~�q����У��߾�VU~|'���D����hǐ��\L�-g��c4�[��{�02�W?ÿ�a�^ME-��_��ƕ1,���Ξm�� ~#m[R�}?\OL~㚰�e�Ia܋�T�doIu�+�&�}Yz�t�����>��"��*�Zp���j�"�U���������k��g㛞I��xs69�ZK�ZC�P�_Хfo��Jh_�rb����hdH�N��l}��?܅n�	E5�ɇ''��RÚ����2 )�>Qc�_#D�=��e9��@z`qc�X��i�'���v u<�'��zs��uN�y %T�!���2���0xh�A|�D��
Y���ݚ��z�O�1����r�ǩq`�n��'�t�E#��B "��3
�VN&i�w�a�^w�`��O�G���~C�g�)���Ks��Wa�bv�^�j�� �>1�b��~rB�˄H��T��/���@���}@�)�B0���~���䕙�Ͼi]��~T0��/�c����?H��ג��yV���Ct����; ����z*��ΰv�1{C��w�-���F��ֿu�h����������{4�χ`��ą\v,=z�%Y��Kec���f��p�!��(�w.�.>�M�`J���L�RCD��.ߘ}��,����a����`�@���j^W�E7��#��e��Sa��!ż0�{�THkHU�D��+mL$���_�яé�����x��mS���ٺ̯L׻w�s�Y��-��h��m�N�����|"�@uj�_c���weH��(u*�t,դ7� ��_��S����顚�p*��?I1B�N��ӮV8!��F�@��=����̤�I�t>��{.��K(ȯ�`�6d��!T�; ��ݣARQ�/�x���?�3����I[$���e�/w�e\c����z�[^b� X��<�&�>�=��-{�HV�U�c(#7���Ϥ�"�[saU:��6����FWky��@^�z��T S����o��%j�	��fV1 Τ%����U�Y���X���٦4��J�$���0���Ϣ0�p���.�����:�	���e��P�ĵ�, �ʨ��]��}a작�{��C�Fp~_Md��4�S��+x'�>xb�P݄p�;����wdC.%�P���0T��� ���r
/��>^�� �\�t��P],r�Z�9��\��}dUP�X�l��>f���~�ß �j�QF$���@!ad6�kگ��)��8<�3^	��.Ŀ�ޯ�[Mz��۳C�'�Y47�/��.~�������r�x�/�E�����f��l����|�6�
�;$슀�c�`	��r�ˍg�9X�&W}�#���`5�z���ˌW�:�BB�Y|�L-�[�	<q���=t�����0��W�X�*
�B\�i=G*�G�'{�*!U`�3 �+$��'�b~"B���(�Gg�(X���bt��?�:���K��$�3-_'Րu{�^�g�G����?N� e�G��e&��Z�g�l�] �3��U�8�$�
=ſ5��A�G2-�i�	����,�|� _V8���C�1��7nt�v\��DH��Ew���&
��A��'�KK��?���s� HI@0:7�+���PQU[��è�LL����V�+P�n|���
\����f5Q�a��߁D��ӱ�^�0Hk���B5D��^�M��F�2��	����F��حbT�6�������m��?{g`�b�[������W���V�	����;&����'{�ӲOr�� ���&�\�!#����MA�����2\i�A���f?I7B����������|Ee�;/��GO�!�~̳~A���5>r�ës^V� �??p�䟓#��Ǚ_��������`�.��~E��G���|�\����pC�p�R�Ԫš�֛z�����Y����۰�0v�  ���ea"�X>M �N�Ԑ��R_�`(y���G�Ơ��)B�É�4C��,ҁ���v>�74��r�aa�-��i�y)����f��xUGŊ7�]�1�0�����%�%p��%0�#��A�>J���?�8����XU�⨪k���8>�a�+��*�]R�G��YC���5z�+��~Ts��~�H�Gt��7ȧ?Y��ӡ�_N��ڥh�� �o)+���ي���Ɣ�7^�Td�����?��Uŷd�=K�۰�p
=�1��x2�Y_�m PD�I.��Yl��,,L��ϋr�<��ƲB����vq:�7��Diʪc�ˋ�du � 5b�D�L�*��/3i �i���u�.j�(��:k�����p���a���Ѩ���Gy$�-}Bߨ��Wv?��ڃ����O��,�p�k�#�7��m�����G�L����u�m��u$<:U�2�Q 2V��k<��o��밓z������T�P`�����P�Q�c����$�k�[�c�(]��D�E�؈��mPG7�b4(`4#H��*^�����eJ:,|�P��2w8��r���t(���Px{�w�K�5��=��gQ��n�}!_1(d������nX�����c�'�'V
���
�lD�f��A̰3K.��(%ш*gV����+��t�(�U^Q��p��lr����;�`�1�'��'�cPp&���)��g~>�s��<�XB�O����}ʋ�Ѓm9����7̀�0���`���O,!u�/�?�!cJܬ?�ic�%w�F�86h��/p��:2 ƹɭR��D�ò=���>�o���q��|�>ˢ�������~��Jf�9����}/ʩcs#LA���H2+�D�Q���#O������.kWϫE>��jJ1��N��U���ۀ��#��?��!������¡'G_���RE��{����f]�Ļ�>R�;
��4���g���o���z���{L�;������X.��P9��c[���� ��$����6L��.�eE�%����

�LY<�Oa.��C������h]
���%-��~k~4N	DI	���:�f�ˌ$u�i�дb��l6�r�ۻ(�A5J"ʺ������?�*�(��Et}�gdM�� Ɯ�B#�>0Eŋ<G�LH,m��	H��R/\� �κ�w���/��l�ה�?X��+�;;)�p�٫�η�rEɃd�h9�6˦�؏TRD�::���f{!�t(�Cj��@݃1-�l�q��nE�a}b�MI��*:q��)�M�¹�:N0@�@�k�����R�f�Y��B���Ǆ�6�=^^��#�V���DWh#8C�T���B��h5�떣]	W��e��2�(ն���[���6���(����[	6��s-s~}B�쉝�$>���^�:����[�F�ˬ���M��q"[�G*_TIi�<�!{;7�.�P$��h�����IK�#X�����Lv���K9��h}�XIHT��/U,!�Q��	�<Uov7�@�8���*ns\��E��|�Pn�t�]</m\�海o��RKE��"Td��n0)��L�۸'ώ~gq@2v���:i�6a%������I�C��sJ�(�^����o���C㩇�F�̛߲Y�����X(G�Z���H[o�5Z�G_So׉��$
��+�Pe|��x�Y>�@Œn�9ほb$Ј%�$#�bq�8 -�.g�%2F���i�䏮l����U�2+��^�j��R��� |�`�^�)���o6���~H.ԯ�ה	�y([������O��߃��ƛ%y�hc�.T�_p馬�ߕjh?�`�>��.Ǳlp�*䴷���%���=�����)/~y��;�i�O'��c`��R��U��A51SD"�O��#=����b�֒	��ߘ�Uu�D&��ÍɁ�w0�CZ��h��Z�pmË6b�p|E��&�h䖇���,���>נ�}G�Etz�B�s�H�\�V�$��n����K�l�䝴\����H8
���~��G�6ET6���y��J�8;�F���C��)D��:H��Y���L:��Xj\���z)?̑N�=-L5���ټ����8N�
U�m�J�=��V+,_���A��{�;�w�V���%x��UB�KI󨥖��h���ޥ��^a!��ꤜF)���vD��|�W!j��b�lG5����94�оҜ������(�����)�y�F��:A���yB�r� {��IyZ7�rK϶��?4@o�ɉ�q�v�9�!]="C��߇p_���3U��]���ݼ
GdX��pl/c�p����9�і��'W�v�k�ݿ�%��!u��?�O�+	'��l?a�XCH�	�y�P���i�z��(H����R!�ܭV"�f%�;����Y��{R�`+)�#�`IM`;Z���Dوh��q��_��W���1 ��cK�}�BOBRź>_�s���؈p�R��`��)z�2��g�a�j�@��b	���[�s�kQ���B���W��%�_@uC�����#��yac�6Ӻ�``�AA$��WzZ��<�<��O=[����tK쬋6��[E��%{��\9��dԆ�[#��U�
d�&����z��7@��C^�4㸯+�X�I
�Uu��lv���9#�h��?����io�+�Tqj��3Y��A�X%g�j�H��\h.��a�I�[��|�����h�J���e��VwWt,wPN�.lz�{��rd�F����0��ZF�VG�]�S���C��dmw�����kw�1�[�
�?�Fh�W��"I� T�ϝ/ũ�����ܲ�$r�ؓ��� �Z!Y���ΈWf�x>6/S�NX�46�޺^(w� Y���)Gp��)j3��+\��K{C~�dS�����x"_�ka��Ş�s��&�n/�^m��V)�6�D|��f�R!�Ă�L��R��b�؜�X��F݈1B��W���cG�d;>�����>)��g^�5Kt���.��!��vN]\���!��(0��[���&��yY���(����k����������y�#�^c!���ȉ�3��S)8Oۚ�q�_:I�~&j\����f�D�d2JW5
���U%� �-�s��������_�w�|׌�a]�˒Df�D��$�.4�-"�}��n�I��"m>�	#�ڰZ5z�[�Qi`cD]Zj&R���� D����ز4�e��dB�����X�Q�����X ��JB��{n^T���S���)u�b&��l����+~Wn�r��ϧ(�W�9���r�WF��b�8�Y$pY�q��1��kz�%`w����t�ĳ�y��A
��VN�k*}��B���;A"A����Gqɦ\����P��^�k��ч�*Jl�����H��0�(ع�DRv-MȚ#��8)s�Un���GU�jt��h����G�󔀙�w̬q����dI�O8A?�Kx0hkR~;&�֞Glֿ�TaWFvL� �mi�Թ|�[�)�^�����=��d ��6�0��w�eZQ:��޲��@��P�D�F~���Fr���_�"�f��v��͖C��>�O�, H�W�c��He?+�|o��
Jn>lT!FHa���/5�EIC����hi�.�y� <@D��N�c��� �{Φ��H9���c��#Cv�s,�Yb��!�ZQ��K`V���p�vu��#���Y�E{s�����<bA��:CL�j��V>�<n*/L�Z�㗊E��8i�?���F8�kYݬl8ZY쐘>�$���(U�4��`Wa��?��G�aw� �rҷ�&/<Ñ\� � Ψ��P�)Ta�;a1�:|͕���%0�:�ys��g���I���ՠ��$a�#|���[@TT�]���T�v^���sa� �ؔZF�����&���y����F�zo���\
~��N��!��0���*J��G܀U�n�pw��6�� A.�̭>�?��QM��unL��һ����oa��ҩk%%�Pq(�צz�C���L��|�Au5*�c2�CHZ��Y��x���m�R�4KvW�TyTz��T��u¸�ȋĉ�����H5����RI�,�9�Y$��g��n���h�K*�6��%�5��+5�G�w���aSS�"�ذ��G��Y"*G�$���7@,����� {�3��v��ް{�I0���+�0�6t�M�Jn.�a�v�2��t�^,���5�T�Uf��c��[����E���:�rQ�Ls�c�����h�Y���Д�t��}4�{,��o��g���6k�۩	�&2��x�U�'�zT���0t��%(;�a�\-�'f���' '��(3]�ki.������b�[ �3��m������thX���_��-���	�ҵ5:�g�h؂�^Q����2B�<#9F�el뉘5�Q�2�3\�A"������)V6���R���l��i��H����uL�I~��;"��3[K��C���E[J���n�'{�;�:[8^����*���Ћv(�A��$lS�ؚ���'SU����Z�+�%��&H܂�4,u�O�e�fvo�PE�V��]���Pۍ_�ze��"���z��ٗ��E���o��T��|?���A���ݤ��xiNڦ��<9�{g�<�zD�3��Y����WDG���V��G�L�Kn�P0�~���*X��f����� �r�[/�K-�x<�x΁�"m�Iȷ��y�h���PV���:T��iaQP�n�t���P�-�'�
����ʶ�-ڍ(�_�?�j��
�;n[�x��E=MTL���~{�_K��r����%�\=�G�^�Z�>R{
�H����L�r�p:o��h����'S򬠽hn� 
�d��	��pGb�W���] ����U�'/D��(񥂛�!��&P����	�N8��$�f�*M�z�֥Ty�������Y|��u2c{l����s��Lnw�
��n�$��"F]O<�$���$��gZ����5Q���9�s���&�bp�p1{[3�V������y�W_���ʳba�K�� �3А�h�����;�4U|ހ�n�tV�����+$�i��B�s�~����?�G@t�bQ��R�r�Y�I�c��Ku�"��¸�O&�e����)bd_ >�q��������N��� ��^-�w�ò{6�
�������\3��ݕ�j����qg  Ym�f�Ȕ�o�;�T̾�+��i��@H+T31:����I���<��ݥPGwI$���ς�6҇��)�?畟����˯����� �-ĉ�|�3u)N�B )��$�v�q�	�Z���d�2F �<5���f�*0�|�n;�i��a���L��M�����橛P�y&u��Rp�*0Ȩp�ݱƵ����ʳ��+iyG%���$�Ĝ�Z��ә�u�+��&9��KЍ؉���Fw%!�0 ��������O�����s�-;�V|R��  �m0��?ZW�"��mhE��VnL �nЫ�3H05sz��p���}�X�8�^0��N}��)�Z>���a���mI�Q�B�I��m&����-�,k�0����}�b�Ъ��4