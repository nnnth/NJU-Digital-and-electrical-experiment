��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��op"~Ϯ�!Z�	�����0�q�(�q�S%�z�(Ha7y����2�m�B2d/{����8<T%7]���[L�P�ٌ����7;6��M���6���}���0��>q҂��/'�<����	��_��:h#pǻ�1g!/e��(w2&Я��@��ݕ��"��Zh����\�N9%���#����폵)?{��d�����U/R�毩V2*=%��:��r��:�қ����&f?�@��e�R��n��z�o	�ܸj����z�������U�ިq�{=#tH�(��7��<3�ae�����۹e�� R���p�oO��!�h���sxiZ��E֘�s5UL���B7J��
��3�|�i-+��VQ{�Y�+*i���9��'���/f�fL9�9S�Q�t�$-{'Ͼ�)�o>��ĂUc
��0FJ�B�;�ࣖ�SĹ��w0�F�SL�<�&�ī 	C��.������@�Rn�� i�.ux�m�2�1�����rdpD��n�?7�t�<�Ж'�~Jt�$kf� �4�[i�??�աA�@��c�<�f�΃/ڏ���1�	3Dr�	���.=� Is�7���A⾘�p�#i*+���k��� �9̥����(��;�>�*�T��}.�����*P�k<����(�L��:�pS׶o��ˀ0�[�
�J�0�g�4���a�3�宵Me��)?J��
b�,%N�:kU���al�"v��<On�ѓJF�̘l{���)8d+೬�L|.��!��!x�J��_�Ԯ� oW�^U9	'FG�xx+2mQ���Y�A[�(3Z}�����HSHd6��R�5�+��;7�H��\)����Z{_/aU}~";	�ԩ�w��GM|��DD��x�H��t%�^��#q"~�6������"aM��d�p��<L8��f����6���4%���Д"tFX��F�p�#3�@��bpW����u�*Й' �Kȁ��*��'���0��~ݒsoi,��s�an�+w���r��!��J��Q)�n�q�0I�)iV�wФ���W\�m��x�SI_�vo�TX�,�h��9�̕�R�>ٽ���[�ю��?.E�
��߷V�oQ��G6� ��l�`�j�Ӧ4r��j�ΰ�G��>g�~boV;���j#�NN��*�K��qD]��t^�y�d�[�$)Y���d]Ba��yf�>6s��Ƿj��O��x�gZ�P�L:�	����c�� �8��
W���t_�X�� ����c�AF��#gB���|8 
�YY�;��jD���hT�7I�"P'b���x)b�[���G�k?�W����pE�ȁ3Iz1�w������o椪?�\���J�%'�Y ���'���WRbk]\3�0�B=�e��/?���^��m9�������v��A-��y�D��t{���%�d��1���qu��5�/�
�<������C��S�Q[�I-�y�j�r@A��YB�����sV�/ �F5F�(rd�(e��O6����3�W%q-Ġ���p$��mAʢ�c#����1Z,M�3�,�+�g�����c
ruK�jލ���t�7�"�p�9�x��L��"��H����5p�i*\-�����͉fu��be�h)���	!
�_���S���5�)��r�ފ)���&9����H��?��@枽�f�:gaKb�㛵-|7��XT��T�iU|p3�N�V���(%EZ�����SF�����R
d�ȚC��q��f����?���-=�S;�L�z�J��A�ʇjw�� aV��̚C��L���]<���TP{���(1:�O���ꌌ͵����Sd���ItL�̨��Y�����A�`R3Ѵ�Բ�gt�(! ��������Uf�d����b������_��9�e�V�*�!Y���=�I,����z����ψ�ڨϧB+fEoE����hyL�Z�@���Y���~h=�y����$��L����D(;�ٍ� �M�(��P���y�l��c�
��؛=J�D
�j���7+N��fD�h�f~���y��A��v%���;o�6�k]Z�Ŧ��*�E�NNÕ/����i@�0nb}A���4*��q̔;�����3r���
>�F6��Eɸz&,��j;N�2���!L����&91�����Ox�)oJ@��"x�fY�-c-�ik���:�}�ى���/�q��u���\!
?Z��T��or|�Lu���)��}J�]�IVVwײ��1�㺼Q~*20��9 h^>�y�#ا��vU��yp*��ٰ�`�LP8�;N�p�@����ĺ��$3��6Rr\����${�Y�Z���ܞ)���.�aTӻ�+�@�T`��� 8��֊+������?�Y��o����/��(��O��#]t�}B�s�K@v����eE���I���o��0օ�$��� fV��*���%��R�'E�(�ғ�vݾ̽���L�"C��4vBR�K�P���N�G��-��V�����O���j��7�O��u\��m�D�!�tY���_u@��L��Oy�s ��낏����D����/E���u�hH}��\:�K���oq�/�l�ڈ���5��9��QL�7>.~��淧���8n��#�O��I6��w^�B�p+���*_���Q~"�g�_�~s�D�|���*;�rHO#@�ۢ��F$�x��;�[��&�/�|'������]w����%E��6E]Lb�l����$����:6,��,:���D��V-���~帬�ʻ�Nsz����cu�^����Fa`���]�|;G�〥��W�C�:;��,��$�7�/Af�*Ar�.�X����7�!;�T�j�VN!�*���|L6w�2��L���#�`b�>�
�[nB��W4h�͡����UU
 a%<�x��*��>��Z�8�Q�~�P�
�Od�O�4x�Tf�s^b�:�M9 �f�P��\ h1��9;Z�l���E�n���X�
L�v�b֥f�~ɬ�^⎪�T%33`�O巰3^		����E^�}�Q[�8|Ne������|�;� ���G�t��u��&u��U�����<À���%���v�@�ԩ�?�(�{�4���M� ��sq�[�z>4�ocM<��w��E����� �MN�v{�_�	�r�kUt֊��[��|�Z9Ρ�Bz_�mJZ�6���t~�����QY�����,ug����f�&ƿ�Gg����	iZ��mY�YH=q��Hp9(ói��M)����^p� nl�D�,Cm[m9���&v��6�a'̟���^P��/�Bޣ��tN��r�H�1�s`(k|��&�7��'=4���>��MBĔ�]���w�r�i:AE�EQDli�i�`J;z!M�O4�К�@#^҄Į��rdB����1�v��P��8������J���M��'倯��owUNs�$B��Q먺���������?/��  By�~��im�#����n6q:��w�_1�̙Ї��h=ٸN���B���0k�pǣ7���iH]B5�����;NqJz�g���0�*��&h��NRˀ�F�`�TpB �j��%9.��X�����������Nt[�o�2�P�!�'o��h�-��*s�Edk<��7�������2΂u��ϛx �Q�YxB�h�G�z0��5�0T��b�� �OyHr���}i�0clg��y��uب/�	��4�b��C�t��5wS;�cwl)�MnD���k�zhdq����|�P�3b�i~�~Ly(O�]�P#3���2�px�:�����TSIt�ᗤ))���4�m�9۷k7����S�l��(\�SҐf1�E���J͔=�f��8I���BsP�2�*��;�P�g�0l'�:m�r��'Z.פ�GH��ힷ�p��a��zR����%�n2���Qذ:q���!�����5cn��'b!P�P�g��1*�+8�T�fC�ܤ�ڿ�.'i&���yߨ�r	��@����ܾ�I�(TN�r����Vw@�Ж(���f��a
vS�V� ؝=t��/���py�'�+
Sz7լ�ŏK�{�X��6�>� �T@��+i�#�a�;L�AP8�hQ̿�T�w-acz��%^]>��yR�̬j̯�A`��%��[䝫v�R":㋖\��%8��"�2�C�`�!�=��K	������x0����<������X���94mL�;J�vw��n���'
3�=�ndn$�����8��OʷD���|H��fFX����@��a��!grN��8�J���,X0��Ki���ؾ�,vS|P�6C��+jR��L�c!�c/*�����G�Cu�8�9�Ι� �A�E=�m�{/���i��^k~s�K���Ix~K�=��V�2)�p'G�z�8�ܟ�(AIcl�0-���L��JX_Y���XY�Y�i<�O�:gV�l�ۏY>�?yt�rIj�Q�F����V�W���l�]c%I��ķ�i�lu�� W� �4S�j]�w���`E��'�A%J�����(�[�E��} �H��FG٪`#��G��_ �b������J���[gV�b}��{G� |�,iC��e��� ����"�go��-��~�ES��ݮ F�[�����\A	c��MO˓���>ڧ9��XŽ"�U�_�R��.�jOXJSm�C��& ���o4eLk���Tz���^��lt�q� J39���4���@!�g�i���a'�j"����ٲz?%)Ҙ����H�x7�Z���J���Yrd҃n�����E�ݥ�~�<jD����M�����O�#��F�b���+6+��e�m��g�a�A�3:�
�I�gL+x7�rQ��E��������󧕤!Uw�Esc%�=��,I�4Y= (����x�q�_	F���,T}�'�֛���J[\��VO_���G8�u� ��u���0`Z;�����dFڤ�<�g��4��ދh�f@���9��`��i����k&�(y�T@E�nf/V�C�F*�Q�·���t����p/�p���F������	��6VkwfH� �\˫��\�T/�yk�o3Lۆ2�zw�lf���� 
=G(�!�}��ƾp`��9͞���wR�C�,
CB>_nOL�`�bhh̠��VTh=+1��s���}���R!g~3��3}#���	��&�X��C���oN~p��Ϯ?���C�"��S�y�l�3�� ��ؖ��(�F�,��@_[�~<?V��l�����U>�PG豯�)K~ô4Qo�'��f��^o?hu(|M�`Z��]�)���-cU�>�S�� '� �q�Q�$c=�8(�O		�G��"��Ҿ�,[J��:h& �m|pDd����JWȶ�4����>�Vާ룎�ܪ�Y�������v���:������(1�EƑo�Do�'to����<��\�Ff��Fk#"����<-<�aʕ�r���#���
n,J���a�A���Oyoٯ���'����l��+�;7�4z5��z?�"��=�(3d0�%F#�zw�'��[�Wi�G������5�9B����)��3���/�M���Zl6*��&E+򪇽��q�J�������`Yr\��YI�y��G��& C�o��C��Q��
P��k����*o�G��5�^rѯ��w�晡�0?%M��w�2Զ�V>��K���hu�|�'����$T~c��^@�m�
_�}�Uv	'���$k������?N���@��G�N�Q���M[$��
l�b���gT35�e8��Y��׾�%���H�_T=:���HVP�(���y2����Q��p��b��UJ�]� ����W̲�-i�}8���
r-7bXVT;kĭ�1�x%�/�w�y\��{q��= ?L#�XS���� �B�Z^��-�c�ka-#�/�Q�ր�����-R[R�Znx�y�}�\�K�l��6�ٻ�-�c�w�X�c��$r؂hf��PCzt�T���-i�_{���Ao��%9^)Y2ɻJ�A�x��EC�ق%V��~v��z�f�d�K��~@�(G��\�U���p��?Hg���=�9�-x'�����0�Dd�����
Y��'�A|y?��:�6�����-x׉��h�m�������>�]1��Y�\;{5k��Ӯ��J�9HH�E�M΅�P��;��\�O��jo{�� ��Gѥ��K`:y���d+�i��*?�^1�ӏI�ǜ'ID�nk����$��H�������,��yh�X���pGᗸ�
����D�r3�;|@O��ՅV�K�G�����o�h�n�^0L������P��uwI��y����oNEh[�����U���ceUAd7dy���֠N�Jq���)'N�
1Nb0�x; 43����}��y����A�����������w�y�y� �z��{s���Y�	�����M噕�,�$�p�B�o�8�"���Zb4i�&ɘ�IGD�@G�P{��@9�[d$�� �ўWB_�:7ׅ�}*�%��W�YW����u��k�¥��lIr�`!^U�Z�46�aQq��yZ�ч?|O>#��˰�Ъ�u���}g����)�I�UahB	���n���l�q�ië�y��C�Y0 v=V��.sz��I�΁{�G�[��G��qK�*ǴJ�}I@���R��AȮ�)[mNn�g�.���0"�|��S;Bc� ˶'[a37[��{�Ru�?���L�r!/R��d�f���.�H���Ь�b�6�U�-hb���f'&�4�fu'h�8 ��/�߿}��,��X�Gk�G2�`�e�U���~�����s-�p�����|�/�S�;�`O+5`7�0���ӂ�ڟ:mֽ�aZl�\��/���^mW����e���0e��31,�)��W����Վ�洈����kF�����WQ�g	%�x�c=�T۫z)���������P99ص�u#��O�O�K����3}����_c�ȕ�g��Q�[#����1�A���I5V�4��_���] ��[eB��	��b;IN�kq�=���d��ĠD�nS�|��K�n6}*��좨����Q��ŝ2j���%���ɧ���ME�Z��mF���ۢ��9'���aƱ��n���$`�>�Ձ�Й�BV-<�|	�S�7[�f.Y ��N&�D2�Р�1�z�$[D�`|p�.H�<1s=I^��blq'�В�v�Y�����SЬ�~<�3Zg�ʑ�.��fl}̫���Bk5���6��."�L�p��؂e��S/{��Fn��5�J�X��,����A��y��U��,�urS���'�T.i��ޖ��/HͰ�-�ұ�:����n�~t�h��t@~���PRcq-��G�53��>t�tƛ��7���|���	Ƣ�m��3�&��Fo�^"����;z9)y��P��!�;��9h�YS붂dw��h8�ҙ���EEA}��B�`l�o�{|��إU�R�Q�atO2"0Β��y����'l'�H*�[�>$vVqC��aO���I�/�,~�F�'W}jj;*�;�x����{`ԯ�w#~�8?��qh� �̽�
~W�(�}��ܻ�O藽4�暿@�����R��w����QA���|�$�����nX1��<�~F���ʶ�]��qvف��V���LR�@�!0d���br�/��ߍ=0�k9�ʞe$ ���G��In18�%U�w�6�T
�^�r�,:��_V�9��҈��k7/��HM�]NQwʰJ1���M �_³D�M=�.�s�g��'+�Ԝ���M5�[0$UO�X�\M�߾XTR%&CY�M��/$
���g�g�.���6(0F�M$1�����*�#x�7���!��>�\�I��� \�'���i��nspf �����U��J �M��>�2��d��&k�@\PZ,�1WlϦ�X!Xj=ae���2i��_��Nde��wj�	���8�G�W�<>���+;A�97�|�,�4Q��I�.�G8�Η#!����?���-�9�y�=�u��q�B��:T�ΰt�1U�$v_���$int@�ƤH�%6�3��G���ݸ�D�;t��!D�BZ�,�Ҽݠ+1�i\�g$q�Q����qp>~J}%������"=R��_��%ux����C��W��6�;1�Ddˌ!_�vS���S�Ě�ץ�?��OA�ħf�
{V8xBe���Y4��j��9l�A?lb��V=u!%�Pv~!U���)�*�t/4%|��)�L�4̵�Z��%��R�B�x~}��ԻL������!��f�=I?Py �_W��%�����誵�ŕ�~��*��-Fd�����c4�Jb�n6q����df2����%D�J���j�X��V&�l��U�/�p+�Xo#�t�ۭ���DGf֎��B��E{Q�X̛�:B@	��NW�O��Z���f�$'�F�c�r6��z�WH7!���,�\�������F�����q�I׊�,��֬K��&s��W����ȉ�;d��[�� ��*��[�M�f�}��%���jcU�o~�js�H��%�RlEst�`��Hm<_K���q�=k�c;���gO��� 2�Z ޤ<�w�t����H	ŷma��b,m8���m�����r�\��8J���])��Z5�1���-m�ı��)����7v��������6s���**��j������*���������yZ�]u"dtb�����Ia�qG��o�q�-����^�/��{��UCԼ�ʅ�(�}�&J�J��0��D�j<���T0l,{��-�*�g�u}�����e��w�s#�_�l��g�~��]�U"^D�&n<�Ⱦg6�����e��ݻ�P-8a�Đ��<E�i�#]���|7��5���u��#_o�I�.@P����Z�e!w��#x��7�T�ݷ�CR#J��+��zFD�Y������3�fN�(� ��qÜ�-/�;~�[T֧/�?s�{�6�Y�|��o���9w��p�,q�%�F��
�m���ω<e����V�56��|�3 H�����������bU��t%�T��Z�h�R�tf�N�][�a7z���`���ry�/�T�D �p���i�؁e��;et8��So�Q�5��B=W*��*O�U<���w�}�M���̈́L٤��2�z��N0rZ`ET��A�-� R}��VُH(��Ϛ�C��ŵ���Z蝎8���+�O����;��~��D7JK(���o�ao�s5Y$nK0m<�$�X���[�kܐr��d)�^�0�k���{aQ�0�Բ����i n#��yW�.T�E�5[�Fǜ\':.hhe\�-��L?+U��"K�������d�b�8� 5^�����

`F-����m�����+J�z��m�3ŊC2�xw$>�Gڅ�ޱ��ɏ�Q�����;��c ? m_�f���B�ߋU�%�Z�y	f��Vo ĭ�	�E?���]�=��q��?�Ļ������
�֛�!����;���$���mf�)!��%e��H:"���!qE:��CU
[s藫b5ʁg�e�[6	6K������� ��@w��F���b~�o	Z��@�.�<Ґ`�Z�*��Z;�;��ت�8��9m����C)i�5�'E�*D����/�O-.�'uc��gxt}_��A��YY�I��t��;2����������у��..�7���Gˀ9�L��={�2��LTΔG�J6.�:O�X��Q�lEu6g�V�r% ����*��>X+��5n̏K����U3�P�9c�n'�X:�ι#��V���'���J?���YqO*�z+��hK��fL��@�l}�u����/�g�BK��=:����0E�� M�ꘑ��D;�s�ak%;1�kZ��RNK��pc����3AaөZ5ۊ@��gl��E�`�v���,�j��0*]f��؅0ੑMF
b����̼��e��x5���e�a�K-�5���)Ӹ�X�c��tL2&��l��2�q�x"T��>�X� �H9�������ƨ2�<[�:������	]h�'w>q���^/C�o���,��	5�hkN���
�/3K���\�5Ϸ�>�����O��������/Ð�q��3��Z�4�Z���0,��՛j��� �2F��.Gz�+��@�:�?��F�_��Y�3��P����Z$1a���k��@j�n4�l ��Xp�LO�-^j��K���7��|/m_/��;B)<G�� ��I�ݰ/��}^�F��%�����]%�����{�0�o2�=n,U"Ń���f�z�t'��XP�z�
�$ ����P�}�])�P�<�$(C1��l���;�lD~l�����Se,�-x�.R�q��h�5{vB�?��tJ�w�[�zm�P�M�J�WB1���2Z��TNɱb��@]m
X��i���ڨ���� �n��!(��q���Zr���k����V6��+A���	\��B�4
��x+e_"�'X|{�	�Tv�eS>�~�0Ӿ���
�S�GS�o���4q��Xmd��tu�-��BG��O6���A�mT�{+�?Μ�`<�krl��l'Ȁ�5�'��y�6���W3�C�8�z�@���'�1ׁl���Z��O������oKH�t�ŷZ��o�s\� ����h\_��/ ���	֥��}[���E����T,/M�oL��i<��z-�n�����%��D�b�Ys��˸h��=�B;f�%l�7�w�}��U�7 u��T�`f$�#�)R���B�<��>]Җ�wsaR����B�@�B�	���,Q�(��/�$k�O�¥3��Ɨ�3cWR�i��&�́\��;��Α���U��J��KK�fUBe�hN,$�`#�~] SPF-�|>�/���ܝ���w��;�G��i��K���#���֥VൌT	?�As��5:��a}���<����#ZnP��Ev,�H/�F�x�M�ׯc�M�?������~xae�!�۪��N�&�x�����7� V���m�Q���B��kf�=��K�l�dSO&���^�u%��@�n�z��,��AC5�K�.P�#+^�5{�W��%�^��N���_U&��~�&N�Ǫ��yi�d�FT)
T�zgw�� �I��C�&H���@��t�Er�z�8~�R�f�1����ԙ:XϺ0�6K�I�K�N�2���8��H\�Tdkw[L3�h����/�	+�k����=;�����M��A>�
�'f��?�
��L�h2l�nN�a|yVH=x�5���_vZC��ɰ��)Ȝ��u���	.Suޤb�#ƒ����r����9���w�˜V�����7�ڑ5�&�G��9oA�Y�1�g��A�o��MR��!���\�k�����K��?�ƞ�.�J�@��A�M/N`fb_1�Zh�A�ȩdo�Ŝ(�b��r���hdv
Nz�}o2;�e�N��V#Y�N��j
���N- d}��%�OQ;E"I���E��V�\&�N^�^�����$��+�zG	�����:ۮ�bA���G�T��~��L��{M|�m�ץP	m��n����}#xYk|p����w_7_�#�������Y::������5[4BE�q�c�;�i��%
��A�A��/~��Fl-���PܿN��6sw�ղ(*l�'c
�̖0���-�kT�V�:��n�d���=;�JYP=b�h��b$u鱵�Գ:�(x[鿙�\�GbK����[�[�4�vg)�g���W�Y��NT�K�f2�����$�DM�zZ�D�{�!n��~�]�>~q��,I�ۮ��yh8����Qc+�j�훅~x�DRg�q*T$�v`�i��f�i�o�8)��` ���+�:���]-�Ԉ�ؽ:���ZT��1h�Q���E4��!��\��d�y�����{|������-	���+pv�3c`LۓH|�qf*/�o�~�����B.\P!Yv���:_�1"��a٦F�5�&'�K�^�+�\4၄�����i��i�x���x���-@: �v3�*`jd��<�өz�3���٬%y����L�GO�6�0�2��kG���ȃ�m��%��m�M\���T���b��I%4$A�K���2�ʀx:<c�Rd���$�*�z\�D�6��b���\���������ӄFA�(:A�a����v���8:�{d/W���@%�:yq��j�.w�Kfic�<��my8�v>6}ÞQ�ѐM��]{�c���If�Ί�����4�����?"L\t�[��)H/j����F�� 2�-�Eư�-�����Q�C.6Zc��WSh���d`P��OVK����(�?���>���w
}OMc���A5����s��8�`}�2�'�P��5����e�(~���{fH$iKS�����	"wE�ɖ#���
kb$���=Lc��~p1J�
�
�6�+�mh��L�p�M�ǂ�&�����n�����s����n�Yd���L]�.c�B�aw=�YR�v�M������GK�mbr/ ����8^V8I��*�)�h���luٴ�U>��d!@Q��U��0	�4��.��p$gvn�+-��8d]�ec<��2�l;�#ģ)4�Ͱy�D#����hU����IG��8	e���DS����M�I��nA�W�}��@��P�������]4h�c��s�I��8��������CW�n5���x}�n��YϷ}ț� lT�}��p�aܦG�
44+(�0�����l^0�=[Qc�u^��^�;�T���7_*�3�� ��	L�U�2u@E���D�م kz�K��KL�.}�ψ�uSD���/Gat�
���!2o���������"o���yNv��t��ZP�9A�5񤐛r�Pe��h�z,.{����݂q��s-�B��h����Ą���a8.4$�eJ�^G�ӚN|�q"��(�F�B���J�H�v��݌ W�'�Wz#V ��
���
��f+2�?�zXQ��H�����(\�C��6XިkO�n��X4h��'����Id�@&��`�����#�bW�y%l���/-�n$����S�Em�ʲ������1<���MY�	�,�o�� Ԏ����[,��ƀ���i�v~���
rl�K3�%�hL[O�5����,��RM,�3L�*_�nQ�	'��L�n$w�u�,w�3�c5��4!�)����JA�t�ek���S1��+ԋ��u:�%n�d<��R�V�U�]�<.������"^&���Z{=��ςKv���P�L�k+ש8&#q�Xg��h!��l;x3�d����d�"��W>~)7~U8�Yy����IU̇�Y�����^o�d9�j���,[��T)��*Bdf�g.�)�|�bLW�kʶn�m_q���|��U��zeN7^��_��JҠ��I�s���Xy]I@9��:X*��bo�c�H�3��ɾߑ�;��8�s#�-�}�|�b-�D1��9��j�7oƚ�Q��Ő,���hO����:�P֯a�����U��7'�ԍw���H�C������x�f�ւ���J���B�����������8 "�x8�c�>A0~����)�x�鿉ޥL&�D��%��&�j&^t�~�=(��l3���������y(Y�N��!���F���vХ����%��B��&�J6�fd���.�a�T��i~/%K��g'�;B�=k��q����lI�Gt6�Νε6H��F�)/:LE��s��k��~��d��;����!nΣ�N����z����a)��x#��]�I�.�"02-T$�WH�q)�?��=(EP_��EX����G)`�^�W�#��I�8�%"���<>0��<+4~�������&�e_I9��2��]k7�:�}Zi�&�Ĺ�����d R�\�0�P2����aa�ң�H,��A5��Q�Lx`׊Sgo�h�8o«;�!����.�p�`�Q���	,s�s)�uR߻���}5��K�ą&O'�dg�~�kLn��8��o��RQ'��0�1ޡ�Y�b��ng]/��}kZ]��=�d/�dfQp1��(\�.��L����$|���	&+����b��I @�����	m�r�o1�kO��o4�Ї�L��m������\�	W�7B���j W�"��s%���r}%�a9,T�T��ڵ�u'I�������&��t��ύ	�Ej���d��O�ķ��h���Nk61J�l8y��@X���b͎#1$��W�TY�v�"���K_��K�u&�T���	>���9h.���QY'b�'.�*��*��G�ǈio������f����_�i.�:�T��uE�%z�^�#�3��.zj(�a,��	�RNS?��$�X��n=���U�
	~��$t'�c�K�P�?�^�N�?��y<�bӊ(�Z�&�e{ۤ6c�쬕�\��Z`k��>[IxX��H���&gt'-���DY�9p�.G�:��u�C'���H	��z85X��T利{�p��eX
��]ntve#/�	|����gJDL�L���4㒝Ty�X������)����q�����vy�$�=�*7%s2{�����8ǗA'��.�6�%�H�0(�o�.� �+���;jb�a��!B�*}��E�W�ez�I�i���4�?n�|��׌\��=	ֵ3:փ#L��O0�+��g�2�嚞7ds����w�)�����$�ӫj��(�P&\��`h��23�:�G0�qE���}�_A鼍.5�+U��椶�j�DyQ�¦{S�f���snF��q`oz�t��C|�!�<��[NAv�!Bm�C��y�<�'���ƊF�k�Q���W�sׄa���)"���+x��ʚ�Y�y�=�b�S�(A�"Ckg[v2T��X�Y�u��2��T�� �:�x]����o��`��<P0B��EIp1�BS6ʼ��Dە�������T\Ï���M_�=�ax�1�wD����ydT�w�-T8�طkzj�-�Qi���@�y��<�SS�_�� f��ϣ5�?`q��:�L�����F���ߢnF(0ܦD:O빗#7f���r){qh8M�7W~w�n=�]�����7i�r!�Ѯ�	^;t�j×�����u���$v�*�*PK^�0Y40�����'�$n�d[[�K���o A��?%�d٩��8�l\�(���hu���A̒0�F��s�h+TZ(�g�餱��K�� �-���F|����ˮ\[�c��?��t��E�z:|��EP�x&��_M;	�!G����nl���ج͟M��Qj(h�l�M� �֚!�x�;7�[��/�!�� �Ju4n��
���6�2� x{��*|u��0g�Am����* �m� ^�b4���nm�1��{�@ Ó�!������.KV��<,oQ,��$6�Dm6*A;_�"B��C���C䠸�����V���#E�iz7VY��]�ь%%Yi+^��ʔ��cXOk�B�7���X�9Ge�c�)e p0=��$�$����e�c(�T=e;t��*7�����RQKK���)�O|Fkȸ��I90:ٔ�%F�=���y��(ϣ�׺�ȌBfO�h[���ޣ�������LH(�!�*��8շ���8��Jg{�!��4������O�W}::�;�BR\�6UO���1�{�

M�U�ԨS=�E1l˼���7-�_��y�_(��d��"�0�a��
�V]{�)P���>ő[����{�B�zY:���h�8�S�F-cA=p`=m<p�Z����_(p�UK9���dȺ��qmY��M6P&�Q3Z�ɚ��!����V�A�b���חkw�|oj�̡H���"4,R���x:�&R��������ֆ�8Z�e����4�X}�O����q��(r�c3�rƍ�\NŶHK}�U��_���,V�?�/ެ��*ē��1*�2���A�4r�����_��\����t�dl�P��J���v]`P�J�����x�3�d�b`�)i��r������Y#�7Q��9O�Y���J�Iv'qW+C8;�;i�T?iɶ$UF��g�ʮA5��Q��j�"p���gS�~��ɕ�[0v O;��:�G�/��nZ� ���� a��h��\l�6'�/��+P]嗀9:2��� h�b���������m]
�y��U�k���c�by���3��Ȏ�\<ܔ��k5���!s�3�rx|'�R9�=
��y�0M,�<E&#N��+k���炛�WH����cEQ�$�t��?t�:��i!��pz�&��G��O�MqT=Np,󨷒�9��A3�D���@i�c$���������@��EWU��VH�Q�@�^/k����u8�Li��0D&����u>�2]�·�<�6n:7�\�N^���2L�+f���?�Zg��|�����:�܂��G�t�Y�<���DD������o�r�4˘$�u����Cp���̄ ��I�K�l׃5��m'TqF+�Sj
ӕ�2[d�9��~�_��^,��3��r�v�Eic���}�
E*3�<P\]������נ�.n�������P�ע�u�}e�[9H˲���ߌa脝pTguL���UX=�;�Gn��ub�_Cx��8�OmΜl����d3�N$�d�.�AlnOr�d>}��:�x��R���0��:����y���O�V+�;��UTL�c@��:V��1#���,�����[	B#,1����0APP��/PG����qB������̐ԗU8hc��f�G��\��B�����,"������S��\��y;��|K�D�V/m'� &5�?���R��%�n�4MYCS�����a��Cڑ�� I�
�0H���2v�#iX�,%��4�|�aG
?���FΐL.@^��fY��%~���D����;��8��=��g/��gI��Q��:c�䥽���Dp:G8dݜtHG���`q�ʒ��g�k�:k(�B��1�?ar��R)�<Z�ɷ��9��`�Zc�*�:=���؍+l>M��7���3 ��_�s��5s��P<?�w-�~/�;"C˖�Z��6XC��e�T1��
A���9ʐ��A��肿9���*������> �	֪m�0����,����s���9��7 ���pNY����?��-��`���'!m�����Q'�ɪ�"W2��9�x�ʌT�~Ui�S.�С��#��TM��	z�Fb* "��{ǲ�y�>���2��[e�7,�W�&�4qdZ�g�}��(�&���oo�fn3��l��ZT"��ۃt�I٬�����J�ШyE��R��EW3ݏ´8'@I1��W{�}��<j]��U��1sZ�2�NX�Bl:�Z�.&���4���o���{�iK�J^��de���w��̱�[��Ax�tdD��ӐR��U=:8wV�ٓp�A�и�u1�v{X[Wf�@Z���1񁪝������G�8���ê�v�?�m���:݈����-��w����Ґ���5HB1دF�-�z�UY'IM����7r�)�I�	S�<c��n�)ĭ��9B�68��	n/1������Y W�Q3\'��M����������8�(ġ� �yc��ML)�!ny��}0���!�?bp6ID|',�`�b1�
��!�����=HW��E�<�J�
�����ϳ.�P'�f�B�J\�F~�(��iӫ<L�W�+�ܴ��#��+��}��L�l�p�+"��✜���'�R�L�����+���c~��0ӦѺ�E�3�uG��ggn�R�V.���mK�B�)1��r�z��@R�g��@��+����@�_���go����u��h1�(�O���EB��$��22�G4��#-1*����$w>�0	��qF禕-��`���ܾ�W+N`���|�Mjg�7S�@��?
�(!0����I��"s�Y�'���x�]��O�"��H�_Y����9�I�֟|l�:��E�"�Q�p�^�y'[�M�Kې�se��~ {�=���62��p�+������٠��隱&�2z���A�v�>	hB�3�����O�/��)�3\��UXM����Bb-b���uB+�K�"cI���pc{�7�XI�h��
��2E��f���B�I0"	&�*jn_����*�шA�����+���JL�G\��w�5v���������v� 3�M�� �D	>��+�~	x�y���%�(��T��N9�J�p�@���`� ��P���8���B��.��m��4������<'��Y_�ȥ�B6�.%�)Mi��^L�_J��&9'S���jjX]������(�"-�N@���v����wmS�cp��B��G�A��P0��oA�QѾv�w�5�2��&������2{7=f���z_�49���o`��s��3���eV�|��d�6��z������-��vW�Z�V�c�@� �97�쯝$-�5�캌n�qPQ���|�Q�E���/��~k��I��78�mE�� ��S��=��duB���P�ͿbN�N<7�w��/�n��({c�K|��S�E��.�@���JF�U�ۦ�y���-3�r`7	���>���E��An6c�o�Ϲ��u~����&��C��/���uٿ6��f���KX��^A�|w5��v�e&9X
Z!���x�������]r���5,�[�H��!��8�TB�a���"�p��.�W�)���O�;�e3��-Z�G3�����Y�^Lm�����S����1�z��=�
u�l	�D���F���"�W�zхRL��(���GsG�l<�dz�@)��{�F��$��ux�r��Xd�����jٻ#�t@	2���{R��R�PR
����x�ic��Ո���@9>��N��R�[@��:�<w�kc u���B�3�PyK�yW6��b�	e7�_�X��㶁�Yl���J��l?��dL5���1�߅�T㦠�"�D�k)6������\��]�����b�7�����ך8\1��![�L�e^(�n�r��ǉD/7��(�m�/��2T����}t�)�}�0�Sv��Ҭ�k�m�K��SsWl^�W��~����-�C�VB�7�8a@����RN�{��9x 5q:���I��,���.�X;�>�i�`���}��X6�A"q�{�U�(/���*Y��̤��̴V�r�|��^x�I���u����:D��bוR��Z�������!0Ɏ�5nX���&�_l%�� !f���\�Ï8<0Ά0P�8;�a�U>���4�,�L��mΩj�^�L= |ES+�x"�z%�C�8L�Qޛ�����Z�U:�W�tSR�;�}\�C����q�Q9�@�B���u�|L��?ߨ~ay5��3������l
׌
�^(��Y���L�ʵ����k!�N+l�a�jV�� �O)k��`��@�4�I�<�������c��v(�uO���#Seȅ���Oԥ�L7���٤�Q,���V��i��Y�L#zRR)�x�ϋ�M����F��~`�5pb���ҫGL~��S[%����	(?銅�^���%���wm�1��To�$N�y�Ve����={�ݿ�'Y���,��Y�F�ˀ[_��q����?/d��ZؑÆ�����ouBN��ߓ_ˮ��TS�j���(&r�0z��֠�0c��|SGI��p��I�������]"GF��b��A-��'òE٦g�U{-�/���H��ls�n���o�M���A��2Ft�
�@ �<� ��
��ՙB�����u|ȈƩ@���pI��y��X<.>8�ҞL������2���<-u������X?QI�t��~g\d�j:�X�G*)p��Qe݇a�/Fi�z��-�L/��;:�X��k�H�s�FH�c��i��ݕ�*�;l1�9�}{���9-{���}�q��f��!Ye�1J!�U���J���Tr��罜Ƨe�ʊ�ZŌ꒰�}�*��l5�i��^t]]�Lv��ªDI�ln��j����}=�&�N"ᓑ[-��;���������<�x�&�|��#o�R�ע-�]5`���~��HWE���_�^͘c!@J��zi��� R�}�o7/�/������oKk�1-�Y�>�2���D���H��{��q3���Q�HzY����ٍD�� �����+��;v�=�X�x�A"i#��14иt�t�Q��oP�!��(�y���W�Q��Wt/VXw�rA�K��#��o���y6�=Q6/��I�\&�1�f�;�vv�eí�j
Q�Jn*�%>�@����V��l(�3�C������Dγ����]�h��}�,��+ë�.��Tv�㟚eM&_�6"���5}6 �	�A�E�Id�<� ��k*#�u8��B3�SN���tE|�@iJ��0u�m���0�"�k�#��x�n�=�;(؄�0��h�k�V�ޭ���~�^�;H91���&�]�H�u�A����L�w;+�}l;;�LyBWNC�DP.~,�Rϩ�G-5�q(�T�c��>�=��I�i�{G2z-1��kWݖq��ͳ &\}��8��Xd'��ҥ�Q�g�'�$D`��JdH��>=�s��2�b��dߊ���2©����U>�nN�qyx2����,D��7�-��]^�%D/�j�� �ɽ��-Uȣ,y{߱\��@��n�/�����k��@��Z14��^���hk�d$W�3����|V��١�̧���G��o�l���9�����f.�KS��|gO���A����:-�J���.?�6�՞k�I��SS���ǋ}M���!�IG]8���TC;�A>� 	����'���Xï7Ika���������4��4'�� ��t�l�b)���>�ܼM�ׄ�|�4�]5�hc�"s쨶�{1����D�\%f�mr���I��NZ>�K���>j��Y��{�Zm~��g8����/_*Ʀ�EJJ���A�_���?=O���v�2

��d��CNlܼ�B9JU�2o|�H�e9�U��A�:(L�C��&���y�!0����F����r�מW�s��F��u���4�׊���[�l�?����1۝R���g�9p���pd_�xl\�V��h1� sx"wt'~
&�������H�(�O����+˜� ?�r�;Ɉ����*l�gm��#�B��q����� �P��u���V_#����9�v���霯��s��堄��rbZ,�=!vo��lQ��(���J1R�m���m�����q��o8���,� �P@��w)�9}i�C�����W�T�ΐ���Bf�������KЖ_^{vrvH�Q�8껓��4�u�?k��lb��(� 
���YI���s�$1�q�÷�L��cϗqk��9�OX�TA��S'W"ðYJFN�T)5�Qf7q�_��柤�	d�)G����J!f��G�%�u����E�!���Ǘ�CB�C�����v��}�X�s��ԌS-<�9���X�2����g{?r���V5}^1E*�����.��K&O�7�{��Z��N F�±v�$��������Ҿ��',8�d���Ѥ�x#�|؎�7�i��N����qb�^���6�ɸ*9�hH3՘*Xo��O���Y&�Id1�ֵ�yj��e������O>ڌ<�W夿�dF�&)��	�G4�?-�s�Nr/�l���k_������yzut�cF,�]�&u��Z�g�/>>�3��VJ��8�q���;a��A��~Bc���
�mfn�)H�K���M�~#�CC���x��]m;�#_;����YE_���Ii��e�6@���z2����fY���;p�b����YOs&�A^%'� �Buર��śxRƢMin&sG����^�r�z���v���2���<�}�1I&�	��0'iB�Ğ���j߃'�s����[�o��� T�:�a]���_S���>�l���A�E[��r�c�(qXSt ,�聴1�p�q�T��)�M�n�;���{x���!;;U%F>��CDe2?�0Y�]�z�퀈�y3�̙�|��):a��!<%�M���z��\9�oF��M�Y�K()(�%�E��������FC��J �b]��Xk��_����u�|5I��#�~Un�=F���� ���W���_D��ڃ����=ԅ6��ꝏ������m-��񗵨�
�,���f����¸{�A�K������f>���H�Qf�a+M�9ݗ4β�M��)�̌ 8d.R�7�o��~r�˞�;C��r������3�_b[DNv�W���y/C�xT
�X��$Zk�۟!`��I�a�]�c���r+	��($͍�āW���U���,ًs�A.ߩQ+��JD�gk��&�U�UL!��LT�	6�UT ��/fsyN�(�+3�dd{'��� �[�����W)+��~��!��L�SM��A����
��ݰK;��F0t�0m ��%��	�������A.:W�-]
��He}FRG�?�qX���!��jPyUP��z�7�Nh��O���{GnJܕn��[ʱA�]ͺ/j,�no�ə_(�4��[���P��e[k�0�Q��h��c��录�j�d�GR�Ӟ�q�{�S0�8X:�fnmi�溧DxA>dY2��A���cJ���EQ��B[���q��a��c��]]@&}��l�\�f�Gn���ʦ��@��(�u�|�T�,ُR�XҰ�P�!%��B���+��[�oY�eX�pr����b\���w�}|gQ�Č���/��3�����{c5ʾ��D�a�`iЗv⟁6x�x3�1qS��Cf����CۧN������F�J�0u��l��0AmAC�Q��xm]�q���#����GI nRU?Jn�T����\�2�9��@�"He�hg���RA�
/���r��� )�>���P8e1�q��k`N�Գ�����0k�OV�a۝���D��'�J���6'��E�I����x=�k�ԝ@�j��Ć?�_}gj�ɐ�Oaw�kTg��*	�����h��R��|�<:s��г�h��V�r�_g8Aau��Ku�[dMSCn�u2�S#P�J������ӡ=i�\g+S�W��GN;�.�L��9�44�@��7˙ȥ:ͦح4�3\M�R��NM,%����9�>�Շ:X|�����ö��Rf�m��$�.��x�(Y�r ��p>�S��eJ?n�cS7R��&�/_gi
t�J�~&,�'aX�A�*I?���/�=;�z }�$��F�dG'���<������e�b��Q�;J����i������jm������$��Y�䯛�cdY�?�j���r�g�����\�P�ܧD�z�;dqt|������E��	?k�Vl"�Ă���FH�����I��$%g� ���o����T]��4���`��A&?k�
Kۡ�|�CR�d�կ�!j]��Y
�B��;�@�&�W��Q�Ώ��e�\��]���%�<��xG�LG��� a�d�;�SK@c#�g�vP�c���%�Uufw>\��>���%�&7h�|T���R3��R�� ���ͨ�U��U�r��
;��G�a|��9tb�4�#t�gg�v��w�Od_�9X=o�qڦ�I52x�	1�-�l�Z��3��KM.�s�}Cb):�eu�`c�]���В"�e9(l�"R�l��DvF�+�2[Z��ݲ }��������P�\����1pm���:�|.z��U��į$����lZ1:R������.3xu�,7��8�t<vzԈ/t�\I���7�I}�)?�S���9�R�c��`��#������`��'h
B�M���S�g��]�c��Mi��`Z�!�bR� E�k�Z�+O��cW�$%T~��l��>j�ءND7��=^X�/]�Uʧ����tX���v���ޕ�*�?�#1������o+��O E��5\�bε���a��z��6��qk��ETF�d,�LCZ���
kֹ�E8�n���A�������ł��d��D㢗r��{d�D+M���f��>{�:�L��"�s���A�J����6B�J�/�Ӿ���\���(�+��u����=���o��3Rb�&�Z�=+sݦ��χ�Ko��`�z;��,/GQ�^���W$ހ�ϱu�;*ucM�K���q�c�4�c��}.|u`my��CU��5�Ȗ1����/�d��\Í�.[��Y=�;[x�)�v!�q��׽� ��ן�% �E���gƇ5x^u�y(�6�J`'P�q����גEB�K�ٓ�s�l*E��'����+"3>ƀA�e�A�Zͯ�m-�yZ�-�╞�
�
-�ҁ+�I���8���6z��A��c�������?|^�)�h1��g'�B��I��y{l�Uܔ�<@l�7�G�9����f���4S��ϫ�w(cXؼ�f�FQ��g�ڙ��6"Ѓ8e.ZR崴P���.����Pi�{X��$�W#
߿�����C�,����W54���s%��m)9?�S�-)�7/�_6ZN��%�ј&E�T4�y[�DbW��7O�z�dH�B\�R
�ƣ��B�[�6����%��B��E��F�B��d���wt�Ѐ�NKQ��e��D�3,�w�L�mp|�g>-��}�'��A����g�x���8QO�O�slVU`"^cӒ�z�����R
-�
}������v��]�[a��m?����[�!��,/@o�8�|o#�H��,�tt���r�T����u���)�+��FG9@�9��)����ʬ��c�P	J����S�A̳�l����|��%Z�P�ɳ�k�[�md�A�F�s^����2���<�w�\2��z��8��[��=�:���[�&��;ݣ�ob����G!� K�
� ̃�s�cL��,v��J}�m�ې�4UU��%U`��/����=-��f͍�v���߱�\X���^�i���d��_V"�I55(�WT��3_���m�dh
�v��u�9�@��i�@̗�g����6C�-^T���x�D �p�N�8Vw�ډ<�|�({�2�]�X��df�=ȣ:�;_�4��u�=�5 "7�������It�u'##�̜}�P�Y����@[�Ю�����Go���W���p��qnï�b8Ѓ���A{_�Q�H�9J�"���FHN=x~0̈�?a&�j	��r�\�b���`�񣰼�����Q	���Y3[����r�3�	K�rZ��m�E��2�x�zGmOU���I\6����J�(���?�:�	���vk�Nr�`�����Dh��m*��?�w�V{�S(�SG�^�H&`�������و0#녅ōӀG˨i���OD�!D�y?}2��y��V
�(X�[�f����:��K4������o���(]��Ƣ#�l9����6~B�T�=�q�̈- �i�A�:�=���ݖP���_��w���)9���s�}��<�M�g�6&�Dc��Ho���c����kĝy��(��>����}Y*��Д���;v���o�a2�N�U�٫]�d�y��b��	�������^�{0���?u[�@�/���y.<���6�'N`���Ka�@����Z�)�d+����Q?�?��DB �gvÏw������	 <�0�Ŗ�H�zɓӱ}�6#�o��5�d�M���R`���֞��✖����ޑ9��� �ų�"8?c���?�ˏ���FLc<��GE��[�� ��&H2��������}D@��cG����Pi�#���� CN�-�R�b���E@���!�J-L�E��4�[��p���a��W�g��H���}�wʙ���nMr!���%�G�U�k�%< �h=}�fA�a�I���`	�g��WWq����x��%�Jx�#r�ˌ�R���O��!�^ ����#����='[Ȓ�>��	cP������o�}=o������ܮ��_��`�,	���D*�
 ���{��g��-��Bd�v���;�PAh�u�!ol$G(�����2p��$��������ۓy��+Z�xrbPN~aW�qey�t�顛�TA.��f ȩ8��&���Ș�6�J�u�U	�/�M;C���H�t�[��2��D?{�q���G�G��y�?�����'����x���)�*����m���~����s."|;Ӭ�,��3˨[��Ұ�n��Q�zc=��!s:�KfŇ��2�"3�m�4[���i���w�ic�<Aߛ�2<���fB�
M�=M�͒7H?0 ��}�֭��R�b�N�M���#t�R��QC�	;�����Ե�*:P���\#}�Z,�/�BaƿT��:�3�|ȡq���AO�F�r��g�dޕK����[�~u��N����y��l��o����W�� H�+�,����X*ω�q�u���O�]�u�nJ-:53!�(�5�I��V�Q"������ف�װr\�B?��U*i}k��)���#!��ly�h������R��P����	�����VTN���<b+��\�LP���r��K��p�Vj3�[%��X�2�m��A�{���(m�C�w������r�	ݗ����$w�u��#�
�튃�8�<�D!���%g`wD0XT�]�WȤ�_#�6 ��|M��sD�nD�P��r��#�Ox'���g�0#4g������	q~TWg���$��3�պ�ۤH�bXN�x+��oM��2���5�-��b�Ry���Alf������`俏�i�2�0 +c���X���Wr\<ks�G?���{eҎ�|.����F�w+72���t�9}�t���?/̷��7���;�Ԏ7��x���|P�ʸtć-���������<�U0nɥ�A{��Bt^zA�^��w{:@��u�v1N�4����[/�Թ9����*�f#-�W��c�!Ⱥ��w��4�<�96��<�@�VJ�_���x�U-a0'��5�HoxM�/9S�!�z�P��n1��t�i�������	}�y)�J��mW���EI��-�6��\^8w�(G�_���<:1�O�G,cW�I�M�K�Mj��C���g{�pi8g-���F�*�=:�m����\���H�a&,�~�٨P����E��0ޫ$ ��E���;���{ @}a�`&����ve"�K�!f��2�aTɕ��6�8�e,;����TN
��z1��ġk}3�0rk�wR��1�A�vE%�"�LHO ��~�J� ��'{�\y�m��I�����]G�C:|�?Vn�K�WZҦ���3�\�f�]@��s��<�.h�������!��?�q�M�����&�!���s�#;2��n}=���=(�5>`1���r{�B�l���=4�JK��6�*�-�'�6NS��Dhk���$k��xH��)A.�*�uu����z?�$Y�;��j�������8EG��M��{��ƀZ��I��9���R��nO"@�S�H�[�� �]��L��yvgz�&n��$���D��'e�L�b{)� ������עJ�i �Hi,K: �^�q����yܣ|�$��۟�0/�u�T-U\Nqvo�tH�fb�t���{�x�[W憓�3����.ť��]@�z�����Kr���B!n�,��(R4A�}��!��M����f�!wf-�d$�-ܼLD�xtf0ޜ��W����H~LoJ�x�e��8�[ݧ�b�#y��d��r�Sq��u�vG'G��_W#S[�Z�?ۏ�/�x�@���I���\x�	qMj�x��%44��&u-o��f�:�.y"xE�	��-e�������^ �����B1��ɛۙA"*�;Nh�eV��@U�\s���a��k#R`(A��L˚������-gb��A���������Ɂks����U׫J�^��Ax�hs��m�A���ʄ���X���w��)W�
J�?]�*�d��LW	J��x֣����bc� uk'k�կ&2��9�Ir�GM�wt"Un!�!����Z�mԍt�Pۗ�X��Q��?GH);�o������HՈ�n#�����_��3��i�L���.}�c7��ˈ؝X�� 3�فmػ��UE��.�-�=T�q��TkiZs�j��r�_���:@P2�.X��0z /�^;R,��%.�>�,�魢h7�f��1�, t��YP�S��Z[�E��=���W��:uM�X�����X�:l�(�"d�X.8��5��&Lj����oAHux�2CS��~.L���ZE�~��݂)r�o��~���d*d���L�sh+.d��M�1�j/"*�Z�CM=>``m��\U<�G��Q���96���8_w��y��M��T���%v�������������)�#�c��=y��h�����U�����,8/��RW�d̩�Q9|��g@�G.����6��]��0�B��]d7�e\�Qg�9zc�$-���H��+�};X��O��񲤢jK>�J�䚱�Ю�����j�����w5��Z�H�9PGy�U�k�K�Z��T1���)��k��t3��i�gQ8u�۷"x"JE�5f�����ą�.�J�h{�*��a4��э
s��m\u��J�Th�9��r|$e�w�D��b��T������&�Us���_ad�DR5_� �e������5�¤^��Uq��'�,��"V\l�KȊ�*τA��s�,�p��~���|���2f��c���Dz�Z��*p�v-���-HE�A������XY0�~r���7��NAy�����tk�^��ϮG��)��'1��`��
�ę����L�5�^�Mp(���6�C3#;	���ᑝJ/�sv�H2@v��|����du#�2��^�@!X����߻9<�)tZLW��B��C*5�+�Sc"M|�� �IOJ%��%�t�2��q0V�������$���j{spИ�~F_y�i:��U޲��!%��j;A��F1K�}TdD.�6�7�s�}�ܸc����2x����C��TZ�*�Er/����l���N�v�=����^ _��"��z��Kp�ǯ��5�q���`���&��h6�Ƽ�0�r.P",tUfD/e ���=��<7��1����S[����rst(c���з,�4I��i���a����q˥�ѝ8�ZsH9�|��d�OXQ��	�j����aȐ���:��*N�
J�"FHtQ#
��_�IU��Q��(��ڻ{����tă�~�,�ד�.4QM�z���"�i#�O��e�[��Ԡ�˚B�t[�''����7������E���=��O�#H�ڗ~M��+d�t��d#�'��g7�5�I	7�}8s{��T���D>������.�0m���|�E7M� Pr�G�:Ƞ��8� X�C�͢���L���7�������:����ڀ�M%����6(b��Gv�R�Kf�����[ī�hp�ͼ��D'2�����7�d���)�ʏ�W'L���9����O"�F��6�3��N~��>��G�\��,���9_7��tVh�D�ݒ�&S�;9�L��8�U��3�_���캤�`��G'��7~{m��?X=u�\�x����ě-捨�7\�i�/�$�Jc�G_��ɇ����w.N�^ &�&;��lO�Zq���� �tD~nW�b��,w1T��+��\k�8�Q@i*�/���L�\.ݿ]^њ�:�6� -�	�{����/����|��sO�/�a����7���w�uM�QT���Ŀ��d�Y���,5��}����o%ΒZ,�!�9��(מ���$���N�}��@p���dP�_iɶ�%���h��bGU���NR�(�l�X���h�f9Z�F`��S}/ƙ-)�[�)h<�6���X������N�v�|5����dTO2�o@P��V��<V@�p4.���m�>A�F����65�>�Q~�ȡ��n�kgIЍ�(-�����