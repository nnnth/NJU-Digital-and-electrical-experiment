��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��2��i�;�3�������:����Gx:�	A!Վ��O�:�''>Ji�u���7���K��Z������G�

H�H}I�H��_YD�@�19d�%h�B@���q ��	�eQ�1;�ޒ�9F�>е�ax��Ȟw}z�4.gGت���� $y�;Y���[�[�a��A@��1Fk}�j��3U�B����U1�����pq]&�ȼ��+��ap~#���@c�,�2VU��k=p�Zz�8��#.�ͳB��̦�I�o��u�p _�U�M}T����o�ur#�����g?��V��r�zNJC6��\ ��vo�C�Cj'�e5���Db�Ϊ2z}r�ҧN"QNjR�s�g�����~�9O�[��K@�g�_g���5j��!'�9�)	` ^�P��3�g@Ujcg�m�#�΁�ӎ�|�%�1Y[��c��jEw��F�8>i\��t1.��� ]hӒ�B���X�'��@�mc���H�(wm�u6ݼ@i�
pJ�ӄ�����o�l��B[��K[����W����������¨9f�#L���Ƒ�&���<����!���9���6΍�`IAT��JEGU)Q4�u)��X�F�ڦΓJ��;���QOIN�m.xt���^Q�6sU�����%���(�}�a tp��,�Ն	8��a3�*���|��ۉ�<��?��S$���������ɝ-���"��7(ʥwAZ7���$8��M��`�U�Q�'D(�����O���ՠ?Jn���,��[ȷ�
�T�E��m��t_T�T�..t�ϩ`y;gL���4����Z��;!XU�~_�3��LJ�v�F#k��GCNګY�H�Į|���O�a`)�#w�9�����n�)x�
��*���懬�>�
o�ȼ�Z�fA�HR���b/�	��]%	�P�PY��Zc	��%�l|��y�e���!F$��!KV�O�e�}�4W�~�V��G[]\��n| ����v�D?�D�Ň"�}�/��_�b���׏(f��tP^���P� ͂��/��\��i���@'aS_}b���>+�.Q�Ѣ�KO�g�HY�T��KRZ((�`���a_�y���Ю��q{���E[5��R�y�B�˺�@�+���)/	��z�|R~��>���(c`Ϭ"�gX���������Ey�ܺ����H�߁��=���d�����_��b�@^a� �E�}�Cr�$�2������2��כWy�J@�:@7�z?���H,=� F��^�[h�Q �N?���C������?f˰����
Q%���aQv�__F���dV�j��x�M��u6@�R�mڸy&�i��r�J���~��fM,@j�����|h�\�Ǧ���_I���QI��$�&�����;5���2�k覐�w&
��d����f��p�6���f�����9X���yuӕ�x1�\�M��o�o\�9�DKh�(���fXM�����T`�ȷ-��l��!uwEvP�`���y9sx�oX����ԇg��w��t_�.�=��F�{0aw�!���I�?��4�C�� ��$�*7����Du3h�)z�lw�w1��ko��ɷ�����F��.I���$�{�4� ^��Y���qKvk5�+��X�)�wv��l��<����T���@��	��*
.��c�����J�*�o9k���fX��/Mu�g#���D��P̹h��{tc���'@��po-�<�{'o���E562 �+(�,���)��F�A�2����c��D/����iָ��� ��m׵�JY`�cmk�t�(2���<j
�
mD!+kiC~`��VY�
Ϊ,�X�oV}��lf�XO�a��ޗ[Vo� ������.�wo���e�K���w�9�3����F�qKm K�푆Q<EC���6 �J��!]�a�eK�\ÃnݜKʾ�<�qc�@�U䯖A�-g+|�t�g��;t|�h=��Yȹ��Q�����l*�e�Z�U��e��9�\'�����&:�l=��D�T�^����A�I[��\�`[��%����'tK4#��r���{"�I`�J����>v���!�k�
�t ��`�q��(]:��c@~�a6u����&�@��.7�=.hO�8Hhi�C�DH���>�����`��*��TK�k�GٮԖ�����nۜDR\��������v����C�CG�]��xڅ�>� *��y�-���I��bX\��(�w����ܪiڡSx��G���D`;e� \:��EP�4+�C���g���C��~f������<H�(����b���l�9�-��ať��2�e��[��f��9�J�K���qs7�.�<����U���+m��xGx���o���;�(�S"g7�Ekǿ��Ք[�*z��T��&�6��e0��YAJ$�~��}qL�a�.M�X�"~O&�An{u	�[)����N�YGc�/*'����B����jXqT�ʝ��H¾�
H��u�OV���:t	 ���$�æ�8U�1�{3A�f�Kk��M�	\r�[��"�U��9�M#̅��6�h�>���	HV�G��C��%f��y��'s�ϰ�i%75���y�h��;�mS�����de���p�C�`u:캓�&�w��G��ˢ���F��mH���9+ʌ�)=���W�>��13��-�ք�5�Be����E��/�����t���d^B�ĕI�H�Q�f�����"]I)��4zC��|�Y�Ư:��a��ˁc£)]-��l�w���� �g$�׮_�'8)ݞ(����C}h'��l �F�2��U���g�U<��H�em�Mv�	�����%��+F���f��nϽ��l��\�<�����j3m���'-��Ba�μQ8�  �n����T?�0�����R2�+ !��^ԧM�H���oE��J%�zYI�M( B{��/v�ɡa*ʏJ���`�i���Zl�+ѥrh�;��;x�RL="�5�S��)��u������� ��'�	�$�ut=�@��!�b�{t�Q�Q{"�����he��,�o5ʠI^����ی��)R�y-���ӈrQ�rĢ�yj��9~q0Yy&ʶ���Xl��<;4 WE�%�)S�xө�8X�7+�9�ܧҽT�R���<��t���.q�<'���1�h��{�Z��u �(��{M\;�s6���c?XG����F��:�ȯ3!!Q�¶���C�~�?!ŎL'�i�P��9O���A�g�����e�x��0��(浗���ˎ�[��X9��7�5���r�imK����?.4ꦏ<����3�����Vㅃ��W�}2�����l>��z�x{'���P����&¬�?�����p��ЈӨ���<eT����_I�~{���]@Naǃ�>� N� �0��&Ɔ��yr)�ZpgmG{�~O��?Z����p�E�&����f�O��)�Qg��G$%ÿ�c��ģq=�
�3���	M:�`�^9�����'���������2Gl���:�y%DEFBI1�|l����*�]Z��V��UN��5*��h�=L�+7D��0���G�W��1_&���y>��-֧z#���Ϗ'ٺ��a�o��#�PTੜ;@e�����jo3b-����Z�0���0��C:�����N��`��]���DF���g��h�@ZZwvڈ�]%w�s�R��4�������ˎ��ߺ�������,,�b`�z]�7} ��S�U�ܼ�F5(�N:>���)5.u��%�D��E�z�*X�c�pe'���W�:��JP�=��xϱ�M�o��v��?�?��87����)0Em��A���:��i=A���^W�,�15~B�0/�� -��ӈ����:�vBn�O`�����q��']	UL�j����y#E(R).�.Et;Rr�6nmQ���z�(}��J�K1[C��]�m�})�et��I��;O���K40
�'�7���(�֣�t��_���l��`�u>v�cAm��\n_r��~æ�f&7�\@'���w��������o��yA��q��q�ݶ/��x`�#��Xz����ik�"?�V5�.Fe�~�� `� ���\����HZ�#[�� ���E�t����-Vd��H
��i8L���h�V����s�I
�h鎟�g�"�H�bJ���K�)�y����m�E�s)>�Z���'�޾`0\ m��ԡ��!-�P�v�<^ҕ�I���o2�P[�o_�0R��Vb���7�θ�m�k�BkMc�(x�q�~e�9��p��c�l�se��U�v��E��f����Չ]��`�\D���s~"���t�` >c�3!]�+��|����z�ɦW)�'��+<e�2!?1�A��0���q1Zcؐ�ڦZ_�h�bRVM{AY0�:wO�]~�ÈN�=�����G(��B�g�8����wB���`���Şxϙ�&�E�D4������%"w"'>8|M.��W`�HSd^��:�ڗ+�;�:v���/�D�9\����YLhk(��݃�Wc��%[0�M�:@VGO�-�-�ZFlÔzb3:h�Bswj[b'g� 8����v+.�$�$o%e�x@������
e-Oմ�H����6��@��ft��f�r'M\��ް��+��������a1.KZ�,��l��#�$�By(z֐��-�D|��62����<���}�Y�f�4�`9�W�x��Yo	l��_  ���1��w�i<��v&G�+�;Wޒ>���.�B��־�>MG�m�n�&��F�.����p፤ٱ&EԘ��q�[�G�:ؘ}Y8��+���W'��+�F����*i���In�p1���@����kXu���Ӕ˦��w������z�@e�ìl�Pp�X�3�����ac��|�c!ߦ����K�7d����}�eH�H��ۢ��=�w?����)���Fzu8Ǭw��?oa� ODwA;m�?��Jr?=a$���N��f�]�?�"^�ق)1L �}�@\P!l&x���f�%�5��r�"�豈ğM�LQAW�}�M�<�������
z\=R�N?��u�U�sG)Gc�Y�ivs�[��������C^��L�;mqZ�d4�>�0'�z�+m3P�)"A�ㄮ_�c섗 �5Uw����I�УM�sC�|h��ʸ������W?�		�(O0NS��#�P���Y�g|٫'|z$��="��NѪ�ŭ.�k�%������y+q�+�])�W7d���?�W�q�7����M+b��AUǄ��e��$ .-�H�l%q���䒯�Rw�Ф�%gQ�
g^����-�B ��9�!���t������CD�/_H�2ߕ�Ax�y���qhH��l�46o���3!��[Zm�|]L���(���\E����J�kf�v�)�ɯ��\��#w�A!!Sħ/A�+��[�0&�2�h/�P��%�Y�@8ȕ~'Ě�u�6�~à���W�I�����ERAe�ZZ s�5�t������[������A�����n6T+��2��Q�J����q�����������T\$k�M����ؤ��~�'T�t��ܦ�K��Ё�T�ګ�c���.��zH
�CO���6--[a�|�'�=�b�A@u;>�_�J��{{��[��@��b�KE���e�w�)!`ﲜ���n�!��� ��:�h���R������q���p�A�3&19��SՒ���<c�~h\L)�*��m�aɏ)}es�n��oBZ�1Hv�d_�G�������8�ޟ'2������r�f'���J; ��	���X�U��|n|��4|�L�yrg�8���#�O%�4�DX8�>	��-�`�ei�z���=���;�y�]�^k��ͱ��ZL�����f+L�7���S�(��F^0��=d���1�O��L�}��~�k���㲏ְE���&n����S�|�Eȗ�r]�4�t����.K���-���%��(_���	/t�@]n� �B��wcL
n���?г�^���L�)>a`��/�9Ɍ��
"{0��E��п��K�Oú��N�MR���	,��y�q���@p6_�g���D[��:0U�g��N`�pG=f� �����W��$= {c@�h�S��K�8,=K�+������U�S��S˶Ք}�d4�xs�e���LW��/�~5�,樐�g���Z¶�i$M��f�Q=nfܓ��֖��� �UB�^��@cB��*FW�}�����.`�q9� S��Z�0uΧ�C+з:XA���v�r���D�Z�b,��R�䡤fw�dE1�E���8|�#��i6�2ózl2����IkK��a.,�ּ}��+_�jV���U�����=H:�F
��|a�ȷ��'����s�#����\G"~�����p%��a�T2�w4ڥ�N�A�4Jm��L�O�	��k=�՚�����
n*BRx:_Y���
6/H?�}���٧|���\b�њ�rφ8�\��f�8�����mP���.�7n�q�\�6h��J2j8���ʟ���0��R���9��G�"�=��PE�Z#��"�J��N �Oˀ��`�)�?��#��A�v}Ƙ��O���|3
zl���6�T=g��� �F��E).�j���y��g\���H�=%9=���z�#�~�C��{��w^���w0ޘ[b[f���_�N���;y��<v��ܾ��e��<������|���A������ �IwhA6j�W�FR�;��6�ߖ<��C��zPܑ��%Ƣ��UZ 􅠥!S���=�V�����u����a{�Qn�~GB"~F��z�l�҂�2�e���F�I9`�'��碨�`���~Es&��]�ndA����=B��L,�R_e�h1u0/�2�"�yۡ�"�4E'<��B~��"�^9��	���J�����WZ܋A��rJ�U`� I�5� �X��|i�a�t�q���f��8��"�������TI���'���v�׀�z�&�#l}����n���}�äLX�X���>h�#�V���.HJᬇ����b���6��{�AF(�*<)`�I��4�r��p��eQ�0%҅U��J��	����\������"�\���i�PӋV���,�{'��ݱvz��
B�� �'�2�}_D_�g���_�2j�rr疤 㰎㇩�p"�=��uZ�m��y{��̟m�r�����,��x�rd�W���,ws�����b��%X��/�o��B�Ƚi6*�U\C�j�=���x�nyR�����R�/�zʡM���F��C�����X�H��1n�q$|r�a"v�4������t�c+F�[t���5DDsǧ+�
�N�!%��^�|��e��m�mS�B��0�<�t`��ǘ��F�-L�f� ��ʫ�:���G{�=��{��,I˫|;���ufn/��N�ޜy�l����2�.�V��ٴ�R�;/du6�-��&,��d�q�O��=2����LN����dy��37*��F�A�H�@�t�n�j7�%x%����<Z�X8�\�w�\���lb`���@(�4r��Y��RKؠ�v@���]�����pB,H�F�����Kj�f �����Au������ȋ�3�q��ǫE�W���z!�f��h8U�2@DUK��p\�LN���;�.H`SO�X�P|h����wgyz���O�N�u�o���f]�=
��b9�q�J8X��

�s��(iW�&5�s�l�<F��M�l<
!x}�y�-}ղ���\�5k����l�J^���l�E�nN�Q��ǩ���ɤ�Z|{���A����l�E�Ki�ꋰ��/N��^�M����O�;�B�֛��1��XZ�!2�Cx|.�o1I1X�����(�'���<\���M';�W00h����l<N�є(Lu�#�H�����O=�ǒ��i�(k�b)6O�:��$!dIi��b�^�|	�,F�y~�²[�i��Ȧ�f���&��}���z�1ط���y��8�������]^���W Su� M2�Y�����):0g��C�2@�9�^��_κ{M�0�B����w�X>�Ul�ꆬ�<5�#F�z���M�;��u���i�~�=(�'6,�!��f��:�+;XO�OeK����l�(:�HB���k��v0yVU�� �tN.�-G_���9���tM�"�Yd� �xd(��ih�ӌ�n ���9>��ʻg˖]��c����i�m|����x;L��@Ʌ���f3����e�жtQ!�/�Zh$b��@�+�U�+T�-:��8b{~`��ðӎ���/�c��;ב�'S����I�BH�y4j$���mHܨ/�z���Ӓ��{��O��Q�Y��A~ȴ �z뙾	Ώ�"I�W���g���O9P���A�R�&�2'��`7&�Ρ).�r�� �>�ӊ�T��P�s���"<I�8$�0Ϟ�&���ҵ���}��[��sKDS���,0����ލ��z5)L� �j)�^�6C�-{#(�9���P��G,��ϩ��+h�j���"�#D�����D����0�얆���>�=J�Ƀ@k�O�}cv�zuS���,�6�O���d�����$|��<�]v���������c-3Xj����韃����	�,���ĉ��~$���K�p�����|�yC6�:̤�ǎt�9�	�<?F�
�G�&�&�gr\� ��(FO���.Bz�1�a��W`��_C�ژY�Uj�~�T��r�I����'�A���:��5/9e�w7Xb���L��@x��p���1B-���yđ8~�p��@(J� ����%�9l�v�� Wt�
>��㘏#f`;��������:��f�9/E�mr�6{���I�h��E�ßT������C=�����l\R	˕Y��(M�����oh9���0DK ��u�@�9�S����\�;zԚq.�h,���K�j׫�GOG��f���b��OK�X���a��-�C��dXaqt2Wp��"L}^q�~�,�!�><���wn8˴w��jT�6�f��1ezΎ�ȫٲԃ`Þ��Wغ�m�n�<`}Ƕ7��̖�X����ݩ	Z
��uU�La���ϛl;L;'�4��v�u/�U�����!w�;"�;3��zFHT�m.(�?h����cciv9gծ& D 3�<�4D9`�V}f�
�>%�	L�Ş�]�X�vX�@§� {�8������ ���������uQ��*+|�S���)����
�]:��p�����E7�ۙ�4�f�����l"��Q��\��_h5&[,e��������,s@��-�1ӣ0,T�gw�F~��ʑ6�\�Sg��@���� ����D1�PT3�wLt��t)Vd�P4�_('��QX�<�[c_�g��Q��%ݗ�	P�!��>E�{Db���F�^�*^ͧ:Slen���$m�Qpt�{}�Ur�,(��/�A7�uUQfdXH?��8��*��3�S7�>Rʱ.w �[�#>0D~t=�W�4G2塯n����"(m�W%ܖ��zW�d<�}��R�������9�R����_�`�p��0��OR��GKN��\��sO��v�a�f��8�em������7�Hz��y�ALPc`��T7�H�ر4�ߖ�u!���uI�r��ۿ��PpB#�t���IAB��X@cjT3�QG.���k�������t�%~��C�}#��w%"�ײ�����N�ᯆB��G&�)��+2�9 �v�氹�
!I�{��[� � mu�����ˑ�/�IF��gz��;�s�T $vhc�?^fN�n)5�<ܸe;4?��J34�}-�Ɗ=�5x�`�Q�=��	�ڽ������0��r� ��8RF�և$9����Q��V~sr"kK�E��;�W�`ε_9�)q�+�	9�4���`&S�	O5Qc�c1X1� ��*kć���w���'E]?����do�@ј,�����
�s����S�@]���p����8��M�����")�R��ʑ��e�l�MsI� L�ǻ�$�6�-�p���'ɑe����a6N����*���I���x4� ��_�+:��.��7/���ϡ�G,��x;�q�59�������yp=�S�x�)Ԃ���/m�%��3�鐉3��7c�l4�qV����}��Ũ�i�k��P�K��ŋ���!��W�-����d�M���B
L�+�_��\�Wvý��Ւ����X�W�:q3h���I;^��r@б:�H�Bȇ�kh1��/Rv��D~7�OaI��v�����?1H�%�G��6x��r1�����l�'������#M5[<�u	o�y�F�b[�G�#�p��%`�ԯxӬ.�<fy��nۭ%���%�bA�GdYb�!�M�%�J���"���]g��caD�=�ʓ&+Q�)/�g�����34`XC+"r�V4���Y�Ep�y3:�\��v]�e����a�~R�˪�E�u�:�-��Q�3������9�Fr���S����1}��MO�0ښ�e8Sb�KPT^|8}8bla(v�"4����.*���3�w7�VTg��s�������e�k��K�I� �*�ݷZ��`>b@�`c�xR-U�sId�C���P�T��W�G��R��aIx?!<��b�f��Мc����S�Nt�h��|r�8��%����`r�8:ѡ�.�179��`�Se�T��|�Fs���m랇u#4�.UR|�ϩ�����T��h
�?���^&�e35}ˣ�r���g��CQ�ܳ��Jg�&_��\[__���j$���/��t�����'��խ����=�#i�F�$9�:���ש 7��/�����l	H����OF;(7
1j�P�߷�����H���E�8�^�mxV�J:�`�$ߊ(@������~�W�Q�:�2�����y�v��,�`t5��ߚ=dY�WӗZwCS-����<���%��z�Q�}1�t�b�x�jۢ�d]^ʐ�UV�V�	 ��h:<���(��~�YQ��L�G��b�I���J��T&W�2��^�l}����X�<��44�����e!完x3��L�-k��A����=�����N�:�d���i��f��M�Po	j��t��� �7%1�t*s,��_���I�K�����
0��<���S�[�S���F�^��<�c���u�4�*���7"�ň�sf�߅���Ck�ɓ��q�D��t�����m����kV�0f��]D��p�e��F8�a�u'z"y�g]V#C@��RU}���Y�p���d��N�;%���z��6���oT^LDN�,�r�]��f[��G�+B҉ً7�tz�[���sI�qP�:�7z���Z}�t3E�T�P-�A'��+�������Ժ�yD�rT��OH�MV�c�� ��g� ��Y˷i)Ѵ���ս9]�A���&��.��^��)~GnwT�tP*���ɞ9O�(��&.���zn�m����\:?D+h���)��f?5��5Og���4߀���U���)�4�yP���ɶ��ڒ�����k�JH�8��Y�ήwV���V�w��{�mQ�e\�I����+�Vj9�k�d��I16�#Q3eG�3��G�o�l?�c�Y'��`yo���2A>0����A�|��ĩ,Z��Y�=����x�Jw�ǯ��eD_蒒K��K\[t�cq�_�{yχ��!��uE<�����a�P{*��2RK�!� j�b�WNG0�.X'�ා��>�*~@��|Bq�����Z���Ff��\a�rJ�*�0��TL���,���>�*5[ a ���6�&����K��W��DBz1�U��G�K~��preG2�hoSh��H�"7޴ޑq���bl8�^�x�G�t��-Xʋs������Z�o�~��Ư	�i�d�X�*�qi��`[b�7�� i*��5�&�ӽ�(5]����$�O����ۚ(����τ�῟-A#*��R:�u�(#&ȟjR{h��%�x\���FR�Ɖ��Pt�(ts2��m�/��� ˼
%w`���%W�JU��O�dFa�s��0(IA&`�E6���e%�̑N5�����%��!��ߩ��t�fCo(YMQ
;��AϖK�;�d]U��R�ͭ_ѝ�z��H���|�=�H����� T�����7���Z֐��>,r���/�)0��)F)�����_Y�׼v��<7��NR927�sa���2�q�VW�OKt��E���f=��WI�h�5G�js�J���M*Wi���m�����;Jc��HcP���D�݃˥�^7��~\�^���1��MK��%,���n^���j����G�!����&n�����<���ڢ��'U�6U�g�RR�×ig^����E6Ja��x;��$[�����������_Zf�ơ������Q���Z�Ǝo#��g�k��𺼝u0t'�V��"ؤT���7v� D�"FI�6������-�����0_�R�rgץ��['E����w]��W4�ݴ»Q0Nz8J�DZ�gsw 4�Q�O�*qڴ����!1w#x�j�;�+}����cUsֽ}�R��	�@�D�r�D��dt��.
c������o�񱬅pq�	�)0�
@0SJ���Ǡa��p?N,E$��i�SlD��J��auv��}�qߞ%�9)8�U���Y�����5�p阞��P�]j֓�P��$Y�fNb)	}БGJ�"9������G=v7��~��뒶���`��Ĥ�/���^���Z��v��m�|A�K�X�H�t�Ĝ� �Y��*إ�D�� ���N&���e��t	����u��e���g5W8���.�[gߠ�;��}6ᜠ���`�5ٳu����3�*v��Oj���	Y_��ݜE����"xv=W$�V���B������i@���ƍ�-���g�U(�>�)��Y<��rO�;��Yo\�O *9�!\2�!ZXm��b����Uy4��B���Oݠ�l(p�;��NqH��jX���ª')z]�%�g�;�����a�2<��B����Wn�qt����̱u�����[�e�4������s�/��ئ�g�X�o.i`�����db|H��
ځ� �ɪgP�KD�`e	G�s�� ,DHeI�zX;�
�"�3�|�V�'(��Fv�3%5@/|�V^�p�3#*�G�U�,���C��V����o<���4L!&�ѷ��`�i����|�(��_���f
�D�^�+���0�Hm��@�2/�oW�U1�Q��� �/sF������c�
���nҌuu_l6��b�r��`e����^^-El�\[$�弡�LM��$���ձ�U� S�������n����ի~��ŕEf"�O�M��Oځ���q~�V�+�o�p�Vntk[�rbh:��6����z��0%eV�؜^�j�M~��h�%k7Z�����PA�&[�=�2a����[V��a���"�_�K�3��z��taroߝ�Bvx��! 2w:�Dh�a�r���b�w�z���������vޜ����T)d��R�]�N�r�U>�������
���C�@Wg:\H�1H��8E���l#���+Q�K�%�
5O��\���l��ۣ��Z��KG��!��(k��l�ڽ�_����&����:�n��I$�*iA_@�-ҵ%+̈́������{��
����<8�z���&�`�6����3N���t]�_�k� qn�	�Z=$��8�xl&m�aő�H;��m��n�'�O&o��/���	q����1�H�;U�D�7@�l^A��B� :Ӏͥ=3�GKW���$I���զ7�&P���9�
��]��P��<y1$��V�w��$�o�v1x��q�|�N̤'ǹ����"��P�ٹ�~�cE�����6p��d� Q�,{�s�`\'��b�DM@u�`v���y׹I��t���ӛ�JW��S��r�XKL}�Fi]����0�]]��ˎ}cԟ�y���b�h�H���6���\��u}�$B�>�xc�<�ʺ�܉��L�0�J-�9�3�t��'֮��/�iq�f{�z�S��4���I��5J�:�+��N��)=u��	sI�]v��qP��
�T�x�����W���r'^�>7[���9#�m�����>ԋ�����o��,3� fm�� t�M�J����lKOl�V��7�n�XX��+��66�?��l�;h#�Rg����#��7ޠ�����{����[��N�/�1p|ᨰ�N�#�s4�̬�������˭�Uo�p&�6�d���� (�m�q��_N�*P�͏&����77��N�j_NI?#�u�.�U"�y��c���_Lf�Pm�#�O&���=����|6@�g�8ζ�huP43��u"}\ d\�P��O� �;H���Z�p�Űq
Ї4n��j�YնG&����1!�� qM�ڨ`x�T�/��=Ս�D��K�ۜ}f+���DWq�j�@WZ�؎n�yѠيǮ�VL�R:�ck��� \��H�
���,�.��do�9��z �?��{R#���X��W�[�$�CcInR2y�Z3Ř���?$�����kC�K�Z��Nf��`�o�E�2Olq)����jV��ˏի�q��ur��ƭ����{���������U����_afN�������ô
R���	�@}띫e%��9x�;�56đ,'��&��v�Dq��f�q�~�-�����.��IA�le�m��w����/�r����Q�yQ���[��"�r��K�i�f݁��=�Ck��X�Qb�j��w�X���v��)��_�jJ4Q�@��D�^Sasr5̹P��