��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���9w��VpL���~�����.��7
���l�g�S��N.���c����`��8��:��!�o�L�����P�Z�:\��P�&z-���,¾��DF�@��IJ:O�B$���nG��fx`x}�����N&�5b̸�Z�*���ʄ����	߈�R�6�N��+! �ch���c�qb�!��,��2P�2�W1j9��n���C�A�05�l����cn��Ɩ�Ur �coGͰ�ء�9�	�ӓ���&2 ����d/�*Q&T���	�@d�҇j�
�w���/����s�/p�,<�;�'�i�ϸj�\og̓(��X�>��y���~3�[Q*fA��m_�X�0��ϑR�.���Efg.�s
�
_FrA�C�&�A��l�u�mm�%�T�v�|o?,���y���s�!+�-�k���.f�<.�PE �lr\�����B��pW���3��
~��;4���湂���
Ռ���č�]��[���"v2�2q�^T���7�-	�8�ƤS,�ʡW9���J�p�)IR�� G�&�D��"�K�2g�j8	H��Mڍ�0�
���j@N��=����>MIˇs�=y�����hy�leGgp'~�L�MSh�`�>E���|�_��\��N��0V�=�{+*7I����Ϸ�l�X�����~f��[�*T���k�f�Eôo�@伷�;@���]N`�y�S�ě�Ȝ:09+�v.P]���[�1��	"P��O������$�:`6��!E��w t��>Wkxr��B���*o���V�����Uy�'�1$�!���v��7 �Ii^�*u��(U���I��SU���"�W�`��Ny�,�A2�;*��!��t��#F�&�F)o����ۢ���T�7_�[�:�d�:a�#]�4���k��0�S�Á�?��<��N����]}i���\�����2)��#�[$�(�Z@��huט��c*���0��'�ʵHV�:8j�Qҋ�������_s���,BP��E	5s*�b�_�I��y~��|����D�ssz]ACX�G��3�n�W��������"��8�Cْr�C34���(�:�s߬���Lƭ.&���q�?�����LY�&vL���_�)Mu����u���h_;�`��Ґ�����a*��n�v�y���M��u5Z���\	�n�1��U6b������7�ר��~�,���|t��8�b�`~`�����^=-3�n���Em�&�z��Yg��������;�ٽ��̋_{�ja�J a*������T��q����1�K�v��
���)����Fj����x C�v��E�!Zd�e�^���9{�� �$�����[��>ݬ�e�ي�� d�5���7��T��V���'��yh��_�brE������$�Î�ag�Fa3���;����: Ukzp�S�c��Z���ͿC�6�Rl���Ѹp84���u���*A�@���;��I)3���2��NH:)����Uk�"�
��?^*/��w�@�2��ST����*���8��2Ζ#9��W%�m��x�\8il.y�
�)�^ˤl�Tq����� 5!½�Y�2�	�ۄ�ՠJ�3���pPJ9�a���t�i�wmI�����K��W��G�&y�"m�N���qP�6��Rt�N��L�]Vp����=��y�u�
��T�z��hТ#ݛ;+=�NO$�%ڈ�/טY��e��7��Z��feB����eҕ�%�(��kr�7|2��QJy0�H���ӹ�x��p�:
B��g�,��$2˿�_u �WM]�����K��(��#*=�*ӆW��צ�~ 㣬��V�I�=��x�!x�B��k�ʣz������d�#h�(�؜�:�߻��D����jsd�A�N��'Jy���	2��E/Ǆk#"k��{�i� s.%��l0X�+��-&=�*co<���zn�)��7��m�{����}��B�v�ъ��+}�B��Q�0�2���X�(��I6>u:c�J�O��0G��
|b�;?1+g|KqK̯�|��l|i�r�c����K�0�
�ڂW�"�f�;}��U�2D:���_+p��'T�j���L1%M��A�&�LP��?�cH]Ko_��=6<߽#)J��G�˗��3&����hw�5���T�Og�q�|
�ų��[w;~�k��h�{��Y #j�l1�� _�i{=��:Ȁ�tj7�����^0�^M�f�P~�/[��iA�Rm=��n�m��7<W	��)�j����i��Q\4�r��6eb�!z@[��^�4��Ǣ9�8��0�|�����i_�x��iw�<��V�S�+d+)_y7Պjc�'Ν��s(��ڜ�L������۪H�>�Ҳw&�uG�co���3c3�.�������!��c����k����
R�ud' �f#�z� +.��2�k"4������ݛ�9
TtN��
�g��KX| N��;��@�&�xw�����q)���R.�	�p~�Vɔ�f�`�.s��b�~����o�w�η�jt�ֽ�����Cv���<8�>���lo���۽�enأ�\�ga�]@�[�+"�������	 @��7&b�*�(�d@�\y?�0��N��.�=~�,�XӷRn��@��ٰ��{qb{7A5R��
"�~˥g��d>�܎ "IR����a���i����^�Z��8jF`�,`�r�aҜ~�P���!��@���}�߿s_�*B�;e� ��z�`���|���qhЛ>	�4ܵ\�aF濞�]�N4ڻ:�"nF]DN#N�8���T�@��_|�Z�4�992ۓ�zVFg��Ȉ��M�ja��*�X�f8*^y�0��<Κ;)!��L�ӹ>���c� �Ӟ���Y5���Q�E��<��9�E�B�"C�*	iT����B�S%� U���?M]-��sJ�NX�?$T�>��ڏ`@{��G��١ZtH��簧�)6Q�O�;l�n98zR�G�$�ې������{#��0*0ة�A���O���_[��?O���e0�n�o������m�f�����1��8�e�U��S��{�V9��.�&�f�+�,�@���Q)��ƥe}$]���y��
[|MU�bL�'�*������i:D$�&(T�� ���u���S�;ծ��Η�Ӝ�5hX�q�q*>AJ�F(vn�T��SYma�/NQh�I�G}l7B��C�V.���I5u�vړ�=v�}?��m�̩O]�N2l�5`]$�O܅�s�^[a�Z��*{|��H��Yp�1�h�D�ӂ�o��E{$��g3�"�|C��(�e8t\%'o��u�sR<[�jc����D>��Jߊ�\k8��:�r���\��2+�#/�d9)K�>�!Β&OM�e8�Q�lJ�`
'�f;�c�����J��L����kJ�[s2��2�v:Ѹ\C�.�=���jY����� CΩ�F1}٬J���h?j���@�� �y� �n���e)�w��V�Q����ůư���q�˕"�*EP��^��Z�1w����P˭ѭ9_�����+��������&��%�x9F�*+�k�=���k=@S�uB?�������t
��0e׶�%��R�&&iǔX���r�f�P²��m˝�����Y�k��Җ�*A��ˮVYA3U�	"�+�%���v��Fx(�c��7U���~��}� �O�[}f��t�cU���!�u"Ho�,A2���]>T��Gvs��ࡊu
I��/��$��?��+�.v#፥S����7���`�"��}}//�S���`�3�~� �q��>e�bO�������/IJ8帱a������dzJ���2r�洷i��o�g"��TlG@��v�N'�N	%���2�T�ܫ�>�Q������MtZ�5�-�y����4m�ҝg9?K��d�@X�N���X�'��gκp�{�u�FoF)[��:I���4%�5,���#�)X�1���/��ԛz8������tc8�_���SM�}��5g�?V������A��S�L�WuZSq��M�gu0�	>׹2��si����|ׯ]k���=q1z벎c��xTj�Wj��}��g��dn�*,L����^pg�yM~���V [HrZOe�"_S����]�{8��بVz����{%ϸ�R��$h��mFF�66�_2q�lB5�cʅ���Z��랈,C|��77o��E���DT��s]%>���m�s�X��y�/��Tg����f�
Cج�f|'	L�ܕ���G��+�,�:�������8­㝙{.��������W.�ɶODH�$���+聁��JZOy���>6�3�.'� ���i���[���έ���h_�+&��y��
l5�t'�2-���=����j��o�?�A�۵w�Iws'i1B�����%�Q�cq�Y�)W|v,İ$)/<���� �����|����VתP�Ze�G�ot�MR0�pF�����\�D�����f��C���X蟃�L�Q����
B�H��0�yN���W�O��q��s��tМt�o�����Ye-u�IG��)7X�p�YI���KA��̴�Ϗ�G�'�bG9�2$i}b��j�\̪�:��o+ K�� ��C��\ġs��|q���)��\葋T5 �;�
��@]������u3Q�:B'�heB����93��#09��zU �e��H�J�>��R���q�;�>Z��y�I���1@lu�A�{���E�T�uJ�:y=�Y��.�`9�b��غ-A1/tw� =�Q�(5��svwu2\��O�i���I�n�[�5��gvE��[�+ɑo��f�"A��iClU������8�}����&js��dUZ��V}V�=D3?;�$���YF������N���y�?J�_�}�ΥΆ�ں��#J9�Pu�-g+�T�ڌ�:lu7�«��J�ݭq�jpȬ����@�y���R��.}�Av� O�C��Y�K��t�EOzoy0Mj���/$)J_�*(0���u�T�k�lU��g��v�o�29͓�5��L��.�8Tm�]%���=���IfU�9G����E����.^��M��aி>�(�y�d%i$ܖ����ߝ�\>�1F�c�1�]�qOf�c�/�r��Y|\����G�{.b�%<1��-5��SHQ���Q�є�"�JVŝ��$�T�[*Z�qֱ�E)_�:�=ӽ3D�Z��&}L�'e����t]��J�q�� G�9�o`5�|4l�����a\�_�MW	=�,c��b���%�O���[��L��5�W��(�R3�n`y����.S=Бi�-��F�;��{Qi���-�C�Dn����}í�Q�h����o����IM����5���Ұ�M�۽#�$%[����J��6(��d���&K�䲨��F�r|-�cކ�&}p�e�zH�x�� ;�3Kq���X���5���N�"�T(��!�+�f�ԁWe�s�Q�N���_!��r��ʾ�e$l�.m�y����vQsۊ���I�ܲ��cۇ�� ��4��3�5�G�A5��oeq��=��D�q�u�����Å�@T��HW<�ٳ�{3>�uK7&b
tuxF.��M�����|�+���6�p��r&�-�{�TY�������nJh�eoS�;T��1ވ�L��ׄ �9f���̸�)Xv�]�}��&\Yr~��3���q6;�9Pn�;�
�U���j �����#�؍�9б+)�G׀�M�{R�sh�~�貜�J3,���^��s ?�"/���F�uu�k��Q�j�b6��4��1A��j+��w������(Y�����[���"?�OY�v�>:s��tٞ��ɣ.6�*HK}�X��|�˕���Q���	|���*�Sxns�����I��2������.���AѦ~��c��R����7��HOC���\�t�����16��vV<�6=��t=�h����	��0J�	N1/�WxQ.,gY:�Ȗ��d�0����Y����T�/M&�w��&��G�8�[��������:暎J���h"���I��H� */��W��z�W^/Ց$�x��13��*R�po�=��M�e��8'B�h*����"�f �7)�@[RS.�ƿ��f�6���{�͵Z���I�U��UJ�c�vRl�����'�F��jXDiī�$�@_��4����](�	�S��A:z��e@Il��q���
�ڮ�Y`�e�-mU�b#d� ���|(�o�F�DL����.\I/x�6;N� qo睱'\Zy��sR���,���1ɖ������8G�7�>���ߗL��d�.��@��G�7�3�>v�sUm�SFX�ET� �MIh���&�BRͶ/-t+�C
�b�}�#GƐ!x��͛ ���'R9:��v廊�B\R����;n���?`���	r�|V��}��oz�wx��9z0����*k�I52bg/����On
k�n�KNUI�I����Y�s�Yb�O_jl�����%h=�3�4�o)8��un�R��|
T�|!�OO�R+�o�7'TO,�{�z��0����4$-VqV�Q��s��LP�N�)]8,h����Y�	��	y�eFQ�ؚ�&Q�h�5�ֵ8��q��`{ƿ�<�#dBm����%��Ǣ=bY7F!T6�jd�п�h  AGvT<�6oʌ�-�|<[����3�.	�@Wt� ��bq��=��ͯ.��C�&Vj�b���"�9�z�`+�Cd�Oh��S��K�-w�
#�n�%6v��<��U�_*�i�&��:F�`E�ȑ���/�xM�~��Ng�H'0zmm��j�9xRSZ�<�O�|2�,a�4&N��l|i��W{
6J�4�h��sa�M�m���%&C��$Ό�:�}]ա3�%�r$�[���	�+�ʚ^���_� �l����[k��I��b����fC��/�5�m�V�i��@�^����*�#VR�j�e�#H)��!>_�A��;�<������@v=]23��.H�ܠ������-����z�ӣ���g�[8��em�ݸ+)W"J��V��f	s��[����Pwm,�#A�HZ�C��uߧ�*�F����uZwH\�Ǘ�����P�HV��]f1/u��T9�W���$\�>�<7W'��O�7]a	(�4��¨'��U���Ug�g{fM���nq(e��P�O���ڻ�'p�W?�j��^�Tx�w��6{,P0�,���B�Z��ZFKp}�`̜�-��I����0?��q��U��P�&�H97��vN{D�qW/qXW��6�͢kD��͸��m��j��W���z3$�$����sjX�+��61�.�����6�Hy��=�(d{X��d�/�}���*�2�־������%� �f.�ɠڷ��F7���R��K���"Fx��Z`Q��*�)�NK?�B��T,>6��T�Oޘ�����{�Q~p:�żq�5 �_�#FFF���1��'�`�;����#�g�g梻`��󸉼�g��i�L`��'��}�2$ԙ>rU�	�� W͐�����Fg�w�w�bF��Y��62b�ٵ�^�}5V��\��I��)Z� �m\���Ub7-�� ����%��oZV� xMv�23�AI�z>�m��2�N�F��&����߇M�Ԯ��}b��\,õ�
�ҭZ���4��Ƕ6�d3[U5�8|B��~:pY43��TA�f���d;�V{Ў߄�^sZP���. �{fLqig�LJ��������eY�p����s3��A�ߝ@؅��J���^�Dvy�g84����'�� ��C��.oD�0��`�B�y`�Z�z6�D�J��璚i��C�q6"��0������c�ğ)ߚ�z�G���k%u7l�.c^�
��I��`�y\b�����W�pZ�.x�޿S��NM�o����h_s.-H4����v��H���${�;��!��7��7�9��HY8�Ow�%>}���Z��.�X�M�~��53��_�`�N��3�e"�Z�csQXw���F\��
�?������y��8`!s���D���߫k�]G�:���>��Q�vh�R�:��u�R�͂�3�5�6;��}]�Tb��ZD���
�C6#N����:6��"g�&�~ɽ���Ɖ,���u��4`NT�]X�����̤����~��߭�B�~td٤YB���*���ژ�m�U'��T����4�n0L��kc25L�����3�Ըm5ݺdU;�!d{�V���o��Wf`B�b5��J�P�8�����;�<n� ̗]�nS�BG�9��%��%�h5}��J�"�J�F+Ph�f�U�R8�dz�Ԩ*n�Q��3-�Y� s`�t.�G�n,�^#1G��Lȳ!'�t�����Iz��N�����t�\�e����}��E_��=������{w�Zn�������n��fr��Y#Qנ"�aU�J��º{�Ϣ`�{]W��p��e�Ϡ���������.<��e\#x�q�'�Zв#p�S�{Q-�D�E W.1�#��	���}��ɯ����h�K|�N�����1��a �B�K�o��w���2��'R#=���V?8�d�_wu���qb
K\#njT%fg��)!���>��?1ɕ�ds��Κ6G����-X�ގ��+}�bA�N>SU��u���O�NW���Mnh��9�]�f�e=׏�1k>x$ur�5�E��ݘ��;]<75�S�ԟG��;����(�(��>��~��3�#��?��8EH����n�٩������j��z��]F���Bz�D1&�A�I�5cc�9��D�Kn������g��NF�so��>��s�x�����T��:�х�
�ؘD2Ą�,����w�L@e��`��UlW=�إ) ��NZ׷[�U�0U���r���h��L`++r=�8�Q��&2��c�
e��P\�Ź%Z 0`BqH�b�5�ʾ�!+���V�	a��.d �]��\=�$*k#~B�P�Ӂq��-����=�pv5&����ܼ��ҺBx���JR��p�I	�Ǖ!t2����- �v��,m��	���R�H����v�Q= 猀����o}>�̀�g+p���՚��aiٔ�0� ^E�����=�ܞO'-l��k���m �*QfS�)��p�ǃa��� "q��Y��0��ٛ's��WӾR��0Ѣ�51���	��#Ĺ����+x��/X{�M㩅��dOM��́[�A&.����������bs�SC��b�}���a��5rɄ�T�f������$�tx�D_K֫���kl N�H�����ۢ�׈n�D�ɦUJ�v� �2�-a�T�̤6f�
�����1�.�)����AI(/3d�07��p��z'�)7�����Y�β�Yg�q��3��|�=�m�&�/dV���������#�;������d��	b�Q��deV �4Q'�PqI��$����X�D��[ٯ���)���l�I~�;��qr��G��R,�`��&C�䗤n=?��B�^���I�!M�_|��j���g��^<c>)��#Q{H[p��H}3~�`�DUn(��H�Z���u�
�<㋘KS���d����n��:�wAz(!
7���vP��Om��������1~�(���+�'�[>��6�4����G�ܜ�s�~���zh�q`��dkYs����n]T��'ѝ�~|����$��9�i��K/֙��������w��:]��1�;ed�d�5��[�
~'�a����mQ��jaE�;r��,Υ�h<%a)]9�׶�����ݕ��qv���\n�9!�?�[L�&)��<��%�u[+�~o�˧�a�S���PC-;��e��ug�`�8��h$k�O>�����0ÿ��_(6H���M4�����dB���L�T�¨&x��c�gX��/�������lE��߃"���^�)�`�L�Vz�_ʁ?~h�6b\'�А��kZ�t}I�y9�?zh���پ���{a�|nxd܄Ր��5qKNn�a���Μ�[g]�O[}�N(t���Q��s��R8�@�m��DT5�Qѵ8�>�'Z�C��_LY��9	X-�$�:�G+��9F\��`�6����Ae�VX�W�u�-E�@M;A�h��F�V�c<Le����d�i�G���k�k�mU;��^����*�*TD~�&=���*�,m.j]ތ1�!��	����loxE�[$�Dd�s���B���/���5pk*���-���8��g���`�L��ϤTSg<�p#�9���1Fz���ᓶ�6$�t��a����N��V@��5_ڳ$��K��D�a���*�}o�x��p�>���<��Ճ0nP�m�2�<'�]��_��ܕ�����Q� ���z��Űg�d���Z=�Ǻ:>\:�*��ݯw�Uz�U��4ذ�w���a��@���9�j�|�1��|����\k���/��� �%�ܳv�3`(��A.�D���(�Wv�E��B��_E�f��?�?�n����^"��c6�,��&�n�^��m"������/���rљ�F�߶\J�Z�ʌ'�//d� �
�Au��BlvilS{<80"l4�;���$y�5�ε��=|��N�viFW�%��"	�>��7Q�i�D
��e���v�����V��d�ikgU�-�jvu�jd�{`�m)yH,�۰�����2"!r�����A����4j��>�֠� �	'e��U�����Him���!��������j0_��]��%���T�U�>���ɾo�Szn�k'�Mş�UIf��������{�/�(I��k�h"�i3��nJ�G�G�"�/�d�|���g�! B毸<iJ�Y��C�eD��8�x�a��m�i|kJ���9��.���c���C���2F�D�Ƣ���JԐ)��\����������V�c�����6v������(:g Ac������t������L;ˈ��+<��c~���ǃ5˅@�')2��`��c{��uR<�X#I+l��G?5l����T������H<g8�ٿ�U���--��J�a��z��$��%��mM��<J�Z��8���,�����i3�I:�풮//�'�C:e����|"���7���xa�}4%[dl��O�p<š/p��U�.a��e�gp��m6�?�T
�"��� ob�%��_PMY��ߚ����D��qY�GC2d�������ONV̫G�"F���sy�ڟD�/�Я�Lt�K�L%�9�.,��_E���Z��`{�K.]�`[Awm6�6��m�nD� z��uI�j�7�H���K�	q�0�@nX�iz��aȊ�� x���=����XU&f~)��rdc:��I�+<׸���˄D��u�-A�0�H�H�UHL�qf؝蠮4.�>�p���9>^����ʙ-&����TY���`]hxq��>�ω��P�����2����Z_?��S���Q^�E�.Dm�C���a��q<9�P0����[O�7�)�����{~���خ��d��U��t<�N z�w��x��� �o3$�l>)����u���.v���Ϡ�	�� kXL^$.�Co�%:g�-ؽG�򡝬(����"W�����D9�Q�aZ{=ߍch ]H�K��Ujv���"�-��IZ���m�5�%�� &�0䫰�BJ�UQkeqa��3i�,�y���a_���7\g��T�N09y�Қ�܆��?��DK<>y^TgpgM�x*�~��%��H�>b:�׻��g��Ӳtc���);:Im<
٠쁛��M�K�e,�@R��gpc��������,��R�m��z�l�E饡��0i"˲��4T
A�����I���&o�:T����e�t��C�t��e�i����$��e����"�e�c З��e?9�K�Β� �3�eM����4ry���g��vVpu�m^��k���*�	ˍ���D �/穁�l�UUW��t,�7+Z��qK��ip�%�\F���]﫻��l����Ռr"�
*���"�q!6/�ZWcF���e��,�T���n{I2S���rQ+;�Si_�9n���M$~Na���ὀ4g �T�l���Z4��o�c�8�P�aԨ\+3Z�lk�]��Ej�ދ���*�Y��N��݌{�؝)=BT�Y��4��ط��B��ꑀ�Z�0�F�	���?d^M��/G�IC�T��Fɽ�q��B:�~\r�wiqΥf�R<5�,%�����|�i�+��혹(�B���Z[�ϧ�ł���+�I���q
[
	�nɴq�:�}�X�1 d���҄�����L����\չ�*��Q����3'�t����n|���9D�40Q4�'UGJc���0��H8K�d^�>w�AI8�j@�,�/z<�'������
<]%6
�op�3�a�u}X�f����Q��q�L�ki����H A�ۤ5� ��I���>��i��<z6���마H@�e%⩴
,2��"�Km�T���vJ�g�th�Ո�\�',	 ,K%(�7`F��wd�A�Kqxn��yޕEP�(2M.�+1ҙ��D]N�	r�D��Sq�R�a�!�n}��	�Ӥfb�L
<K�d�RW�N���0<#AG�Ŀ���,G^l�y�3�Q���e�Ak��ۣ=��^��1�2���B=���}���$�"3�u��m��i�k�y!H8~�c���Ǐʰ&��V�Gܾ��f,�BYU�s��k�V%$���e�ݽb���;�X��lh3Z&�A^ߟ��yG��x�̽��!(t��x��4ӣM�[��E剿��V��[Χ�C���\Z�� &I�~��b�2�UVu!#Ll��&N��wa}6��$�:��[ !h�V6�V��N�L��>�{����c�_o�����댆����:<%t������X6w;(���dқf�M�t�N���h0a��u0��@S�t��+��<�T���:��1M��"Ϝ蔯�ho�AO�>*1#d��x���ses�)��_7;�In5H�9�m��bi�:�RP�M_��u���F<N)�C�=��)5�=QFߕ��J�㊨</���K<���[��5d[���U���������M���j~j^i�L�[R 9��Y�ſ�	W��،��Y�tR�F%�d�Π�ׯZ����7�N ��*�:�4�H�_!�U�#D�.��@��ק�?�Ȑ
� =�$�4���i��ٽ;G���Xv)ز"(m�JM���d�_Z����Z9�G����?�:������T��"&���.F��miΡb���z��?L���|_�*���|���Pղ�-^͌n���aUUf�әˠ%	J\8[���:E��f|S۩�:�@�kLLS��۬+�� �M��@V#�4�1���垗f�z�O�Y�0��О�W<��h��ı!]���>���?���sID�w�&_@K�D��'K�2y�9�W"k�yUq/yK�P2����ٗB���eg��`�ܫ̯�����$9�����.��v��!��ĳ���L��I��V�:ˠ��`ņK�AǞד�e�M�4�Tݗ/�/H�ur�Z$
�����1�ȯU���g��("}�+v�m���&8�O�Tql; w�0 �Z�A7�;�DL�|��Q�7�h�~��ʢ�X��9�(m�j�8�kWxn�|�k;kߞ����l����Y>]�FS\˛�{>��"��?̑����ٓ0� ����q����@}DE��O$QB`�Vy��=����%�pI+6���Fځ�ȵ?&TZ0�z/�_!�|:��r���.�����(Yr�8<Y���ٜ��Q��S�M���#D�Ȝf�n;ֹ;3{l���ͷ��{��5�"[�E ��N
�x��|�o�}�K|��� ���(�gg�P7�}M�K�4
+%��Z]�^�a��Ӆ�Z]Y�a�z8��H�(
Z�z��Dhr4=+��0��p��Sɪ�)<[6��!��&�G����gA�m�tߣ4Tˆ��B���i؆��}�ij9{��m��c�V�����W`�����a�;���[t	�%ܵ���R���s)�/9�(Nm�����'�S!�Jk>����S2�t�r���-����בJk
���� U�y8 ����+r�)DB�{2m-?"'5�Y�X�����$���`�H�7�¯hU�ٶ�IZ&P�wsٔ��0FXE+I�?^�N��O���
�ĊELY��{@�^�ܵ(t�ȼ��x����m�c�@�>)���]�@Á�@R�d�U(.�N+�M-�x�������{��2BBG����q��Gd�I��b�;F��i�$��%�TՂ�$�hD�h�����p�sv�P�N�
�$A�';2�C�v�v�(\{ 2S� Ÿ�W���L�}�z�>QT!~����2[C���.�r��`f��ݻ�7-�J��W	�h�@�i~{
/����eܜX��qW��EAO��O�9��G���Bu>�5i��p`#��I�# ��Gh
�#]��d����hH/˓j�z�@�*~�(������Ÿ�Gc���H5���4�
�GK�Ra�1ºe%:yi7�"Dj2�۹�������<�ɀij|�^A�9�AΗ�KE�Ƥj����*���LE�*hD�a�U�/��~Bb<e�܍�2�R�~������ϣq�n�i�РM ���3Z�]�v��F��I�t�dE�_U[��|e�10�92lfHX�=��͉Ri���f�n���'}�Tִc�Jķ$���g� � MFMٽ���j6,�0ٔ}�L�㗱�^��S�[q�q���W�O����1S�Ӈ2|�Sg��Q� -�i��A�EC'}2�Ӡa�8�Q�V��x��d/�f��F6Ē�s�B������&V��S}�]I��Ț������HN8�*�U��DnY����)��96I�Ql/���܃�ܵe�g����f��0)�S�t��فK��� �~K��5�uv�ܚ�����u y�ݑ�jjLS��^h���H�|]�=�x�ب��m@!}��DR�7'�	4t�ii��t�w>�M��}�'�(]��BK念�)j���8�C������
2y��axxl�R
܀U�e$�ｧ#h^�	�=����g���_$�15�a0m.$%�I�5'l�Z�@B��t��6�aE&OV(��`���K�6����{�[s�&HN@�\�L���X�t_�Ԋ�1�/hk=�s~(5	�%*� ����ǦY���5f&�s/����*^����,�3`e�%Bu�b��+����e���n�W^��X>��ؑH��e��覬t��eN�����	|,��˓��ܛL��������m����xz�1Mڑ�X����^*i�w��d�%�-<�Gi�?"rr)�(Ⱦ���J�� ��{9L��1r�CDA5F�!�� 4��&<-��,l�}��n�C�2��C]�-W��~���D���� 쵃0q�d�axOat��_c]6jE�5pjv�4,�q�Y��p6p?b���}��SD��`��[��'Z;'��lo��MM�S���ԇ��"ޔr�7���%/�õ���V׷2�-\s��v&N��VdӦ��_=�g9�X�SdB&Ʋ��d�"�+���8�UU���^S�g�x�Ox|[@>W'��=�IS���?G�}�����0i�#Y{����0���P]�b&n(�2t�U��w2���R��K��:�Fqǵ�4��_��ۃx7��;�f��Q��nD�� �������/P���L����R��[��
�9K�G�fb�W�f}W���_��jt�G�O��H���=���D������.�]6��Z|k��Ū �*�˙�7���a�������(��()&pK/�,k��JM��Jߵ�<J�ٲhZ�� �T�����z��Ս���:I��.g���tX	���������E9,�e��ET��7f̶��j��ĳ���i;�2�I�����o����UOI~W���"L�PʸG�� C��r7�N[��HK_�^�D[�}�mo"E��A�P~B������!M�]�ى�������u>$�sx<X��9?��J������i��`�R�n2_��s�Ҍ�̆}�'S�TQ�AOdAw>�i���Z���|�o�0	s��PWQB7�_��x��3����p�1~��j j�#�5��(�j��1s:�8��u���8�N#\����\�F*G��5&"I��*�ša�'��l&��r�ᖻ�]L< (��oJ��LΩrp�I����{];�&]H3;[tS�-d<��[�x�.�p1�$6>h��&؛�:}P�.{�*�m�<�����p~,�`�?,�E�͘�'�K$�;��"����
'��`%��YX	��@tIg��9�!>��WX3q�� ��C?���thDs����Q-�>L�z��j����d�#��x!���1���Q��e�|
I�?����Z^�11��a�����n@C����6� u��.螿B���v�o�E�{��?��W=�T^�`?,x�������no7�����g��
UMx������ى��1���z��a�3�p���i�\�.լ�W���-Wd�(����a�����{RUl&W� =���aR���vM>Nh��7$��l�L���4����|���3�q�S�
�[j��w�A�~�M04#A8�뽨��7����_E���MzBi�X�ASS�7��j��^��� 8�kL��\����,�kn�o݁ݳ��^i_D��MO�� 
�i�-���&$���w�
gWY��9~����9����z~(��4�uX:XZ7�/z�tyq�/}������	�.� N�Mh�Y���(������u�������lFD9���St�����c�,Ϊ����}R�'@��v��+q������3B���0���:Q�N���s2�85]D"����μ|E�|�(���@���qQeg��ߑ����m8.5�-�`��j:�;�6��i��rM����T�#I��w�wÄ%��YCo��$�MqTӴ��*n�w���c���	_�z���} .�e�-t)Ĵ{���*�k,���݁���n�A���f�����}�?�,yߠJ�KZE.#H'5���t�LHy�Vy@�O�8:yI�C2A���t)5K���`Z`�֑RQ�|�n�?2�@+Z\�*���X�2Yk^]f�8�Dy2����x�Ԛ�kZQp��g{U���!w��WU�y��e�O�t�,8��53(�S�G|�)^э�X��ü�b��M]�����7�d�
[z
�|׉��ט\�I��fq��y�Wx/�
�+LH����ᯠ0r��q-���Wgl?de�0:Y�k�k��B�o��(�ꗗ�o��s�X#�?=e��� N �F<�<X�����}}��D�p�;�͓���������}�&Hi8�]���6&��gw|8��2� }��&�h�	Q�L�=C���(ī�
�5���6���S�:z{ig�럭b�)��XN��XS��ad��6���t#dL��s�~S_����ШY3gU#KR�؃�b���}���Wm��+��H�Yr������5�H�*m9�o[ tB��ay��<=�!�鞁��7Z^Q��,a{�שW1�@��>+�Й�O*֫���&��y�TGW~����Ens�ü�Na]�n��y��+�0��3�z~�#mگ������;����vh������f�k��?%Q�)<��dr�y��r��u'm�mq�V�I��>�M�Er{kX�p������ �/�X	ܷ�_�ێ�7���X�B�Or=����(UUn�9n|ph)��z���X>y��{8ۇ"� A_��#1���;&��}��
qq��H��/~��LE�`���|�C$a��V��V�՗6�������V��_���(��s���"�b�ַl�Z�F�Ҵ�g_���'���RD�NN>>���T���B�fy��(�mt�aΛ��?�,���%1:��[a�b;�Bz�p��6}����&ɛ����+��|A�UĪN���w�ԷO�8@��9�'��L[�R0���-�<q��N�<&(��3��"����lL�U�p����p��n�LV}�'�N�ߨ��۽��}>��f;p'IX-k��kEJ�����Ǵ�>:���Hf���m���)��S���uL�A^���W�M�����ӁV!C�e�a�Qj�
�x���:��[P��h��3a~u�H:f�8��5�����P��IN����]��qa��f�_s�x����<�y���Ge�Hi%U�
>�܌\�-�;���Q���_����a)���%9� 	RdX�S�K�����{���L��ia�mhrZ���0���KDX�p\~� ߊ��5��Ei����,����r3�x������MI���R��Ӥ`Ug��k�T��#�f��HUW��� 1�K���>�ҹl˫�]`����V}��v/T��D����,�_�ti��MQ�)&i�q��e�Gn!�:�Ě�\��ս��6A���FO�+��Z�?���2^��Oz��k�.ء�	A{B˰#LK.d+r�����0|[t��7��/�����Fu����^���"�������l3��U �fJ���6���a��0A�B{�;��&�R"���F��,�)y�9��x&�FBU z]�$�S��v�	�F��E��L̛�GRd3�#9
`����t�����P;7�䴶7u�Tsf������K�f�r� 7�f��6��s���V,��5P��q�:�)��$�F/V	(��3�P�3�t���վ �6B�7�E��������btK�F@���C�g�Œ� k��^�XH𫇋��^��T^����$$S���bG�l~�Z��C)�4텸H�s� �����p��� ��8������7�8L2�|��>|�y�)2P �2_)��B����r.�Ѓ}В�¬t��q<H��A4�-�T��?���MJ�{P��'��ƶ��"	�8f�r/�ه�.]��
)6�?������W�:L*��y�#'=�ƞ��6��]؝	D�暖K�{�����˓P\~ó�] 8�DqS�_��YdR�/u*�a�ȃ�=>S=zfOH럱M�p}�!��SA����Ц�����=�o�h�P۲����;��-���p�?h\TS�̵�xܶR����ݯ]�F���C�����
��������#�ᅁ���̸�C�L�gM���{z�#@�VN;A褩��Ov4���������;�Nc69�3�X.�8A��5��(� �� ���,�'���qee��Q,��~W�D�MQ޸9w�૝���U9@�^��'��4KBߢ<<C�"8�π��\
ʢ^�NY
)����s:�Υ��$uسmt���e������`�m�c�)��[�NC]2h��G�ʢ��8Ѝ�M�-0B��|2~�ۉ�w��@&�no1�=j/�S��`���p�IH�~=������1��)J����*��?��r�Yo��|%W�Mhb����d���-pO'L����9�Q��L�s��ǺX2�Z<��4�K��5`a7,}>ύ��V65k.iu8����_*�*1�W��I������kt��G���6(�u���Y eWA�Ő�}� &Z0���oD-��<=�f<�Й���>\�#�g��] �*�F���c$�o�Y�1����?�:p%Tz����"m���`�@&W,bP�yܤE��V�� �y��z��`�U���ı_��
ӕ��\U�2��;�,�t�u��c͖�lqP/�����q$@j?T]�� �Y�!����R?�vܦǈ5��'Q����x�c�h]���ڋ.����z%����Q����]��� /Z��2����D �V�;2��5�Ĳ �&*�=����7�菖���R�B.�,;�X5�g�9�� =םe3v ���Q��N�3>.�藡 \{q@ۡ#��l����H�AC��#���vt�y^GP�_L(�|�)�~�0��l��<w�Ã�~E��o&{W�G5O�J�=����h�����W���%X-��x��oȥk����)��",_���*Y]�F{�Q�`�,9�O �Y��ƶ�	��|�q*��"�#��D�_#9����{�����"9!�Ṣ��2�	��bQGI#�A��=�H�7!$�H�p�ᄑ	�]��d�z��yg�^�`�v LȤ�*T_�K�R�u��+A��3���]�Ɉ����"�r姻J�����6�vcRu$�(��=�-,�DF�p�2O}���z����m=[]�\���R��Z6ϡz�`��;	U�?E�Ӛt4�U��J��{�?x�yw�ǹ�Zi/i }��2Y�06��GT%�o�@c����<����~�i�tb���Wq���� ����۾q!f	�. �\���d/��3�	ݾ[�^�ҦU��YrK���������흴�-�"vD}V�G �tE-��)�Jۖ��R�VW��g<s�e҈kX�����U��<4�Ή	v�v��|�� ��C�HⰣ��G�Eښ�@��Ǔ�V5�6�:v:& h�\Yq��R!R?�p�in�v��@����ѣ�_K��rS��7����ec��(�aX�16L�+k���m'љ)��[��{�g�w5�;W�j�Nn~�(�r�,�t0�ZAL�Уh�n~Bv5@WV�@\Ò��6^�9��;�{��z��VG?��F���q�!s�2B�����@G&��rɶwt'�O�kZ�諃c�@s`®5`���p3�������F�����ӉE+���2<:�n&>��\�^1T�?�@DQ��a��p)�G�ٕ�o�<E��Lgd*f�]$1ɞfQ�d��Bs�&l��nV�JFD񉘠z>������?_��_d��l�gX��9ݗ��ʒV�4�=u◁BɄXe��%G��j�%�b�Z��jH�h�.�_��-^�b�.P>��]e��|ʷ�oh �Ni��xժV����g��<���{���K8$5�d�����B���P+���{f���k�l3�۔g���>��yCJ�������{޶�����%�I����^�w�
�D��8����F{<�Ч�ƅ�^Z5��/l��mla�3�ć>fw-$���G'Ɏ�,b���i"�6�Ay� �D<&�L����qpQf��4�"�a�61���w�Lgሥ��૊ǽ0�ئY�?�N&���dJ��d���(jWQ��"�f�+�q���ѐ1���S9����D���c�
���:��kU���Ot9�XE�w��	/�wA]@Vp���p"A�ҖӅX��j�%��
�����<Qؗ.`����v4U�n����r����b�B xv���u6$���R&먟&�ݣd��Y�_wV�
e�$�$r��1C��������M���$y�k��1��������� �e�Ⱦ� u���i�dQ�dX�fP�����]*�v�,�9(��~E����\'��h{(>6'��q_�N��*��"�.4�{:�� qy+jS��S%ʆ�"�n^C���",ig(���?��@�-N@��F��r�jhJ۰Zl���lT)}&nO�fW�ǍW|�3�t{]�h	)�G{�}m�8��Ï�{���B?qm7 ���d�5���F�t^0}J���g��稩�JS��#�
�D��:{�]�t�N�8�I}�vڰ�_E]òs-[��p;~0QY���N�s��\Ζ��I�_b�=�r�L-���7��R�%b >���w!��H����<��)V5b��!�/_5��������Ȗ��g
��lm���.f4�QU�#6\ҙ}�`��w�=���ł��M!�&m��.9�Q�g&�C4�>���=ߥ<iTe���5a��L��u���F��e$iq�FU�	��CF�x"�l���n�>���8��+q�[�.`�`�5L��' �)V<^��1������ȁb|B�P0W��;��ee��2���xp��{<3'�{t#$]����.�)T�\��+ԼEҺPl��oڧo�8];p��2���8VG%�M�S��l�,���͞��s�*�tؓ�@?��S���;a��������͈�>��N^�)������u�s��^�����C�1ܦ��9�I��'4���D��d�O���b����*��-ԁq�i;/�Qb6�s��P��Pe�F�)l����FNt/���D��y-�>ȱRD*qO8�D2P=�qU;�\�`����O�~q@��,$>�:�H̵��9�pe7��U�B���wY��Eq��z��wZe̈�ʠ!�n;w��X�8��x��iD�(��Q?�~�6qa���j������ʹ�Ē8�[A[I�C�->��C0^���AL��;�;�'{�}�ֹG�ҙ���_�z��o@����U$l�CCUݵ��-�,�]�yi�� d-~�mk��4��ߣ�4eyO�N���_k+|�%�1t�w�d�����P#W/v*"Y'	h	|d]���*M��`���@��ݓX_�.D��y�>L&�����>� �xt��hs�FP��~�R O�I��^��Y\��p��N��<U�'	�3#�{�%��d�l�	2@��xn�_����V�V��b�@��V���ٺ���&[�?��0(<�u���*�_n��P��9�����{�>7㚨���c�������Dh�I8���"#�=�������}q�vxʶ�ՠ��:���z��DH=��{׫w����鰺$�ci��&�Ruxۍ
��^��/g���8��(n�G�Z��@� �
���� 1=�p߻e��G��*�?���h�EO��垞L�����������������!!,�b����T�b.t[;F���zn��<�A+ӆ i�P���
�W;�#�v q�T�Ђu�������$������k[�����@�(
h�������fǾ:�"�a����RH K�;;���Q*LxI�ƝZ�r�4JR<����NwS&�o�y�B��p��;��E�NH,i�MU��8������%����|�BІ�U� ⠞9&~B���5%���d�l]�Ga�=4��cw9�F��<�C`�q���W��f�����p��#����J?t%[�!�~��j�V��H{�A�ih��m�`ʐ�/#�E�Q���{���E8���K�a1���[�X����2S�SOcv���t-3�k��/4���j�F&�8���ɸ��d����5Q9�rCeV0/¡F�z�Y�,��ʹ��IĦ�7��ҙs�CL��ZcGz��xK4y�:�!����K�!zf��I82��g��v] �nS&Պ ��?��������`�И�`.��t�Y��;5eϞ89�y�<���|o�y�#��J�g��l S!$u�٣�D6�@�ھ12n>����ߕ\�u��&>2��"�����MU��$�:����'���_����j�
d���D`Ň�op�[BpsCXG}~wd��3mHX���?F����$���'�$qc�10�u;�-��iD���fM6j�ާ"�и��^�d��������������sx�5�e���Ш[|MZ��XG��7����<s�MI>�8���_�������^cݙ�Kԏ:����=�����bN��d�D0r]�z };��վ����&W�A,��~������	HL�"�#%����5��,A��/Tl�x�A��i/��j�V�mQCtK�tδ��!����q�U&��J�k&�v=F�)<�;Y��o�<?����Y|�:����C�`ڳH�"h��g3n�v
��f%����YQ+��N�~`[U��>��m��E�W+w�]"ý���fHP��q ���}�~݌����8���^�\����V��U��& aR`�,I�>n�>��G֟�O� #���>��m3�R�m'Ū�,`X/{ �8��J�0ـc$�}}�E�+�[E&	�z�8T` 1Zrm2���<����LǾ��-1�*syɉq���<	�#�b(�xAO��q�*Q�<�h�Q�M��T@E�2~=��D�T!YfGoܻo0���*�p��۵|�供C�ۧh!_ ����&���+��(�7�D�6�Ƚ�:a�g�^�?/f_�X���Hk�$�`�����T�j�1��;���ɒ�k�&��l��4�-���G�����o`}=�����µ�I뎣:�ֶ�p�8�t�TP����-�X~�<&�#�HQ��YUB�	n��ؑ�}��%&�/�;YZ��`ߚ��?	Æ@�R��f�/E���">�"D��A���Jx��|��3�n��є�ՂV�����?x%j�[���(8�S�܈sK�ก�C?ۛ)�2�}�gɵ��c��⠇�ٷ֍���Mv�ڲ�9����Y`˘��쬆��!Â�S�~ ;^�1�M�zj�z�Po��zF+x�}�׭�`;�(�h���z�;�=k�A��u]E>��� �(`��Y�w$�z��7 ��I׼�|h-a�C�H��0ѓ(N���oʾ�43�=Xgl��^������h��f� =��k�Mp9�;���N�#{N��3�6nA%�eL�?AL$nz;�S]��#ωxeJ�	ꦄj�R�����Y3=ѿQi��y�%O{X��� O]zb��?�؝���:��b��6;��91��dL��,ʋUUʣ� ��zOD%^fn�@�t����kAM=�+}A�)#��μ	"	3͒�&)���B��+�� mn�Bemv���y�2u��s�6m�·P�{N.�W�#`@�@���V�1&�S��bV���qpop@����o
dU��E5�&P�vX�S��������&��L�0��2�wl>�"ǎ���uu�	�Lat|�A����a���k�����<��1��0�k�� 5oŜ1�<Q�:���X:6��Iy��h2��]�H��]7y�EDÀ��+�������:M���jM�B�z���A�����:��2�>O7#C��R������N��4@�+�����R��TÒ���>�4e�y�w���=@6��)}ˊ��Q�!W��A,��;�����$�_���-gU2�.w>�	.�D�&�$`H؅� 0�5��8-8u}��P(���;�:���<�Tr���e� 2�ل��m�į��7q�K��s��>hdy�l���0��B!�Nb���O�G���2w#8����l�yTr��D�u��Q9�WX��I��D-� p�$'ʈ�s���u���������kw�h��t[�$[qg����	]��|0����[r�te� ;o�<T�G�+,��!Y��7��ձY���I`�����h�m���Ϭ���V_�>F'�ҁ_oGV+�dcZ��gIy�����Ln^����Cr���ɑ�V!,)V|7+�Qw��X@q՛�)���k&�kΕ<�g�֩�2�/R�cg�Z$4�a$V[������׹�d�kQ=��������ۙ��0�<�5�I9W�wi2�)O].�v=��؟�yn{���W~�B� S�<B��~�鰯C��6^<�`������/���Gr�`�g4$��S��rV� �Xv[��.�,S��"��P&ĝ��
"���9#�do�~�laĖ�����6���pO<#�VN���oI=F<ky?�� �k�Y�\b[��;{�< �	�>��LCn5@�w��O��

�� ���f��cBa�;��(l���u��ڸ]��^���Xv�pH�я#>0��H'�RWNvw�� 3ak[�T9H�U�ip�/.肖b�_�ޮ��?�v�G?ڦ�{[�TnG��x����֐3d�����c��MW7�l�$��(��-��f�!n��˟��̭���.�d��i�v��Y��$Q!�Y���0ت{�Y�:Q�E�߇.�xUV��@S�k��w�����O)���U��FM��x\SjpxA(Ii(j$S��h�*��.t��z.�@�U8�0g:��+ԣj���#�6q.���.�K����nQJTK���M�����ā���'|���Y&IP�>��Q������quޗ���>U���!��#�^�����(5�v���%�ϲD0t�y��tN�W+��䛇�U��Fq�Ĉ
�a'"ZrS��i���)��z����Z��5_�EQ�/?�Ҍ	�����ڑ��������r7N���#��*r���;v ��9�u|b����34� @E���� �WN_Z�Kqc�S�<���wm��m�X���yG�HN��2i��,���V4P�R.�����������S����w��2n�\pO�m������ ��,�C�VL�|��G�D1'G.�3q�g�B��ukՕ	�����mF
�3�z��ü*T�fe�f��Du�VSv'�3�(̀�
NO�W�M' Ay�|P0�.�������Dc�npI16�e���18
��T-Gr�T�?S=YE��}\�U�,���4�J�����,�1���v�P�60L���.�]2l���:�QBS�X����L�}+/��Caȝ5	��X�h������v������7N���Z��������iR�
k�w`3ZJ	\��R�%1PQ�ډn_� 	�S��W�=��f1��9O��x�X���+9���t�ׅ�I�qRl�XMhw�' a
���R<b����?6z-�m��'����[��v��	'�<T�x|{�D5!k�J�No/Ud��}u�M�y��Y��t!�z��J~��Z0�
RY�H�V�#`�Ѥ"M7�<����PI���9���a��=}L�fl�S�����GL���߳�H�*N{��Ю�o2����L�����T]�߫�A~x�P6,h9���fP�dê���].�3��}�A�6,ՠvB2rJvEӆ��6�bw?k�h�I�eXf���~��!O^:���iz�,|�%�>�hG8XC��0����� �ls��ͥh3�w�L}lՆz&��/��Gӿ�-���_�	�