��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��)�-�қPc��dڂ���6CƯk��͛���-V�q����ـ�����_��.���̋$R�dSIM�5Ǡ���1��XQ�.wh|��ʦ4�qS�ք7O��(�(��6��7et[��A�`+ug.��ڪ 0d��wN"��cZ3����@�r^;4�>� ���۲͙���II�������P�
�s`XO>!!�R:�Ť%s��B,���E�(�"��q\�t�<nvD?ldG�N�]���Y@�Jn�(��Xq�������e��}����`q_��zV���=H�IG'?����7��z��*�mm`�}�LTM�F��_�\k[��iW� :��y��]Rف��fA�#�Y������N�G�%��T&��JmIg\�v�i�ҐLAR���I� ���!L��~��n���.���iuz�����y���Q`�9��67�|��c�Ŗ�7�ge;)�����=�j+�+������	�&D�:d��Eʔ�O����,�j�G��8hS��D"o���m��#�xx��	-fXf�`� }(��{����Y�gS˕�B�%��*M������W�� N���|B�G�^ݦz�Y9t�)�OJ�r�|��\��M��y8%ė�6���-��# �;7���u"	LS��9ڠ+�R�����4oi�%H=o/���`��0��彫)@�ي47\C�]>�@�B��FDJ�qT�'߽j�ghx�h��$��A�y5J"�·�Y߷V��V�t}10����
�M�ҳ)�"�|^�bVY��<�����1�O��c,?V��.�]|�5R�!�لZ��e���f�X���-M�[��W��,��������*Do�T��0�4s]l=���T�YRk^��	�L��VVÉ
VZ��ЋZi8[h������{�O�}х���HΟaU����@�����8���1g��q���t��`K�v�]�� Ŕ��jJD(�0�!�ʧ���<��e�..#��%ђ����	r��j�x�����B�3��xI��_
���h�HC�2F�&@�7�����I�v��
��8��mL��e:���>{�����l��7���=S��.�^� wj��k�-\�?�u���Z�.����� �Ӽ���6��[���~52����F(47z�|��,�rs�X[-N�f�_�_��]{��B�ZK�rQpt�櫅p�r�l�ܟ����|,�W��'�1�ʣ����������0l:��HTQ���������+OD���h�����[�!+f}��#�К/���ʞT����8�T��'��k�D�D����ȐXK�c�Q{�giT�f:��K��Ñ������� 1�LIr��k�7ћ��u�P��L�!��>Ӕ�+ؕI����(Ԥ^�/�����	��n�4�n��'k��\��v?����M!�vQ�9�Å�#5?w#�|�"tqw�4����J�������5y����
]����(���;'���	�1֐�;���	�Oe��F���6t�k����$������J{��:�A&�m�3��;p��K~�M~Xև��#��0r��cU ������.�+�/�"�o�'�P�<�I}���������}���G��
�9�D^KN�q):!j1���oq萟GS��[r�o�x��۴	�0����K��ݷ�E�)P�,Q��׾������aiN�<
�r���K���C�Oq?�`���S�'5�)��篸!�0�/7��Q���I2��\��(@��$��Hҳ1{>�/�뿲����蛨	h�2�$
Զ6�3�������c��W཰���}V"W��EL-��4)�@��mKU��NRf�6_�u��L���'G��I�i�t�I1٫<��Of����w�u��ԏ`���Ki���װI���y{Lه����jb3�m���Sź]��)��L�U*��S����݋�����ͤ� ��4�D�:�$��c�0��ض��P��Ofd��\D[�0@H�-�&t�H�����3��d����s���C����q�0��<��.0)�.@���|���x�u�Ge����}K�#uƟ�ۡ�O� }�LK�Un�Ś��)M��}��{=9�?L����NXY�$Oyh��"�>����!��LU��,�����[���ԃ���AB�:;jTwͥX	ٹZp$A�9�y��op3]y�����W���A���+;�f+�c��*n �lA/%!	��O6x`,��3�u��ٸ����-�kC$���_�r[=^���G�>xDV�{��+a�b�4)��Ж�7{0�����ڜ=�0�F�8�a�������|�����x ���]쑓�Y������Z.ʸ&g\j���{۹:��L�+��#��0��F���t*�'O%ŰZdα�B/��ǋ�(�0Q@�H���/oW��9���� M��v���/{l����>���W"�}�?�N���c��-zUr	-�^H7N��c���0P�o�~sl�~#�.�'��Z�U��o�2죴	f�>M%�Pa��D�i�g��Sp��q�Y0����e���h�A�H�I6�Sg����\;m�\��i1�7��Vu$�l�����P�EӔ��It���7Ha(j�"m���Ւ�s��EjlB���+�����i?�f�D%͘�Rt��K��h�W���?x�hR�x��G�8]`C�[��x�&Ҍ��hT����O%����{n�c񼹠�*���5NC�iz���U�Nhr|ԓ<��9��	��hVL�w9k��*�p�J��#�d�M"�� ��!��e$�2�����p���DV�MQ?��;��Jt�=b�7O/�₻q�]���"]BY��.���jUŜm��M[аDI�#�.�VBs@^�ͻ�'��[���"�O ,�A=:/C�j5�
K�u!נ�(Y�[���1F�3�]p����X�S�=Kݿ@������'���L&���x�'�|�d,�+��B��li��1e�(�N'3��s����Z�co�w�����{O�lx*���ݹ�.v�L|������~KJ��|_9=O�����F��#�nM_���P� �Y37�u餘��0���e�:eh�z���7����}��%�|d�7E�"�O�G�#j�������mcl_�/3��;HH��SE�εdZ����!�k�Ƚ�|'��N�%���Pc����k���/�k���L��XI�i��X3g
�9&�T�R�g�YV���h�Xb)���B���),J�Y��3D�c���U���_��lg�έyؚ�Ҭro�����Mw����vO!P-��1��M�f��Y�Y��پ�eL�6�<S�D��	0sBrvt3{���KF�� ���y�{�X���k���;��S�7-�S���l���l�ܲ��Um{���$j*\��&��d��N�qK��?W�Y�D�j��
��Ū���qt������o�����,�w�>��m�,�-x&�薴�S�,�� ^�z�/��jmAB��,�қw\3M���(.�R]�"]��L�I`���t�1�� ^�ǉAv�{2%�/<�[��I���8�g[H���C�D�ȉ��z��>fY�Ǔ�}2��gU���Y@�^y/#鞫�F~�%�rF ��V�)����e�J�X�a~��{��@�iV�2ZV�s��j?sH�;�0E�[r�R._T��=[W�� ��*I&;j@��t!��@��f��)W�1��jY�����/��l�=�����tK���<�g�b�����?j�� ��ഫw;j���L�S��
�1�˱'R�՞T�f|�+Q��#��[c�n1�wt�j�5�h���!\ �{��:�M�o�WD�m�m�8���@@q�'rO���p�گ�UQl�ʣ9�?.!�1X�s����\i�*k.f�+.s�0c�����h�c��_�^�8~����vpF����]}���xh:� ���,�ȃ�Q�"P�zj�<2W(gñ.SH�HDz�Ƭ��L�X�U`�u��UŶ�(��t�O��g҈٨�]�n
N�
�"���|��B\����bn@��և=�ӆ-��s�����"�����رh��Cw���mI�7P�hE�U�b�٩��N[�æ��%��M�[��.�*��%]��pR�ť�ȄZ����b��,��ع<����2/uH��=��s�O\�;�A�� 	&�5�vd���p	q"���FJ������hYv�y�)fC��1���~ɣ����YH����9��VKG9��KB�����`^���܃�w�Q6��<X|Ǣ�	�8�:$�5�8��caaogg&�b�[8�b@,�4�.~DA���?�
��	���J�3���~�;�$K�N�1�*�7=���c�����K9<=���n��9`&rJ�A�,��ھ���R�}�xp`.��\�A(���e�#ɀ�Ǭ'�e���r��F]Hv�;.�=jn<5D��>s����c��A��_߼� ��*�YP܍%:��)@#��@�A�:x=�;��h
J�R������?�~�ڭo-����������WY��z�����(�/�3�w��v��[ёWڞ�٢��|&�9�R?R����x{�
���H�����\�g�(M����C}�zl�?G�j�?AE��r?A�j,�B���+�Py���f��c�ڏ�Pug�NMr!P�����t���ބ��P \2Rp��d�w3��UT���06�6�<�}���gO/@�a.y¢eg�b5_��r��;��e_f1��	C�����Y��.�����������&��JW�`V��%/_���H�
r
��Ab�ŏfe�M��3Q
�Ƈ\`&w'J�Å�&�ڝ�xNy&���,�Sڦ�Ͼ>˼S�w\+Zl�dk}�%}���F�u�t��d����=)�?ܾ]V����������z���00�z���s	��R��uM�4�'���`B�m��O)SX�)�;����~)��Ǎ!f,�b$�^ª���܃U ����e!�Á�-��~bk�w��$�Y�H�
cC@`%��s�J�3ɆD���}2�����z1�NSR�#���F��_Մ����s�"�ɧ��F�@�ƻb-x��2e�~S���r��/��:�mY�j��B/9
U�B�����tOQ�6Џ!A�Lk�=�-�����:�?���eם?ׁ���ڪUL��L�(B�=ͳ�i�������{DH�R�ò����
�ċ//���q�P��]���1��T&Zr�̈́E��pL���IL�G[�N)�2�i�T �TĀ��F<:��zL�����V���k���zPB�$���d��v�����H
m%(�ٴNU�8��.�Nh8����������O��3�M��6��a�!�7k{�:A1��;�����@� ���J���K'ۢ��I����L��>Y�ʺ��g3�h� t�+4�2��+�b��
ZY�VL������N2O�8G��f����fq�X��9?�O�Q���^r��uqi5�������D"02K����y*(����T�I�3�C�[P�֊�9���G V�Wv�K]���-��ó�ZD0�����R>���#9wu:����SlRr5���:,�k�!���XX�.S!�ـ�
6�=��:���k�(���]�p@�l��
�4���t�45jhZ��6-F9,��r�������²�o!��Q$����Y�s-[���;4�ʓ'�l��.nwaP/E��_n&��!��|Q_=мlw	v�p�����4p��?dg,��w�vZ��d�b5����v�V;�<}S�v=��u�n1-�N\5���V.�>8�EF$N��}8��Vɔ���#%+\6s{�f�/:�'�9�vb"�bx��A�`礩��}DDݞ�%dפ����������*Q�v'[Hi�p}���;/h�����1����[m$���Sw�O�%0dt�xm����k�6��\��j�JAs�%�,��ʮ��[;9���tY�]�3V��N��h�c�!�w����^�Z����a�d�+<�
�F���]mƖcl@qX/�A靋�ݶ��й0��3@�W*w2���)�a��%�B>�@�Լ�9���]A|۬�����b�M\ɕ��ďmmc9dX���%�i^CN�4bg�,s������ە�[���}��y��JU �>�^�5?;�'9[/d���ɜ�n��S�ǁ���?�E��e�4�-�h�����d�(��_Y3�RJܔt��uB�����۟�FtcP��t��|���2����疨eYƦh]�4|�P&W�
��h��uq�D��k3����G#�Vtv�|¤넘o���9fjɻ˶�/Sx}�U:?٫�'����׬���33�mێ�,��0��L��{1�]찧q;����%u��Dr�'�c�y��=A���p;.r�{\F/��u����N�����>4�*�4�#,��>����:�d�"p[˙�ɗ���X����0
4C�&A$@[E��S�q���$ߊ�F�]=�j�j�U�����_e���1�e�z�q�ᬜҔZ��W�L$�r9|/�����
��p;X@U!9��U/T��W�������?B�`m������O�UT�*@8(#4�ǒ9��������l�"!L�S�K`@�?�'ْ
�",m� �j�L�����W4��  �ED@=�I��[��f���z�`&�&��_�E����>�O�p����-�[�1����b��A	)X�O����X;~[͈��]p/�ק}*��)i���QL��4E��v��_�G����J.=�ж�N���լ�ǥ��
�WAM@�W6�bش|2i�9Nb(s7�:�j|Kldv�<����^��#���̭*�W��CNK�g������±-5�%��_d���P���v�iI��
;�4������	ȡ��24�HV�b��{�[^%*#&�_�)�s��(�^�C|�8Qw�A��>�Y��uɍF<��	y��ζ���(=,� ,G/�|�|
x���%��>c�]MR��Qĕ:y�͎ X�D`T}��tb�
�Y�����؍4���3��*�?���U��,IS�F����i4�Y�9�_��=��
��^����|	�1���X	 ��ٖ1�<8sQ�D����en0�ղڕz�m���!��`��a�[:�yZ�%A��p�|��r�D����4�c�vd�s��K���B������9�rj�X��e����[,f��Gs�b��YJM�P1��	�yd�U>�U<ߛ<{m;-��^�L��H&�B�ھ�.�<g��㠟T�_`��&C��}��R!�~�$pik��<x���;�ǖ�C�H�ո;�'��Oz�/���~�5ʶDP�?Ez��n�xܴD�����I�7�]�s� � ��vpk�`d�"�F}&�^Ƶ��vW��/�^�cɃ�7������o��	3��Cx��1�����?6�3@D�H���j<�=��Q����O)�(�ݦ\D� ��O �I}M��,qV���+���������nK�(�
����p���X+�7��q��FP��b�7��Ey}Q1//��e\��bV;�Κ�K�x���v�O�: ]s�li����߀�8��R�.?
d�4�l��B�.>���ώ윘���(�7��_�3����	V��tq���G�c�&K�U:	�D�2[����Π�kM�:k������d@��xKC�&�Y��F�X7�ƺ� 2��]`x���I%^��SYq -��]da�x�v1�4-�dI@C���i��9�<Zh�vwl��Wh��C)h�z�z�l����Lz~{����-�Q�Q�i��:<�X�DQH�	�scPv��:�w{�"��+y!��3�u?vđ2�&��e����c��4��tU��]��&�ë��Ǖ��7a�l/$X��'��)_Q:^�BK}n�"���)w{��F�孬kBq�jiw6d���3��E��\���e��_	D�O���9
H�*CQMsyd�G2��jr��&D�������U��Ig��=N��Za�n�������ڡE���7�<�s"W�A�d�AM�ǔֲ[�t��������a&�8f5�#��c��7�1c��,�s�(��"�m��wV��v�U3���%I�HM�٨��J�°��r��A�Tʮ��#:g!�Q��V [4mwi����r��s��e&���D�JV�?��C�ڨ�\~��~��S"�H,��L�cޘf�Y���8HEf+�ϋ��aJ4�
7��K�� �tX%�6�Q[ڲ���m����'	?�3:�1��]Nn��uΨ8a**[�x[:���b�"`����aN��5zr�Y=�T�m�6�&��7�0'�߆S���0ҙ����|2^(�1o�p�������z����2���@+��g_Z�}�XS���l��w:��T��P��˻�n1���|�\jd�._�V�`1Տ	rk�,�6��_NQ�D�O��c�y��:{�y��`��Yt[�-lxc/q̫�]εL��r����IGu��ڟ���f�r-]�����KZ�sϝz��o'�U'2�Zi�����D�zj4�NF��r4B�̜wU��_�T$��ĈZ�+
�����BUݾ&�B>9@����gȨ���:(:%�����&�x+�l�w����ŇP�O�5\&~*����e���� f�����bT�7���W^ø��NwG�zD��1��ť@�m�ƣ~���C����Q���oУӌ:E�Mz�����/��ɺD@N�p������� �N�F���({�Ai�*M*�>PY��U$����Ɵ�aɷ�&��A��4�kt���Ơ9FeG[������&`�CUX�f�I��T�D��ѩƆt�8,Xf��Q�HY�'y�Wn�xM����M��%Έ�8�ס$���✟���&ґ�nd�s|�s:NS��J��Ͳ��O�b�[�W��z�.���e����'o�/��uQ9���m�I]����%v�(�ux��')=qG���O�4��6��Ͼ�"}j'D��<�?�ۜ�Ūi������<�ĺG7
r��q�<Ți��.e��V�E��*z(�Qʨ>#��/�;<V՟{s�'MIwI+4��Ƈ��R��U]�!�,�O�/`����鱯c�!pi��S��[p���S������.]AT$���
iX,IG�٥{�{�7 ����s�!<[�	�MP�a�UkDS������X蕍����B�CY��б�+�rv=#v��~��#�5�~@O�n@܉�X��	��v���i�CI�ѾӘl`v�q&fӵ�E�>Lo�7	���S��S8Б�^�duԊ��ff�;�Rh�	XThb")�e�G
���
7�ā~F
sp�l8�T2��z�ºAk�������0q1%��6O��N�}�-S;3}��|��C����Qڻdy/�֥���-���4�����͵�k7�4C�~[���4%9����a��y�or��=d4%o`�m���gG3��ս�D��>0��?x���bw�mi�A�t��m�ہ��3B����A&9x>:6ֱsi7���DNW�t�yA�3��6}C^�1%M�7��6�8��JSk��l<g�\S`���@�=�و����	-l`��k�`�H��'��+ݔK��G�f0����x!7����ٟ�E*��y{i�q����q(��#,���
���r���;�I���zv��!SVͨ�f��,g]����p$��koy�,�z������)ưz8��R"q<!C�� �}��8�㿛�Q���3,W�,�d.�Ъ_9��;I`6B�_P�2T_ɫ����DSp��"�h�!o��$b