��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�E3�hoA�zFҿT�e!յeK!�����59��\<1z��G����HS������n�z�*exd,�D弚�ф��bJ�l{�Mm@�w��Yd���1��N!q�"���&�<C��Ċ�ˢ'�z���(�\���5��	Q2�I iƑ�sN�Z/�f,v�˭K������� ���R\�@��G������E��H���MY�!��/϶jV%i�����I;{�]q�I�_lk�^dԆe���^��S�1k���*�>�jK�HLg�l����fk�{"����H�!��0"�j�@q	�!�&%!�$:fi}�4|��F:�t� >�q�_*����U���:Fv/o?f�p�T$Cɮj0�Ȁ�0�l� �v��Ta���xόE��q�_�|r��g�;�IVh 9i��j��3r�DˉU/R��"2h&��Sl]��"XaU�����׀P�΂կ�OsHK�i"+�*_E/+Q(��/b���Nz�Ǧ�X��S�ƞ��]w1$'*Ƃ]�_�%6k��jj��H`��.�@�m�}�nb�wlh��ϕs�)�u�lzZ�#�ͳ��B�3:>Μ�<�R2���*o��d��� VU��~���� ���wm�1��Ml��	q��:�v�3 -����ĵn�LB_p�|Z�XX�o��ғy��s�(�d�SeGmaCE6)���N)K��],ǆ�[�~5��J*��1mk<C5�a�����$�}�/��{F��x�L�cT`��~��M��#�${�#¼w�/1듅}����~:����/�e-�Oח��!�XO������/��a�jH�R��߮�]s�0�R��pU+�ǣ�-�Д𦟛���|����253-p*:?azc
�l&f|����܆3&�݂������)X�S�؁�,�2t������o�
�,���(C[$�ؠ$d�|�F�s<�ʏ���w�b�qưߠ}_Kt�KVCJ��P�뫊3�F]��^�'��7�{E�(1K�eGTY�Ȱ���Q��w:��QV�5~�k?*�5���ᗠN�
H��8���NH�SV�M;�|���d�YD��}t�1&=z}j�L����b�3(�ƫ�	Icm��=�2�|g�6AFԟ�%�O��#]�7��`6�J��P]f*K�ޯWo��TM�;KIs��G�`�o�c׆v�9Rcp,�KP��S\����Ql����K�U2CЭYx*�P�}�����5Z3���G�2���&bh^'Լ٧V%�P!)F���]J���1,��*�nm�>���%a��[��t���NSAT��\�ߐL�b>�]����OBꖻ������{����ez*[�m��f�0u� ���,��b,��Y^a�O�g����y넿�/�탼�%�!�����3�o�xѾ湋�S���E7_�"�hni�uf5�%7����E�̙9��f톇�#O&�)8ծsMW�<�E!&Ϊ�Š�D��{˱ݚJ��u�|�����31
C�:�r������6��d��;y�{Ϭݏ��,�u����S$�����M�M��ќ�� ��D�P�}Ő�t�q��7��|�<��0)`��؜�YǺ���eZ7��b��s��,�T �\V;iT2��ē)��1���|��f��_ ��QY#�Wo�^+�څvt5��c���f�0�~dM<��s��Տ�-?�-�Z�0�b:])J1Q��C�t�BǦ�{P�(J�����)���[  �:!?�e�C��ZI�A�'�����X&�M�[�����UGO��5��z�{�|J�G��_�&�y(H�^Ƈ&�f�&���	�	����@5.D�Ï�#v�K19i���2����bi�hJH���%��q�����4�Rp�k)�f(WED�ޭ���SHn%| ��o(^ �:�bIi;͕v�7$�q�)x�/.��4Uꬸ�N��M�z��c�L$G���r����-�`��Qop� ������v�@��N��}���N ��p�oذ?f�#;��O�1�'3y�s�XrbG��|�!f�]h����UN�c\ P�WN��*�#����?Ŕ<�$��sd�ݖ���5)��Ѩ(ʋr��\���7���Bd�\';��ͻn�0�o��ۯ�s	�X����ϟe9�
���Q8��iX�;��l�x�
*�:jb��ͻt!4T�vXd��k��U���%ؤH��v(���s��8)k����ʭ
�����wY7��͖g|�O�{)���n�[�-�k5fm^��a�Q�"%KX(n����G�1��t�]����?S����l���^H�+�,=�GΫȞ3���du�!;�Na���n�X��o_\\��4��D�&���.���@���_�A�,�-�v�#�5zP��L�Y��3����y�-�V�a�V~�\әp""pf
\K<G�n�;�#�Ź� v6vpbm�ܫN
��.�h��E��,���l&��[/����$#K��{᱄@ʒʂ#I��=9K���z|���8�����̹2`Q#��z��I&���g���Hw8G�~��Pe�!N���_���X�x�� �����O5)���@�R6>m�|Bc�s�e20���'t4�D,����1$��\��~�YN,(��msf��S~q�~��u����5���O{_�����'�G�W�;.#�J�+��ɒJM��˕�"߻�ڔe�c(C���*U����\г���X����
lg�y[�%#p ���û�X������Q�ofW��6��<�u�,�^�[�QB�еUު��=���N��OT4�غ(��3Ny��_�$NA�@<P��ɦ��PA�F���ŀ����Q�@K�f��9����~�F�.s�����ޒ=����K���"?_K��� #=+���޵��beU,,�8�Z��s1!���㇍�Z,���1h�垍OP&���i>�7\���ǀ������"%��f�%�x
�g��Z�,pM�ոygsH�r!']٥O3��-��i�ص����0�"�<Ҽ��\Z�M;��8k�Pǉ�w'xb�_�ΔVZH��}�0�S�I����Nn��|_u..m. ��w�K5��'���Z��{�7��y�M�7��7'��nu�޷OYH,?P�	?1L��]�>ۀ�Z�^�6%�_��'Ի�i3q�W�@M�8lE�d��%S��
��y���=���4_��>vudL0qŕ�{SB�*O�x�>�^2���D��:����9Z+#�[���>ar�1��Fjߴ���L0C�
��,��T�m�*�	l2�c��_@�+	�B1_"�!Ț���uo�gW��|@>)��x�hso�rwr���Q�lG3Ę��4�R�0���?�;�LR�Ն�#\PU�����x��j�͠�ތ�>3���%�5,�Kt����kj�D��H
�L�Ws�T��ֆ���^+6w�Y��l�]�o[��"��҈]���s'���"���ֽ�A�b�X��ke^������t!�SU+�����+�1����[����~3�������R��cz������G�o%�M�d;d��=:6��a��PQw��8�'G���ӱAT~#�+S"+��b�-�j�Q���(�a��E���q6��MIzG��ȇCg��H���X���9���=�`ƒ�)����܊��׋x?����c�BD�:��1D_y}�cRR��3�Cݫ�ԡ��q�
��46��,1}4R=��5r�����������B����
K8R���Ҟ��N$�K)3J;��t@`�-V&k	U���HAA��R��8ؤ����SEDW�U����nq4��!�Š���>�u�t�ϖa50$�Nr>U��tMv!�=�In��u8.p��4y���U�v�Ӏ�bߝ{�Z	����ҾD,�#K��SNO�Jw�9�UbHalƾ��=H��u�)ϢCL�BMSi
���$ϫ�;����s������Hdkv��kXE��f�;i�$�@Q�*�k�b���]�zJ�;"	�˷�+����?�F���a2�y��sM��S�2�O_��&)��Zg��;m�� �w��
��O�����޻Ѫ\�#������1�G�\����c����;y�l�����U����&��_b)����7v��#Z��]ϝ��߳
�2�3�l��J�z�ֵN�'5^�O�?�RГH#��Q�H�z�����~��F���=��?�CZ��/Վ�-H�Y�)�@��)P�m�躙��9�a�}Pɱ?hѺ�9��`>_��9�.�Lqay�Qa>䉧C:]?��v�u"v�'Gb5�Zjۙ��n;p�}����`�5ǣ���e�g0Z��|�y��'0�S��hL�o}�CCV{o�؁�Z�=��g���<,Ҥw��1jV�|���,^�*H�����&�IA�4�W��(4��s���S�O���5h歾��q��菏�-B��Ґ����:v�ˇ����[n�JZ�U��4��C���5$[�В4?{$+1�OxZ�p�P�9��=.�n �>?�a��$���!�S��J��~��/�ۙQ�r���<3�VZ�r�"��@�#&��������k8i�5y!��eed�M�Ȗ�٬�?�.k3���K�}��q��/�K� �g�M�ӥ�%CJ&^��*z�8�c���(|���ŧ{�Q73��:�~��Z�G����Cn����PG��Ԇ��0cڿb�[��ι���#)2�3ç��Ǐ"=��)��O��y
��S���P�2�:$��!GQ���Mg�ҺdBA1{,�њ�M�,���`}dv.h�5k�u�ƙ��J��s6����?�Ⱥ��=�d�3�=�\�6� ��B��� nm� �av����R�0؏(+�B�Y;j_��X������y�v�T������^3�5H^�����/O�\��)�0-9� �����>C[_�^�Ix8�������6�̝@_H��m�<�Z���R�l��]��d
�y��b��c��v��B�����~%=-<��,4T���Q\�]�f��|9��p�րC�U�K�(a�sI��qqڌ~9'Dn��K6�Wwq��:�b��JC;���2k��xp c�C��/L����?t���E���� ��Q_���&�������@g_��ұ{�aC�֫�f1�ٜ�X���a���q�<K�]I��$��}��zf�	/�0�kq�޾���K�h6�*�R�of�{������*�tN_q���RU�F�S�w��!�n��>�4�}3�׫&\
�ҏ��DKBx}�r�����ڰ~��8�Ji�{����cP��Y��kr�R��?%�\��:��!�/��һ14���/|��'�/x:쳉��u�{�n�� bp�iwkl;���M1������v�e@�P��@�fX��O��eP�F���n��<��M�ɓt]�[�8�P�B7����89