��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�÷!�J�T 5�h��dp5�oU�)Y5���8_�y/"ɭ��6X�xYY����F.�[a�1.'}��[ ��.��h|�:_]��ό�m���>|��c�|�3��_a<1�Pn�~z�3/�5_�$	�o�*=�>�nd3��"V�d�/�24<!S��r���'k_q�x�R8�^;�"�_��O;�*�3�p�W��y�o�0�y����0R���}L�͉G0;Bwdt�r�k��S�ټ*�+s�q?�~R�!l�%�4ƒ{����7�e�K���ڪ�x녤2�%&Q�Q��B�q���X/�D̴�v���,P �/���,�Q�y4�. �����XDǘ2Фo����ΧX@D�����&����S��];�e[��T0P�֬�'͠���!���J��2g�l`i�',�^�r������x�Ed��x��,��jM�Ͽ�� �$��K2$m�7��p7�N1<S���f{��|4�1���n�����T�I�����~���&1���L�6�9K+�ֽZ�±SBL�i�)�����3� �DK
8�����A=�|�!Y+���ѩf�?�}����ͬ�D{[��(�6<�V���ٸ��c��`��
�o}Pg��_���?!��^��S
ӣ>�6'dj37/M�A�$]+�
�!����s4�y�������S��5��m�;W�wa%�q�� Α����?i�@h�� P6aq�3���y�2"�B:��=K��Is�br*�Q�9����$,�(c�4�ɱ�6U��C;=�q�ɐ�g��	����5$�L'���� �7�g~��J�pp;3^}�4_-k��}�^�4Eݡ5�����r�Ｘ/��g�Ì�h����ۯ��1�����S��4ز@�!��	9��
��S���$�PZ�B�K"!��8�Y��lG-B�C�Ό��ȕG:^p��.<��F-�]^[*�=b�����܍�u��M����'i���'IT����i�3s����cP��:\�[ct�+�h�k�X�c��\��v,ҍX����7KxUC�1 ���VB�ٱ���5���V�#�K��1�`#&���b/�7ŏ�֓�@��"��R�)yn��݁އ�/�th�[�ԮPMnFv9����Gh�i�^̿�� �J���#����HK�L��]�F��c��$GѰ+�`j�<���v;M������n���Jbw���S��WJz؝n�l���vG���
�k�s{����|�Ҕ�X�1�
E�h��蒃Ūy¨.�}�ެ�� �	�h�aFFg�����I��{�����-@�I ш\/�c��̴����H�O*($x_h�k�[�"ti��Dͅ@�������G>6ٰ*T��8A�|�գ�nҎ�wN0�Xԛ�:���>�`��-њq;�k�u�{lzLK���UX�:��a�pP�p�53x(#qs"S~�����&d�Ā���dNď:�'�񰨻^��]�)r�]�#���K�@^vu�@=0xިc�8�~�w͕.ȹ"�~��b���0���4��8�|\LS_�>pK��Q��Y��d^����/�T��YnD�}�%TB͉�!$����	c�A��y��r��̞�����2�T�"����Jm�JS*L�|���3�'�b/�e��>��-�Շ��k�e�;�)F�{���}�o�ą����J��c*s֠��ջ=2"�9uT�T!�RK��ĽwL_F��6%6��Zڜ
9��#�AD�05�v�,iwOc�c��C5��]>���8Q�gh�Aq�ҮgƙIk���;<�f�շ�%<�<��,�LY4^�S��oW˖8����'*�la r�A��_E6��oC���^������<��h�5Ҭ\��W\�:L{���&0L�~l��).Rߜ�z�p��"�������(ZFq��fyn�r�3��w~�p)r����w����Մ�^��B��&����xmB���?���*a���B8g���W�	�ꕹ�m�>��S7�0�jo	.��S�G�g���mQ�iw��ɸ��{����\��LdQ�tx�c#d���pC��1g�;8����٬ ΂P�	/�R��5����u\?k�M�m�<1$����	K�`u >�/��}�P��B��Ǩ��1���2��3~�5�ap�ǍJG�TQ�j�����a˯Z���9�%M9����U�
�%m-������(E�&��Ua��Z_H&o=��
�1=2���0�G��GI:�[�9~!�}/���lz�%Π�U���49��r ��Cv���X\.kY�h<�Y(���?�GgL~7kE'B�H�XT�P��4�;g���#�I�� �C&�s�V4�+��mQaj���c  l0��>w�����w�&���
Zy�S�lv2���l8Upw(&��B��[&d�Ǣu�>����%d����W(�^�;�OS���A�y�È�p���2EdA����>]��f�K�� ˨FBO֛az�-9�Ph��WR�6�-��{����m��&�ҿ�7R���W��2G�V��
���W�s���]��Yҩ9�.B[�&hű=�~�@�2��L5���DI}��FV���@S �ToN�"���q�5P�46b�D9�O��R˙�Z<���}z7�;Sz�xB��6p��-�H�)ÞL.�E<.�耙�34W0�$k�����ʮO��z�ֱ�n ���5�#¿�����V|�t�R����*r��ev�(��o&L���o�V$rw���К�W'ha O�W�I���D�3XQ��o�ƶUei�I�*D5�ڸFzi���lk�Y���|D=��$�e���K�LGR/k��
�	���?�⎷��=�К��	��\�ym�tl�8���;�V�T觴E���"�3.ib��|��U�����k^a���2��--=�!"7������S�E�M����iI��%
��G�<3��_�$�E�Y솵-+"��{G���R�����ڱ�*��~�[{�}^�£FU%*����ؠ-#لѥW�v��]��V�i�T5e,�3���]O�� G)4��w�F;l0*g{�t?E#6��پ6���]���<v�& C!�� ��W�9��覒��u[�R7A�&�P@��ZZ���=���6V���.� `/�J�>�h�˚=�cA��
\���ב%�#w�F)����j�T�q8[ܡ+�c��=�? l=,G��S�N�fa��Pd�7�u3��b����߿*PI���N\�As%�e��}�r��PUS=�<ٻ�_�k~��B�ڞEgKyg�=l���:a[�H�I���;�q�5S:�N�ڭ8x�/OE6X��^�A�In5�WE�*�k �V2�^�	��1K�g���>"xc�q�N����R��r|L������q��~p�D�Ҽ�G�2��	`������!�@T�l(x�RݴY��Pk�k�� �q��6e`ܭ���5�Q�X�����͸fŨ�;Zܓ#�C�'�eC��v%�����"��v������.\t�,���<h�?I�D�	S��kcM���n�S�l  @��y�A�2E��јs�zD�Y]P._��R����t0&�9�	�`TmY5���gټ�Wc�B;��4�m�I`��	��{|�2��?�C_2"�IE�/v�J�>���3�9�&i���ō�����'�]'a-ǋ�e��B�ּ��^)�N�����tk�.C^#	f��z�#5-ҥC�����ɖt�`�1�P����?��Z�kn�'*��6I�����,�aC�m��wȨ���⏿`��A|sR�m�9rd�;/�&�{I��.;����O�m��(Yʏ��p��gXScnܠ��jxsR7�3d����� �ʳA�� ��5�;w�VZb�f�{+�J��TU��!� +��ɤL7�`V���l:����u$���%���cu+��dg"�EbT���n18����Ƕ��U�{y@�5^�;��2�s;/s�Gݸ^t�3������_�����a��b�yU�v;���j%g�3����E�`j�Z��}�tl��	a��1SR�g9v�?��=��x�rF�}��<S�m���{F%3p�Z[���(K���E���t:đ�l�ҫ6DF�ш�x�d^[v1S�.@'�3 ���֯<�ѽó���\�o�o��� WK8�>!Tg "U(��'��$E�&����f��"N��_���Ȳ�.Hp��e�>���撰�q�G�xq���	kBKR���c�i���VY��kiO�p;�$�70ڳF/�����	I��s(LY�Be�U���C��`#��GN�i��{-�`�iY�i2���HWۇ�6I���)~�� �ga�@�("	��(0o����`h�:�ɀ��j���k��a�X'� Ec�h��<���(}V������+긍��.n�Y�x �c�z��6����>�UT\���kn������
�0�-wo|��e�2�츳0Pϧ�+i5��R��6y�JSS�uے>ӷu�VјkRc�tP�+@�[CG��t	"�K[뜇��ǈR��[!�;_?�-Ml�f\)�
�+f�1j�_��=�H�q����+������%�X���yX�)U�v�I����'��(8����@O���6�#�MqBF4���Q)����_�ߕ�=K$�-�7:d=;�X��ܿ���؀]�5�X���$�tJ�X�*ZvDnc���vImw�LYO���h�j�2+T~*l^E)Lo_���ω���9m@C����D����qmk�wҚ�hLx��{��
���=%Z��ܻ{O.P
t�>�"]�Zs��q�%�;:��O������*|}Jl����l'�]��]��5BMpeÞɞ�����'�M*2����\S��%��}���|f�s{�>���5��,��%/�T��S�B@թw38���x�&-T�T�"��[���[�'w�!.*=��f�T�ۀ�6��"?�_��6{��hCB4��F��a�n��L�2��k�[��C��o���u��ò�O��|���D����������n\xWX~�|i
cp�n�`�Q2��Pq��#:��|�D�QѴ
���������	�F���b��D�Q�(��K�4���жM�hN���W��}(F����(DiX�JX�����E(��xt_�%�hR~����&���#��G����lau�htJ�-��j�$��76G�[t������ŀt���fS��
L�Z�&7Y�/�1D@���ȤI����!�i"������
M�Ŧ�T%�]����t�ZE1��a�g�/���X�u�5O�t�J��B��I�	[�o7��M<�8��zI0N=�j����㾮E�:'�`ʰ!�\՗�oSm[J�QVW��?�0W�k��y�ɏ�Z�f`��/9�:��&ox��}�"~��sx��f�d@�+4[���?T`p[4��4���wL4��D�T�X���PAC�����|�	���6d�뫒�Shq������A���}<زփƾ���Ds��T�PŸt��X�`��e9�v ����!	�|Z��7�<V��L8�.�Ow�p%�*��y����C�jo�lM��D��W��.����@�ksYe��$@�$>�ւh�
o�]z�3ݐ{����fyӋ��Q4�/-!ck�!���j���� �1Y��:��k>IaR�)pq��_�95O;�x9�kx!:kp��7�
�9����"6���j��|����Z�����sOq���/2_4���}��j���g!	X�ބ��3��Ҹ%sVv��@��]�s�U�^�:�~�A��=�M���ȼ�ַdre�ķ���Z��0�uľ���� �h�OTL@������@.p��o�_�d��-HÕ�.���!|.�K�p�����[�����$��v'̄����m(�GM��\X3NP���׵���^z�8#�O��*)N
�~�~�ϙEv*�����_��:-��0t�z�`�SP6U� � �X�㻭P��t`�o�*�So�4�H������s�������Q�t�N�;	Z(h�zcUhSb��S���H��t1Fh�\�����Fh�")a�D;�M��y��S/8l�ȂQ��T*�������:+�XU�j<*j�QZ#^�=n+�6��F����0�<��	�&���(���+a�'�i8�L�~D?J��:Q��F�*d�}����K��zܱ��ſlω��T�	��(�e���9�Q����%:p�mN�jzH��'�
��Qq��o���\���X�[���3~X#�o��T�hY�n�hqO�>yB�� �x��X����qx��W��~�����2ti ��o�bY�Y�X'_������=ug.Uz��e0��J�̄n�{F%�/-?���ǿ`��s�=��� �:�<� x�hPƍ����?t�2�>�.��0
i��e�V�����×�*�M0J�ֈ�槅Q��/�E���M&I��H� �"�
�]߮� ̺dH"�i��kȵ�&�1�{�������(H}`3�4a~ ��z��� 3����ک������dw�S���MU�u�K�
ꦻ'�{�u��>���t�NA�I����?���K�$�{�ң��F��f�2_������).��1`��_���Ho��5�oZ��@�w��i�rU*Ľ�F��<KK?��0Ǐ$��_TB�-��L�u\&b�C۟�@�^���
�Gޑq�M�At��c�r鞻K@nv����6�O����.�u�W� }�(S`���@���Tƕ����7N���]��(�W��ieL�HO���`����b���MQk��eE�ʄ��0���{�UW4��sx%7�60X�uK`�������t&�=�ǩ��j�/�a� '��S��
?VD����?#taUV���˒��n���0�8�R�N�s}�k4"L�N2 ���Q�CWc9N]F�
b�-��Op=���K�N�F.g��=HP�)	�nf�ei�r���teC*ʗx�x��2CQ�c;�����d�ת��P�#�6����A�<Q�͋�����H.�0M����*�#-.8cp�h�@D_�<[>GY�27�r��f�O��!M��Q�G��\�z"0L6�R�c{	���ʉe���З����&�k��k�%��f��s�2�!߮��"4���S4�5|<��#���o%TvØ����\1���{[�I4�l��Wl�^�$��MV��ʦO {����6Y�go�����܇=_h�� �@��t�u2��{E��и��G�W��/3���%_EdX0x��D�I�pm�����.I��s$eT~���ӆD�D�ؽ���x�����
~ݴ,��ԗ$�<���L�US���_=�.��/����	m���u6������Y�I����-\�v�(��nC������������J8Mh�`���{b3��� �EK;�Y<6s�K�������Ex�s�^v �*�	h���E��lp��D�"�&�d"�ji6\AΞ'���H�G��Z�m�Ml�׆0l���2f�qA��K�ur������ ��&vSg�\���� �Ig�4�Cg�Y"��J*޺����p��)H�(,P{r7��]��V	�8/�Q�%�����k ��Y�:M��.M����׹.�]���IU�Xל�35��n!��/��N��1#�`�,��^��BI��'��x^B�s��p����x�K}�����R�W��g�� -N6�|�������r����NE˼;�Y?�-L��ￕzl(�<��1�#����9M��V�A~K1"�jP?I���x���j��%�!�N�h�+���x�	n�#��3e%��F.yJ��ט�2W���6g�{��@���X`G3��T,}c7�������i� k��3�̌�ML�i��yE+���A~S-5\7�;�ܘ�?1�P������Tr��t����x��S�J��H-k��6n��0��μ�q�J��3�nq���aw V��[*�^�㎽H�f���۵S}�J�\t�ND{�Ŋ��S��[���Тgu�_a�1�'����D��9]���d�X�b{ES3��
��i��Ʃ��THc��M�mĨfi*�D#�5e�.���Zz�I����9�B�~�i���	�C�4͑W�ӽ>��b,Ϩ�"�!W��D��MЛW��
�{é�����o���J�k颌���N�[E�ƃ=�&j��x_���b�-k�a�;�A�s��0�r�$e�q�s!IE.���9i�3?+8:l5s�^���w���ց@y�Vb�Q���
Ͻ�4��:���ޘ׀Q�;���њ�1�jU@��|�N��ܪ�_7���~m>}�e���Vѽ�aw�J�(+�����K����������eXȌ��/�f��M�E�R_�F.!�%��!vo���qv�O���J*�&NR��t�V�)jm �4��?��<�7))֟-��D�9�:7�:{�iS�,�K����Rf����F��L��D��^�şf�j��B�#1�/۝�-�¨|�n���.�w!8�mc<9<k��;�S��}�>�F�FF|�Q,T�a��Va�F[��}�,�E$�@P0c�\��r@�2���Gfx��`�ll��?"�r�K@پH�vT�v��?P��[j�D3�瑰�>LN��u�|��ප��,sFv�����9�S�Tbقv
T�j9�N�*�WX��HP����(����3�����tʮ��S�Y�NГ��"�l�zK%S�Q�B�����e�� �c�B�,y���K��;}q�`֒+m�����d5o�Ci��ڈ���"�B�Q9pɬ�>��R ����h��B��ڣ��~ !��^�V����G����oWJ��*#��<n%�`�B*�7Ժ���N�E�:r��LI�0rMu�����j��h�ܕ�[S\=���#�ܧ��{T���A��A�_�G\���'�(��;�x��e=�t�pD#f`[B>��фG�s��Pa�M���nۡ�1�ؚ_���M�t�2�b�*��7��E|{hb����|G��2�d+WIe�y��`.*�`�Ǉ�4V��`1������`��<k$Uɪd�i��[Ī�Q����y����F�����P*�\�G������/��巳��%��F���U��,��2I�lj~��t�S�`>nsܝ��k�1�b�\���t<pI}v��`bL���}=���������J�+�Z��O�Q`��c�_`hϥL"n�8L�?.�}G0떘����ϙn�zFr��1rNp��x#/����ixP+#�5»5�Ӝ��l�7��wl���ZȗxQS��׷�ۭ>��87�RDmĢ9#��{}�ۡ+��D�C����|ak�w��y񸩑��g�MG�Q
:=*��uZ������ ���1Ö)sT��l�������BEb���`{��^�\���l��?��x/��]&�����xI.�:�Dz�fgѱ�u�zlf�f=Q�ZY��<�0q��S�i,��mOL*Q��Wm���x>���4�`?i>�:R����V0MֆTŵ*��nZ7p"1yBAur�.Jw%�~$8�=��?dr��n�.�*d19���O�J*P'{M�-�gϱ(a5n)#@��t
?���Bc���w�s&�X�^���Wh�����h
ߘ:G�x}�O��((σ���̎�1������\_�;�^J\w���>}��T�Ɛ�����&�kl��w^ =[蕦jm�ݐ�JV��pлh`"�\��C�7���3 jF��>�y�oU�Y\1B�';,�(��y���,-a�_�]V>Cs���PJA��5�ݕ�����OQ�*`@,��/�Q���Й��ʪd��@`�Cc2����ך	�D?��C�1,���^ѓZ�v �@1X�wK�j>�u�܂��sN�2��T&f�R8oa�t�j��*8��	�pN%����mfh
Z+B��^Ӌ�+9���H�"�}�,����ri��<_��g�;��Qe+�,!n��r�I@�Y���F�t4u�ťTO�����|����9���HP�yhΪ���{`�u����9�(�a�$>�� �&-��E�r��0��c��5cg�*�,�V��Ϛ/x�6�X��6䙋��`>� �f�L��,J[g��yOFJ�þ�U�p���|�!$���C5��}ܴ$i�GS�#� �P��K���֬$F���8����Pa�B��h��M�KW���196���֦g幎.�ϐ��c��؃�,h�̱a�L��������􌵃7�'5��~ouB,����T�*�
P�����qZp�	�	�`��h��Mų.�W݌�qW��W�����N�N��ϕ��x�;���dC�ӅQ��� l�\�b{y�����
Ee�J�_��4��v���`���J�	"�a�g�@-0��Ы���P�Քi��<���Ԯ+:�ɕ������ȷ�7Q��9���٠��Ȓ�6u��� �ųj�k� ��0D����b\�mRݵ���.RkA�f�Ì�ebE�Tj?,�^�!m
~���'�v+4�KW��~# ����id��R- �'����j/:&�M����k
I�2�������j9r^��ʖ˟������R���N�Ӣ#D�O>�ic���~˃��}�F.2�"%,0��$h�S��0��c�`�BlxV�h�U8�t$!_�(�ȭ>�M�6/4܌鞱YlW���z��Z�\G&K$lǭ\������n�Wo$���T-���}�4�W.��#�e|� ��ѹ�]���փ�恙�����*c%[:�R�W������|2g�վ5��A�|Ύ���5g,<�0q$O`Ȗ)ia �'U�X]ؘ�5�3�k$k�y����9�͇���ny);��n���`^�/��
����~\U��Io�(N�
�!z���a��G�WϢ��{jB�HG���ȥe�5����"w�<��3��o����k{������n�B�ȭܪw(��4������Y=���.drf���PIɪ>il�JU:wNo�f�@-�a�FB��][�S�Q�I�gʁ5̰w��Z�$.��KX������R�x��v��%�����\l�T��Q�q��.X�Gsh7�+�+/���x�Ww�� _�T��d�bQŐ.���ՏJ6viq������b�$sN�T�^��-���qV�RI��"NȀ�  �}��(��u�B��KspZ��+�����|W�\OD���ڴ�j���`9Ⱦa�xlA�lVvJX��8���3��mO��7�6vj��%��+���p������l	AQ�4��	���}�o ��|"�C@!�����+�ٕ�CW��9�Xꢺ~�B�����JZ?Cy3�y$'�s�Z\̫f���\ת��g<]㋆��� w��AS�p|-)�Û^d�,?R��5z�>'KT?�{:�38ڗ���oFA�%�v4��dr:FSoM��Z��n��q�}%�F�[d�N�@��
��5�z(:�8�cM�efb���ˡ�K0/���2׃���z1�^4���$bVdx�*�iW>)q�ePfi �8�B��$fa�@�N��cm��=���2m�o�<�d���|�@
���D� z�J��H�qG6�h��H��+�����p?[� vK�B��e��j��}%�Ia�;2m�h�g�aw�Y��`�`7/�"xA���:��<@�7��῱�  ��QO�y���\�z�&����Md&����[�
G?Y%��G�T��z;&� (R|�� u(���]�=$ƴ�=�nx�X 4��r��&�����h�ZN-�kE++x4�	����5O���/}�r�;�,�+ :�Ŋ�7kj���[��"Ĩ��s��+K"0��  ��o����J-����gf��h�T\�s�؃�_�Z��b�휯�IX9-�"��
�@o����`M�.�bӵ�/���� <P,�ICB�\�o�Dص��S���*3�W9w�z�o��������sl�r;rUs
R��O�!qcBE��mM� C;�Fn�NO4i9��+±6�X� 3�X������j�:h�	���h�Z�<@AAO�? >)�V���p[��~ر��dD��fֆ��-=r�L5�:-EI0�NS�4�^�w�e�����Z���$�� a�T��3��X�x⓱�?�3����0�
2�'M��jܥPY�����PڱE^Y�"\�j�!d:�~���%0C�����F(��@�U����\3-�VL���H�#���H�����'��w��d@Ē���>��k�);~t�>ν�w�埃�x��Q�5si�]1��Lf*��Z�I�qC�RF��zu/�����|�ͮƇJ'�9�Mo�o���b����<Ǭ�>�Ip<w�¶�k����snW�e5����eCD�����������'�jKX|ȣh�y�|6y���0kx�=&��������	���m����)�����_��������@�C>X�6���&�g�&���h�w�,y�uQ�B�#��	���m�L�`HJ�^��9k��(t���@���+�����������7�����Ӧ}�C���q@��E\Ym=_��ؕ�$I�XI衲����`�wgR�~x�5��i�[��5��MZ%.�)^p�l)����th_0�	��cl��֕}��-7)�a�2G�fdޫ��P(�.=����4mr�P���/D�$xռ���	�&�?%��ۜ�����\|�uQ$bs�I5�"�*4M��rCw�2�b�r�Uܷ��q���z�X�J$J=<1�St�m�7�?��W��yGpW-�D^�ǎ�tEM�Z������"~��]�N�M�w=Zh��Ii
�l�Y5#��U�.�z��gB�^��镾���e�$K�����r�ʶ���	+�-�aB��0�����Uy\l�8����ƍ� "�Ϊo�����(��9Aؒt��.[ø?�鐨,����	I�.�֤="gfφ4X��d��3b��PL5?M �u��D��0�S&�w�l�V�����e�6!��7>򺽥;~��T'N'�R��0��x{\d�3��iS �a�t��7z���5�4J������w�a^�9H�;�Sz�����A4������y�y�$d��E�wnl�������'K �Bd�[����9��]y��DX��D�j/����(i}V�8X�ݐ����lN�<s��%`����F!A{BBM"��|�k�uD�M��3�.��8�IS�3��%GĿ�sn�;�-�	.���xZw�d���Lvy��Ŕ�|���@�@��(/��l&/)/+��nˮ�3� r��w͍��}��V+v	���������f$��l3�(Qڗ��_ˆ���9�q	�}���X2i�`��/c�Ӛ��c+&��g(~�G�#�OD�� ��u�+r�"7#�7雦�*r߁9�g�����}W4pe��(�5�'�g���ܺ�¬�X�M���
� ���R�#_-<��ŕ���Ȝ���$�[xᐑPM���2�K�2����h
����g��e�'�C�D|��c�~�:����ӂ�Ȃ�uR%I�X3�Ӧ�&�c�I�D��Y�p�[�a���Z;m}����6�	X�Myg~F$Dұ�c�u��c؄����֬��ؠ�MkV�D���c�?�<�Z���՞+hCXc�d� (e�`�T��-s
�x�,	9FH�Ɯ��_����D�{/�D9�>�Y����a�+&�r�D��������d��G�ݜ�����2�!Y:��ڲ�cF���'��Yu�N5r4���5`gq��8��0�u����B8֋F?�����
��@V���k��f�3s�D�O̸w?��7�΁������ۿ��p纓�U��P<�a\����w�$����)�<@�*1���g1���m��T��75�IK]����iԽ�ݤ����E��ܿ��@��4�H���XzM�������ñ����?=g���VW��z�>X�,�8�^6~�
눫�`d���z榡Z �Y�6Y�T�rR�����q�=�-�L�RM����Ge�~I���Þ���>��2���Hô+aU�~�
��Mɼ����>��_���%�� F�J�l��DJ�*�qe�ZXYU%�x�P�"4M+C��Ԋ23b<��x�^�����v�%�@l�Xz3�7eb��А�8ቮ^��u�n��Y �R3����Ѹ�p�E�Z�:N���ae��2��o$�^/S�0�ӗ�u�I_�z��
�8E1^jUWt⻒�D�*Q����!��Kq
Z�3Ԩs� .JA����v��&QZ=����s�d�K������*� �qD�L�� ӈ�M��|���8Ze�=]2�2�\�'(s��z>��|�����ֻ�� �s��3M��iN�K��@���ѳ�Ψ.%x	�40a/�����}G���}�@���Nx�6��&V�NP+:{%4�� �A�<^M+���o�[��VZ�H��%l\����f��J��OtE$�'���Hd���\Q��6�yiv���,r��O�A��s�� RX0�-�a+��8U#~.E"�]�M�J��AI2���e�׶�s�*M�	��%�17Z���j�S� 2>��05(l�i�{���f�_�f�=�Q��	�-B2��[�����<3����m�&�	m�C
�o�*�H�����c�=Bf]�-���$�,�X�-�N
㦵�R�V��,�1ľ�#U0�GO���ꛂ袤0���}�躃�-��*�������=$v��_����Xfn��E��_���'9�z��%Ƈ.lЮ���ş�)O�hs �����n$�6����b�����Zᯮ�;�@4�:�*0��k���h���U����*��|�g��˯Y�Fu��X�l�HL�I��/�1x���3���!GAҺ�	7rgf��a>?&1��nߎ!���-��E\���߮Mv�>���h+O���*���ww������P�P�;�B}�EOh*�0�z��e�����g&�1ޛ 	WV�{�6�y/$J/�a��$batJ:p��-V�Vf�o`�\��^f�+xd��G�LWb����ǈʛ���$e�jlFCd;�������ш�݆"M��naXs�a&���R��W\h��_Hr\���[u�G"�tV���� ����Z���'J�{���BJ�A���^���wbS�b�*�W%<�� �sÁ��@����r��՛�2��-��$.o��EE�b��R�C���x�k�H�P�#���q��G��I�����U��B��B�r���O��D[���NvG�
�TեfI�oQ^���D�wBI�#!�+�QP6-'g���R	UoU�C�"X�9�
w��;w��FW,�x׮Q�zT������*ou���k�G8:V\4���X=�S����;a9
Ww}_��{l~��y O�/,���	">Z��d����d���W�� 3���E�msiiZ=��	�mFǘw�JV<�4��h�L!�&�o;�+�+��1*�7��Ǧ�Vi�A�����i�40쉛K5*��i �zb�ߍ��ކx;���2�w|��S��ȁc�wd�1ur��U��56��/a\(��V��j<28�(7T=߿��p�0����L��-��$�d=�o`����a���Z>|f��)�?򎖹>�_'�8���/����x����ov��ܞquH Q?����ӣ�ٞP�{7�?���أf�+LOL�;���̌I���e��ϲ�����,3����H�KV5�q�&VN��c \=}��n�]ޖsu�Ø<z><%��,!�Ǧ��߃P�r4���)���:����O<&=1�=���p#���[������ܜ�p�l�
^�R�z�X5q �`*D[ x2����S\�FVΥ���Qӈ�MY�k��ۧ��
��&�x��v��E��Vg��!�z�\ �Q4��FS�M�'Cw���ނ�ԢՓ`�tz��Y݌��C�K�*�ЭB;��]��J�g#��G�����]�2|OQS/a �N��M� m;d�y��v} <�j�T;�ggsm��9Chr�s�b�c�&mǱʻ���{?���:K��.��rbJIƎ�m�P̣#�P��C+yُ��;�&qx(�ᾃg3�.]1�@�����E{�I���R��:��0��Q���踩�k�Է#�j�)i�P¾�Kp�w#ϛ�Li��`ھP0�.�\�r.����,(MOc+C�pj��a���	X*�cЗ4.�9lg����¡�
��q>+��j#;���R��Rg��v�е���V�	�?�9U ����M`Hz���yo�N��o~C�T�*�-��4�WJ�/��+���)dm�5_+�5ݢ��^x�#��u�%Q��qm���]Ơ��]HW3�b��I(V�x�i���m�:�.(�o�f;I�]h�h�f��:HM���S6��o$�ɰ�NAN�/p��\�_�A���#$M}
T&��..�^%�={�K�/��� ���ҫ��_;2�����^�)��& �w/1�p�W3�>�D�@���H�3-��%QJ�q>
IJ�䕅2GP&w���7��ˬ F��PbQB8;\s1��T� �*%�}� �+[�,2�"BP�uV��A��Q郠�>`�]��s����#\�!��O!�.Y�2�%�B�j�!�Md��>��jJ�h�\�]�� ����y(�0�U��}���-��,O,�ｋB��{�q"/�����^z��z�ǍE��e�>��I)��y�mO�h�Z�dv���9�L�L�t���}�27T���pR�k��E�2��Hu�M��jR�	앾b�։��}Ǌ�[��^�P��t8����l�fw�3�x�*k����5��Es�|����!&Ϡ�
ֆ�{7��T�ºH&a�(�b�y�tqQ��߅I���"P"�&!�c��b�
uTA����M O1� �*U���ƨ�2��3YX[�=�t`��m�`�g�	�DL�o�@��� �A�x67�u^�4���M�Q����kb����v�vF�mKy"@�O�	Bw������ ��xU��z�ý2\���|l@240�0�{��&JO^����'f�XV�&����$�4Y�fbU?8���P�a�vi���u,�5� ��/+��V0E��8����c_v�-�G��z��}����W��u*[�!_���[{��M���f�O�s{c�����{+���w)��ဪY���^�g>�B��h�;yP������߾�Wb��e.dB$�^!�S&۠*��~u�9Gn�'�+XL0I��������6�і���(��PF��=�Z;LQ^�+��62T ��o�E�"AA\�Ä0�!�A6m}�_��ۄ;�۷�������<O�Do�8�B�Y�R-'c�Ϋ��<b:L6��H�۞����_�ywQ9nF��n ��H�:v#Z�Ê���=s��.�H���m��a\���Ȝ�!0]��#[J��#�෮e�]���jJI-����)V�v5S�����N,�E�&�g�t�r����Ŗҕ@��֠ف_A�]��[M���Eဿ��Ӱ+��E'��a�����~��*Dd����v)"wA5��I�T�t�ͭ���u�	qwϭ�_�l�g��ͷ�J���ů�p�D�|�_��9��ہՖ �W�
G*�8ѐA��:c��E�A/�)lϦ~�D�H�X�����k{�BƠ '�WB���Y�q,7,^p�Y-f5:K2nu[����c����)�׉�N�nbt�~<�
�z|:�������-#�7|��Ab땋kK*n��i8Ӯ|;��ٶ����$]*C�z�	�����`Z2�L��$��P��]ȹ{њʹ%��MP�V����nA`n�y'��7ǙP�.��$=栈?�t˭���Q�V`�� BNQ���������_�Ụܖ�ֵ�u6j�~���D ]$��p��+u�Q� ��_�5�{L�q��w���QJ�Y�uv{�����j�jM� :~�'���v�#�� �9Y��P�Q�8��Q�醒�h�t��v�ɶ�ݓgR����~i��9��f%��¾�`ƏC�]�ﶇ��&�|rݥ#�<͸+:�K�����4�RFV��P��\��va ^CG���?j��2m���4Hq~w�|$L!��� �8G�?���<k��b$���\�VE�-�·��LN Y|4��u=��^lnTl�!���.���/l@E�t���[�0G�CNB��ګ-����"T���M���P߰�ƈ�!�sڳ:��?�RE��~�i�w�İwſ%E������Y��V�_����k2l��{x�t��A�}��Y�9?O[׽����
ኻcC9E���������#��t�y�m��B��"��z,_n��tH"��h�"�j��d)���W�*�;��L��u�4�B5J����ٱ`q?{k 9v��y��X{�zש�2�+3Q���Qab�Bp�WLї�-�0����K�X��#�F4 �˩>�6�0��ʚ>�F��P�)�Ǉk#�A�p����cfj���w����J�׶�Ԑ��ɷ��ܵI�bFJ�Wpn��Y4?@����M5��lZ�<5mIg�O�"���"���O��u��?�֝����0�m���[��O�H2���2�4� �G17 j�5��%��ZZ�`� r5¡�/�5�S�A�`�b�lˀ1����\���nX��j���k�:^�~�Xb���B������l]rO�����"8����=_�6�(���^���qg�`U�I��J3^�w?pObk�;V���	��YмZ�.��h��w������,A�AԖ���J��l�6�{���H�'�X�ɬ��Hҿ���Hޔ�nZ�?��#�����;LI��2�H�EF34'�򟒘(y>�p�퓁�.�"��0��莱LtY�J��@T��u;%���b���<}+kP=��_�Ph�F��������=�O���x���/�Ak���5A %��X\�Y ��Ҫ��#g�D|W��A��1P3m�����r�~��N�Ψڙ!@qȦ.oxRߎt�Sx�u�蔴��٤�+vDՑV4�vZ�אB��aV� K��~B��۝7�-.�PT��"�n����ZX�V4T ݭADԝ��(����	�SH�ׁ���)�HcI\d���ROʆM�U4�xg/n��P�����ի_[+��g}GX��D 3z|+|�y)Ǫ��%kR������|��O���t��w�_�6q�x�L��ԤQ�����W ���+@ �R�5��up�>�ҟRF�?�iC]Y��@��;?���l��N�7-�w!YX�����OX���ܴ�dǙýH���BSn���=��U��d,'�i�ѱ�hh*�@���u�I�� 6[�HH]u��q>6K�.6A��\�sORhI�=�	5	�[�\\���.�.�H��S��~7+���*�/1��՞����X�	;�@2�:��ao9}�9𩪢V�v������S��(��n�e^��zbo�n�ȯ���o�&�h��0����*�����"o���Iݿ#|q]�#���H�X"�];j���u �� Hg(0�{���������#�Q�s�<�x�H��F9�C��{g�i
�@��}0��;µ��Z��X�����M��LFY/����t���a�xS@m(�=$�ld�&�uu~��#���)���>�hk��,Q<�e����09�EP��fp��Z��ǅ/�p<.�:��O��Ӱċ��1�a��vb�K>��ي�^�c.�	�38�eg�d���<\|;9Đ�6��R˗ ��7��{�'��g�,?\!�Jwa^�JJ��6�ĵ�"���D{r� W��R�1�2B�+��w/*����@$B����Y�ApI<�d�H6����I@�0%�+u"��:AR�˧b�q��^�}d�di9�<���ft�-tM�ګ��9�j���1t�QH4^�%�/aۣf�0��D��:��艂���9&�6���m��&*�\����O]�f=�2���_�-[u��G�bs�
�e��D�;!q�t���K�)*���b�����{�� fR�/<=}��~��lA؁կ�����zM��6�]�-ײsK�R �t��z�{��|�U�n0�(���J�"��E�xS~�j��U��ymU.�V6M>��<��	p��ꚰ}�j���.��Ǐch���r�.�=<"��{ U�=<c/�/#�l#�e{0G3���=N FN�3�0�K~*���n' 	n��6]gg����1{�����JG�0�E������2�D���^b�gWӜ �-���zΓ���*%6������]oZ���	$Hh �U��T���HkrZf�� =z�h��V�V,�o��L��FRH��+/+"��7)h3?Vb:�5�<.֔��Z!N�PV�@>�AUxP�v�����]�|j;��\�rI��RH�?K1�<�<0R����ddg�x
��C��:C�d�~�����a�kv�1EM� �_X������c����FutH�ӳ��9NJA���k,�Q/]\d������f���*J�_� V�:l�l,0tE7,�F3��}����	'u�i��O��}���Ça/N���S���� ��0��Q��]^}���d�p��['��'���r����F��N�v��?�m�+�N�Y��q�"t�X��_^'�lda��B���Ah�;�\M�7;��M�j��A�c�� �v$!�2�Mìj��]ͱ�j����)�o/��$?�Z�%��$�KUC�s^y.��b��^����Pt�}���1�ʓ%a�@�- �;�>&����������7�������s/Tj>K���R������?F�QWok}�R�<�}�"��-؜��`��ېˊ��iqz,?v_Y��۰�;�@���j0Í�@邘�z>}�l�k��^E�X��9�?���O����;.��Q	��f���ݠiJT����x,,n��Y�8r�i	
�Q��
ӗK�c->��v��!�!F��/{��%��shY\�"%5�CCGv�|�`T��i�5���4�{kS3ʥ�N��H�٧d�����'M�ѥ�������8Vi���@����c���O/Kc��������͉���,C����Ua�בR�V)��nș/����谋�6�x��;��k-������;���+��3l,yi�H�lNmֽ$�<J=�-�1k�rK��q1��A�q�ґޜ��(�Y��6^�U�X���j��n܊���Fh��$�N.k��*$��z�v��-ڌY���S$5�AR�o�"���G��������43�"��M�p{.���T�:�΂+�E��}�iM�N��o���1�9�~�C^��%�h���zIb�O1������&#H�� [X��a��e��l�����N�{%v���]���>��n��wM��-5��HI��Ѥ(q�����vdǎ�Xo9 N���_����R�r6�B��O08	���Va�fWR�k��v��Y#5���d����$@��E;2��~�)X�j*[���@uj�OM5��əqqhL]���O]oY��)JĕR�-��:�a��YL*��FփN?���'����P��{&���Y�W��p]�������TH]D��tm�ò�ʃ|� ����B�)�*U��4�}�t)dLt�W��ʺN)��
� a�pSưK����>5G
���{�����=>i�;�3���s��T�_�N�8n����[b#8]Cğ�����{J�>�4)n�+)�sF��Yjk;��}ز��|M�������`�� t��p�M�'.y/-q����n�ӌ?���l��"����s/�CչI5/оΓ�挵ԃt�mP����@��囇�59��\p.�sY��]�t��EE�Ũ���e���~�na�{/�G����nJ�r����絆�)I��2`�RW�[���e6�H�~����CM)�L��#�����$���M~��8S	F��؏�H�f�W
�g�3#�����Y^�ͫQ��4�JT*�8]>`s4����W�f�J��]%��ϥ#{Z�1����*H�}I ��x5i�H8� 4��5͗�v�W��Gɣ�A�/���V�ȿ���,򢽀C���t�9ň:/��7���Urj��Z-$�|�����m�FG{\/�N&���`���lhL��P��6�`��d��u�k�,g���̗c۫�j"����L_X��p4~��wc׍yv��3�4�Kx��HzO�'e"�t�W&���0��ǌ""7�W3������	2�~m
�g7����(}�X��Ĩ<UvsŇ"C����Ԉ�'v)���t�o�ʮzj7����L�E�9  �X��Ś�?����X��V4%�])9�����f������&�heɛt�P�!+��*����f�Uo���6�v�ͬ/�Z�Fi�Fr>`C˛)�H�?�m�|M�*2�%*&��.��0�P��6h9���I�^�z��W y�6������K��lDx�7�r�8��I�]f�H�K������,�j����IM��uki/�iyiq��|L����Cy���çh�Hx�󀟞�j+.R�D.,=ز�9{��,�S�A�JL�W���<����z��JG<$�0�ؿH$��?b����o̦�qݭ6�O�9k$�3�J�������1�WT�#j�ł!��!� ���������f�h0��J_�/hѴ�� CW�j�7�i�����[E�p�2A�🎞�(�Q�|h8O����M�)��@UW.)^`�O�&��@�mT���Q���S�Fp�^
��0%�U���^x;�eĝW�UA���L�3��R�g�����q�<����Am�����ݭV�w
�Ɠò:W�Ύ���ܖމ�Lcc��6x���;�������,+�\����NZ2Z��9vWx��FW�oK���i�$�w�(�bI��N:�o�a�������o�
�����y��mn�Pׅ�
����k�FH�P�wס�
�� $�8�[�d��4��Aa�씁X�M�_������Wt4(^�е^�"�&@�˧���mI�n�����ݵ�h��������F,,��G^hS}��ð�64�ҟgU�{�[�3.t�[������6M� �
���I=P,.=�� ��&�Ex�B�+S�"�ġ�#R�m�.!���q§�e����o�t F�[��\Z��G 7S�A��&����޵�Ȼ��!�Y+w:��K�$6�։��p��l�4yҢ'��ڻx�Y/����UEy�G�cZ�����+ǁ3����N�bH�QU��E��\3ۨ�6��D`��`0^��|~�ˡ�D����:�M������r�I0]7|G�������ar�Qۮ�&BշOT!�X�"��$s�eEƚ6�^�2��垍8�}��f94fN�y���e�:'���ʅ/�ԩ�w�0l�.�z(�^Ad�f�^l!T4u��ݱpo>}�렛#!�D�-f�z��߬+Y}C'c��@�,N>�B��Cf�̟=J�[6���Z��
U{��<�(P��^��RZh��u�ǍN-*s���~��xd�2�	�u`|����0+.Xp�����*�w��Ў���U�t筃�O>�S�l.��U=/���5N��ډ ���ed���J;�
#�e��\�8J��HƖ-��9��Љ~�f����+Olhr��%2��b�1���a?WY�D6/+2��FE{���S�H�E�J��*Z��붮�'�`���fh��t���q{�QkE	RͪoR�#r�Hƅ�����M2�o�"�n!9EZ��s �՞@�üD�m4���[�o2<Ϧ�xu����sc��P�i��vF� ��"#�D�Y0l�O�5(�{ݍv���u46\�~'N|.��Ҵ��Z 2M	�k�s2�yH6��ʇ�n�9I�vF��$2t�j%��eDf�v���KkO�K3k?�.��V�ZM��~d��	*��q�� Ru���y�~7�u>�+�n#*	+��|E��͝���>��t֕-�_H>f���h���qe����˓�n�x��L=Q
9��Ѝ��(Yvc��<}`�Ǵ\)!8�\�tNT@���$lJЭ�22��By�y��w`OwyK��r��e�u���\�E����Ύ,�pP�����پ��r��zlɎWd�ko':���ݽJp��a3R�\�~����h�&�K�ڲ�U�LkӼ������6P��	��A�wVA�sI��T� ���Ŷ˾���F��dB��L�:��W������J(������F5�d�4lA�r�r��M���	<�耠V�*8�d����s'RZ�a�������[���i���识;Fպf�Ϋ���㕁��z5��B�����+�-��~�d ����o~���r�aq��3Es�y�����S�Ns��Q��b7%xy�.oen7���(�8k�.M7CfS��StO�q�(,� ��Z�rQ��M3b�q�i_-\�=�0�����ϥ�tŻ�Ё!�D�j���qT�����r�J�n��x�=C�\��
�?�3�e��C6�uY�a.�9odܛ�����>gg�:�+���^h_��aҬ�ˢ"�	�<�E>��rq���T�u'�p���}����h��?�zB�d�+TC3�F������Hpq�)��;"�H�DX�f㢮�<��w���Jl*�Pv'�?�g�HNA:o�5�7�;��Х(׋i�f���t��%M�dqxn�<gu�,c��C�1O��x��}���<�2}dg:74V�c�c�8,����� 9h���8�]Ͱ���-��ROx�YJ�A�R[��N��G{2NyT�kNL=�h�����H_6��b�%����^�H d��f�1q]*O�?�{�u�0�)�Xҵ);ޓPd�0���v
|u�ɐ�v��3��2�0�|�U���	P���>*����2�6�2W&ΞK�ON16�������Cg*x����5*�ߵ�-�8H�H���Mt�W29B|�d��I �aI�	{�[L��9�p��UC��q� b.��0��er�DV��Xg��w]_���rzo+���'���>��f���CkE���hy	�or�7�"p�pPwT�}������t�Eb�&{?����O��t�$7i?�Ǹ�G�����W	6Ǯɛ&�ap���E^�Fߢg�������s�� x��6;~&�ș��*s,�C 7��M^����l
��v�XsI���J���8d�3�NV~Z���S�Φzc�y]��`s�=� �ʮK� $�(�;/Y�h����΀��4�E�g�&6ѹ�\��5=�~�������Y}�{f�֑Fg�?[�[��yRYp��P���{�o=Bh{���'�QI�z
��P�Y鯓�VY� h���	Z�\�.,	�
t�52���
?dv
��OX��K����ovLj�$@��lL_��ٝg��;s9	�}��WM��j�]u}N~pa\����mY�8��9�w�
�WYE,dr2߀��6����"\����t}��u�h=de�J�� �1��f��x�&Ê#����8>YVu���b�O4�+�;���hZG�(;(�Ah��<��nn���5(�#��G2`�ڠ��½)�K3�Ur _���$�bp=��[n�I�����k1m:� *S`��$��+����1��LH���\B'�Z�[p�@dz����Q;�p����*�׮�|������D�hu���;0-���?�;8@N��"�$�� �_:9�K9(�,��L���>��>	�g��M&X��+q^�9�'�q#���&T2�n���-=�8����=��e�w���E��+�0���ʏ�ɵCSt�*E�.ʷ�2�h>+�Ѐv�.��9���I#~��I
/����D�%�Ckk��d�ˇ�n��l�H��r�7.�C�~�=0��/χ�l%�ުs��n�0I��� �B�čc���]*2�>0b ��:�8z��T"���e����b��]�56���oX���kI�y0züC~��8�5�,����Ƿ���U`׈N��S����.]r��
nK�݁���UD�)30�Ǫg�J��0�Ǥ5!�������W��ԕ�[<��Ĕ2G����Gph�B�dy�}�"\�i{��j&(������}%��8T�,?%��]h��	K_�"�QP#^�AI�M2�.o��".�R43Ƥ�D?ݖP�#�0�-�\e��XF�x�2�8�<+1�M�$-2!w����E;!�'#@q^aiýd՚a9	��<��0^�t-�oC����l�v�J�#@�`Ugѳ�/F��4� �s�	O�@�вm�ziV܃ܣ��p���L�,��z��	�B����)�pXJ�����^M�)
��q��%%��]-5��_��CAK�i�r������8T�OTQb(����=�A7'h�k�{),�I���;�~�+c�q6EJ�J�G���l�4ϳ�x�QN�@��q�H��m��B̞p���AJ���Z�%�&�Ib�Z��>X�4ba����n"r�[�Rvh1����1�h������;%�8��ө�6 Ďm�h�,O6r��������+�+�H%��6�W�������2��7"kg��+x��~��#�U.�����ߝ�K��2R�Vag=�<�)���JEఱ�i��F�O}� UH����[M�K����^����\6���jb���cZc��C��Ш��M߶��(~���(��^��!J�_�}�U����j�d��S���8Ż�s+�3�u�)���q��&�$��a7;�j�����oo&�O��P��b�W��&G�QP�4�r�(�~a���'��t�.�,��Ǭ����]�]>'���<�fR9j��?��;�fWiIi��!å�K�`�`l����f�[4CQ��{���>w�D�lMH͛��!� M;�Su3����0��dX�a#��2�/Φ��s�ҁ�[��b[%�A�����d@�s�=���[�UX�ĮG���t�X�U*�v��l䖯Qb򷧳v.��ڳdTD}��B�l[�n�)�o�y���T��z| s.5��O0�%5��ڴǃ��]>��Tv"���܍k�д�j0��ŋ���x�P��6��7i!J�@>��DϦ���<8nJ�[�z(�k�K��U����1|zF^l�����n) �>�q����!��M��1zO<���B��3r�ik���r��O�]v��Ԓ��#�+S��-�o�vʍM6�|N��&����ϱ%zPy���j* *��V2�Ƞ��\�l�پ_��F�[|NeN_�v���QuH�u����V�*_:�i��ƈN�L��Q��D-/t
��8<�X(�S� X�~?kD��:x�:��e7��)�v����^���&0��@%\'��ώ�_T젫z^�\�EeƓ�[�}��\�
=,���dQ]��Z�Z1����=F��E6��Z5`x�-P������r��	w��y��H� �O��)޲7�kN�\�&Κ�v����
q]�t��ݛ����L"�.#1~�ʦ��3�8;i�ŏT����������2!I���E��~�R��2p����u��r��iP��y�|ж�M3Z
9��*�9B��W+cM�{ ���K!�`|fn}ι�W*�`�HA!;��X��3s����a������l�СvSD�T�n�ڔ��:D�ߡ�A���5��[0fF�x�sn�z��(��ﻵ���o���T݄SP�XH��P��W4 ��m��7U�7���@:�y�]���VB+�D�h��}S��ca��f��� �ᔪ��mn�<[>5�>e�^���p�����:�e�[׵�B��Ӏ�Ŋ���#!-��Z�8>R����ĭ��p�����������Z15;}�2�Jp/svk�s�����:�Z��Є�`�� ����eIS"�E�l:5��1�[�C[ҮK^���rDݭ�B�j��I���I͝b*�U �M�z���G���@�0�;Ǆ�`a�E��v~�M��gAt��P���*s��K��:�7��t�]����y�#�H\.�F6��ޠA����QU���ܿ��K��bw�RT�R5kK�Q*W�>k.��\���W�	��'��L����I�G�1���H���N��>b�	��2H��CF��^`PE0�_���]YƳ��RFw^���J�՝=�� |_��tlQa� �591�$-���0�\'Uv��$���%I��ؿ���q�k�ċټ���<�,�e���{H2�JgV3��Ѻ-f(Q�� k蛃�w�`<�=��(Z��d�Bk/#A۾��ײ��7$t݂�;䤏X��_�K3���h\w�a6����Q���.�(IOUّ��P��jۓ�.�I�s�+!�N��+�7�^ ���T�`s�װ�6�1ξ���PȞ?|�	��N��&=+/���-JybM?bz �d!@�%C�ZkV�Cl�O/͆�D�?k�#W�ؒ�:P$���B�`Z�/������(ڥ�t~J-;. Кk�a��!Xc�+g�p���>5�~F:��\�1w��E �:$�.!΅�;CDl�H�V���["j]��z��s 8�c	X��VZWE^k�&��G���b,�U��҄P�t��7<NO�r6�66}`�y6R>�sUs����EΧ��������R��ށw�1�V���������o&1ن��?�ֱ)�E��ݖ!�ʨ^�H�x���@S��A�"C�	t`q����E��>�m�Q�=F�D���+��lO�El���᢯F}��4��[ե�	d�Ԡ0;ZٙӇp��۽ce�E��Ԣ ��%u����}S���l%4'-yH���G�r�7H�y����J���U(�~���\�Ǒ9h&�ι�{}�����F��Bp�+&�	V��=)B0�ajD�z��Χ�Y�{�FԾ"��w�R�2fk�2;��#��\�}��������32�~��4��w��h[��s�5Iu�3��WC��9��^�㚦G� ]��b��?9OƉ����9���9?W�1�m�s�\�����[h�{��У�G�XT�s������JtM�L�qQs��2:��#͙,Hc]�ɀxj@�Ftj43����=��1���<�S:�13d1��
ܛqS�L�������Qv<�
����B���a]�5����!/N'�)�NC�5��4�(������@��H����1��7���T嗹=�d��cC�s\���������5�`�`B6��t���nɕ)lX!���J���h� R�&ܬ�¿L������U��_�?{�ôF�U L���J>�+�_���W`P���~v�`DO�Yhu�y��}T���P;œz�`��ѲB����)�(5�)O�G�v��;�>�P���f.�q�����l��o�	���� I�IX���p;��&{�ĥ�F6p�s�F�����c����k���J�l ��W�FU]�ٞj�iE�\$�� �8"X��Ρ�s�^x�$t�1����(*���5^�n�]tY}8FN��G��t�I�=���^�¢E�z<��J��C��X�,��16׷4xX�52���i�)�#�ŬGƸ@��00��y�֯ ��D[�^uhF��w!c���7R��/.O�V�6@|��|�5%j��I��~,i�]<�m����r�����C�!���I�����~L�l^�"�5e���������.s��iP�Z�ՠ��$�tO�>'��y\
-�wSG_�����.��C��/�~�_T�}����2^��;�)�׿�n��~��li�L�x1�޺�%��>Q^����Э�J�Aii	�I,+� @GpM�ɻ�Ʉ��Ϻ��|F��]�F o�$���b�U9��nJ�F�J�`�"-k\�:c�Y�?���;W�Sl�G��PC|��
F�*	�3咀��b�;l>�y�+r� P���M�Ɏ��D�R��R�"��yJ������(|�q-X�}h@�T&�ؠca(r���_�Hz{kf�r�^HP�1�3�.���P��asΑ��@����ƹy�2����!��=�.*=���K��s�x<>L4� �=�@���,�2o^�3�\zE� ��L]���\�5�gH�	�)jp�;�3��]m�����y"��g5�����e�������������ǭ��o�<�$$�ؘ�bw�s�w���t;5z*�@!y�<��Js��V��� ���(#�����.&~���,�Ys����!4(d�����XVx��'��X �3���]���L=zf �9��8�$�ge���$@�<DfRP �n��auο"����r����>�;J��6�O��v�*��]����*�>]�M�E����>ܧ�a�XD�cH���u�:�+
7�P��D�YׇC���(�-�]���K�8~�Zr ��(mhc��߸��]�|�Eh:W�4	��,9}�S�t����|~����0݈�Uy1az��kdhQPJ�����F�q�m�,<�Ρ� �׾"�T�¼�"�GE�o9�J3�d>|��5��i�7C��-�mxT��ə������Uƿ;�b?i.�e�c	JO�!��5�nt���6�a��.�����J�X�4�V�ϔXLה��o2���kl�`�'φoSx滜���xF%�~,'(�?��EZ�Xq������LS�<ע��o�{���Q�]A�cc�ݬa����z�Īv4*�g�������m&�yMp&`W	���&�;ء�ʚݹ�!?���Mx�	�}�:�R��� ����M�dU�H� e��<C����������\�VX�=���<./zk2X,Y������e���^+=�d���	:4P�[���@kp�q��rDϖ õx���t!��'�x��%Eh�#@�0���r��+�=��.�6`�C_vP���o�gw���������)���o$�o�c�S���uK�Ƒ�v���L]@�b��i}`WZ�,pڒ@� 2Pև�-L�����A	�f�-��\��P�;|��(Y�p+G^������>�>W��bG�Y�	���������[߬.- �W�sP���G�C����#���̪l5��=C�������F���8�6(Vt��˟�-����I�~�@�e[���Ƀ}�x�����4�b�s��89�������[$ikDVRq?�lV�2�
h#���5,��&��fZ�:��rжJ��4��LA�<�(n��bO�+'E���ϙG�!H�ڢ��Zy32��,��uu�D��e�7�����^�/��h>�.$��9�=�!�H�Q-�:��4�-[U�E��)�����^����>b����3 �ņ���ݕ���@�!��v���A������LT��yNJ�M�`�ު��e��/�6N"�������;ޑk�H섾��sJ1��T\i�Ý���E5��{k�k��bۏ���`�B��d��ѐ�ߊ{�7��(�Vv:��Oqx�~ox�f�� �p������q�!/u�v GE�L��ł���M�E�[�3�s�+�s[`ӥ�f1	OA��ff������RޛE�' ��X���P�crAV��f~R/U�s�&(���}�	�c�
�7�CՊ�8E%ѣi6y>�L9zT�	ǅ��=���S�[�ҩكӧ��
H={?؃ӟ�!�<+� 3�AR���m�BN8�t�9��³�����"��oz���w���)w��*���D`�O���@D���*�� u��:�vT�_��#�쯈|�d�i��4����l�6�����R�|��*oz;f�lo�{��k��Y<�������<�o�-����H�p$3W�7&�GA��;]�@	�Չ�s��>��[���#/sDcm�������.>���Z�ϔ�9���x���S�JD�Ԗm�_�RAgv˂7��I�vc���{�U氊.wO�J|�k憃�Wm��g>?&�`R)âd�|�V?	��e8�<����1zz0���K�$ee�a1^ї�i�EƐ+pIc�] wu�ä�HsFQV �}�+��+5�c,����%�*��I-�ezs~2��h���]`��b�o�ukX�m-�<��^����rn�Q@��*T^p�N��\��� ?s��_�9Q<�NjT��:�2Ӌ�5�w0���e��[�^����K,}'ʗ���������$��V,j�)�#Ӂ榁g���GTu��^Q@o92�:�w��l%��� �՝�<����q���
��xo�.�TlD�gw$I�X?���$y�>'����O��K�#�� �{�tǼ��ݨ�m37�Ŋ�{����5��q��C��;.�/����;��ڶf�X�F�[Uڼ���|�u�K���#�B*rY��ft�?h'.��<�6t�"#���uV/����z���A#�s�Z�d�?�!��@'�i�lXs��������U�f�~*P��g�A����e�2�"�@5.���N7���d+�E|m��<̳g�xFr�]�M
uߖ2x���[��N��㭟�{J�{��t��"dwr ���6����$jm�!�
Ia�ǘΤ�B3���?�=yj�.������G�uA��liq��_k����u_�c�nJ��Ѿ���\����ͧŇ�^�xaB����WLa⢁b���4JuӵFW�x��E�?�@�2w�0�;�2�z<���Շ�dU�Ȫ��H[��}��լygXׄx���#��}w�!)��������ƒ�;c��Ro<�:v�[+�$tu��9��<c���;<
@���$�3X���GE���7:��|䲂3�ⲵҧ����_�������ܤun4��Kh���_�P0����ǝ\	�l ��[�����:E3���{l��f|9����W�.=����O(���-���q�g�|��h�1J���8�~-�6��*/�e"S=ѻW(U���*M�,���k�c�yEKv�����=����MU��ʹv�I �%�*���ٻ1���B���;�1�jg'��;t�r�a���UXڎLV\3���֯�"Ԋ 4+4��Xp��f�%����%I�:1$0Q�OΈ������;���J��	)f�zN���:4c�&�c�G�&��WՉȉ0l�3�RP�Xv����v8f��gp��V�H�Κ�٫zx�=Rkur�n�8;��W�."f�/�<w����،TM��������3������lĽ�����Hp,��)#��Ģ"��]F��%��̺ݶ�B�@J3��F�*͇Y�=�>v�mx]?|����r]�6����;�Qg�����x��(\�g��9~h�k,�١ ��bL�[��grH�* w���]���6%r����b%���,�"�R�b��Y����N0�=u#�ZqIгf�AKt�'�e3%�V�mp��l%_&�W�`r��L����qHf�'��
R���3U�����K�\R��,V'�T�N��lph$�sE?R��n��ߦ�Ax�;���������!r�7^ׯ��l]׉
�$���;|�F��|���*o��qA���k�R�][sK�)�9�
K�v�r�?�.�.�[؋�.w�?��t�
kg�:@%�p��\�ș6��ѭ C_"�#x�2oR���6D㿇���$Z�.<e/��t��P�w/Q������������셖v-��y&!�k5�ş� 	�R̋�V��E,��7J��:�w&�h���5��V?���B��6�$�yW�Kc0�M	���[�ݬ���qD3�5�S��9�⤛B�G%�=���A (ͥ�3������[�BċF\h�{@E�h#�z	.��E�=�+��'�B�<�jz�:��>������i�[�׃��0F댦��˕ăw�¬kY�����(
���׫S�r�w�%�h��Tu����X�so�ɨ�l�uu�cz`)�u���)���@X����d��;�7g$��wR��9cuM�v�,,cu�V��f��p�~G�`�&�����nQ�Q������T�A����}Q`���j_�[+M��J�x�����J��>��Q;r0z�Y1A��Ѿk�ij�����u熣!ă�Q����	x~-���O^t�xQ���ShCc�l���MF�x�*�{z�H\�������s���{��d����e3�΋����\O����.I-*�Y&��d�9��۝��v<k�MU�_�	%��]9��w��`��T�_B�ehh��雍��-�X��v��4�Fa@�)7���M���\Sh���������M�����6���EV�kɋ�|���L� '.���.f�99��^�=�׾���/���R�<v��Ih��aݓC�3��q~:��x�܌�37܌�t�KY��7��xc�$��J���B�B2mc����m+�G���.
���`/�%B��_c�)���Ƴ���S�Jԟ�9ZgR'��}`�]��S����$Oa�u^ �$t��mV�x���2e���n��iM#���-�]J3��Pq9!|�=��JuV��;���r;!��f����Yo@^��;�<�O�96�|�`�1j��{�ȫ��wR��jX(��[%t4(Z?����2t�	�'�ʽ��(��(� ��`f1�PX)-Ch����ǳ>�y0�D�t�)�Ծ��*��]����B<�?�X�3��'u���2���+�I5��g�	ưFmKN[�V��I)�W�'��	�ђ����=��}es��O; ��%{dYV�k���GL`1S��b:9��ݸA�=�g��P@T����e p�z���VKɡ��V�IoA>��9���f���m���J�g�F�c��H\vA�b K)�Ev�M�ԁ���ΛXKHV��m���	w�ď�N�RuN��/�؈h�iޓ>`W'F��/u΢�h� ��e(!؍
 �H�Mk�(8��Xa�q$նde��v�-��4ΘD,�m��ȇ����a�=�0�pK���C��������10��B���<5w�q�����Ɉ�F��73�gl�%&�7C��B*O����$�dS���.*�s� 0�bݬ�� @�7d�$�`���,o(1����i�}�KE\ĳ|*�݇�*�X�+�uE0�\��?�6����s�}4�P�y�F��* a��Z_L�$��������]��,=/��0�D�V,�!~���][�n	��_H��4��`FHo������;�{�J9M�V��QI&	[b
K�@�x����t�as��2AF�
���SFa�t�9�4��!�(�ɽ6��c]�6O��5NO��I��6Rz��L�8�#xnؼg� � �a�J��$I�I� ³6W�d�c��mz�FT�>�ϴE#>0���r7g�J;�f��0g�|�J4�cjW �t����4:����Ϝ��"1^F�EtH��8T���2�'�O���%��7es�hLo�~���o��.��W�M9��_#K*|U��h��}������r�F�4n���)e���x�,��j��}��֖ ���|����q�c�[� �WÄ�i �Id��\���I�"��_B�3�ݼ��bZ���1�C	�B(t�������e�"�a%�jӇ&|�u��yB�#!Qd즪멄)�>�Dva��쵰O�x �rR87��H�q����;q��T���aʹ�1�)��� ���s�� ����Q#��K�T��@����߂�n׳�%_ᵃSZ�3����(�k~b�^�e=�������P�ٷ��}�@E���Y߄��5���q�� ?`�B�+Ψ�!K��ԛ0k�
��՘�l����IL����(��@��
xrq��L��rHu9)������,��/^?���fg���#��GG�Kl�I�Tw��26�;�9n���%5M��������b�@��3b�8E�"%�j�(�͝���4�|oZL�c�
�e�3�N��l;à��o7�<��>;̐I�Ԣʊ.�`�_����
^c�-��+ڣl�Ʉ��e7��t�Q`�s�Zi��� ���j3�&Gł�	|�܌��j¾�*���tNoW\�b���.�\�����T�r�?�(���?g�ʹhЕ/:��W���a����l�
y�9��u�����P}.Zg��nFfW��)�H�W�s'�rV_&��- �@��5��MA�WI�G�/-k6F�m�e!�w��0@SR�O��넺[Ժ�4��}M���RU�׏~�}d|)��a���8���o���(V-���.�T��&�-��rg���(����s�O}`S�Sڸs8V�WGƭU>͟���PKhS���$��7)�GU�G0�I;�b6�g�E���IE֙y�5(k�"e1�X���l=^�/�_Sm�՚L:�w���ח���h��[�Y�8.�LoX�v�x�!�3��g���=�6�;�')׎��ͬ
�x�VV���e�u�zz,p�s4��n�^`�3��	�; �+9=R���є��.�.�R�C<��/[J8����һ���p�Ө�7 �w���#2��N5
U� �������\��D�0g��[���!���1ϑn�=$��$u��V�W��k��kB�$p8�`�D�ɮb�ê �w�O~�.J��I=���V��%��l"��Y�v��#o���c^ߌz����U�T����v\k� V�K�fGk4[4�1q���s�#�TN���1��iF0���	�V�-��Ph1�v_vN5��bS�=��'y��-%�#�2Ι�On>@�4(���]�u���� йc�r�	m�� K�/�$�qBC�D6+�]3��n�u)2Q�^:���l��}�!���s�����
�S��-�g���N���si�U�Y�a�UM[�IA�z��X���4�b��C%����;�a>P][im�]B�탟�2����}	+���t��
Z�d.6�hv����r�z<$��WEyy��!��X�4O����	-�$���aD��	�@���j)��"*� d
��6�1ʖ `z_�8Y@��h b4��p�(ϒ�jv|ՠ9Z*P��\ī���h��&��{���/�l�zH�����m� ;��ҩ���}J}7�X�0��8����~���^�	D���d���Nvv��-��B߆<8R�J��@2�.�J��2���OG����yB-��.����G�Ϻ�T˒2�R��m9.u��`�1M�Gtr�����BO�)��U��G*(4���j;��t�v�Z����#:���:w��e^��&O:-P�B};�4��mu+:�t`�ͼ�7�a��������)��CKr^+�p"Y��\P�Z-�I+�L*�Z���h+>ݻt_��m�S҆�e�Y�v5̛�
��>�E.����B`�v �6�T���?ݔ0x����*��g(��'��W�&�W�n᳥[,0�tc�S?1ȭ;�[��E���Y`�g�.Z�d��؆���Ѓ�Zf���h�"����[H�2X��{�41�B6d{��h�ȇ�р�|��$��w��N�6c�%�T��G��q�ZҼ�:oC�/��<0!p�ɖYQB�!���Iz�9�L��rA]�N������A�3��w2�^�u��C�e�Zێ�8t=Jh��|G�h�ވW^a�����(�}��@q���Fã�m�֑�W{��'y��o5)FK�r8�2��T��>$)�������a��[@�k�`�����
�܅�!f5�*z'M��a]����������(M 	�W(N" �a���~*(@�}�c�=�22}��lD��e��?I�7JDW'9�D��N�o��R�P�'hӥ_d�~ٞ���F�1���ђ�2��;��;iƃ^����ṃ~^�3d+29_�H�J�D��4
��� m�bvH=Ln�F�"�S�j����<�`��}0�2;��A��3�y�iz��E� 4���Ǖ�)	�sћ����@W�����J҆I����j3������N�a^#&ٛ S�=��t�A&k��)���-/�� �\��MJ�u�ǓUk�`ޫ��u������5.�|���`�>܏{{~�l� g"TFnOY&!1�}�n�D�(o}L�/ i��Q6o��]7#��\�m�,E�o�ձ�h����?�:2Ζy4���~�d�4�5��D���_G���%�o��[D{�Xk��D� �F�䣲)R�ڧA�Z+{j"ڸ�gh��@��
��jzm��E��I�:�c�ԥ�eq���`��"	j�M��P���@#T���1��i���nE��B��SR�-.�� ^>��7 �-i2�b��=�oj�cI3nJ.��{���������"�{�q��&�b�o�]��]p����y�WUG� ��Z��r����QW�N���7r�����Z��8J��A���)C�ߔw���^��F�����W�_5��%~?��	`F9�.�ӅQY(���fs�rd�_�sn!�h��+U<h_=�6�4���5�O�́�~�fc>a�~+�aq����v����x^��3���n�yN;5:������#%�W��e�Y��b��`�.�C+��G�:ÛU&���O{Ĭ�b)yz���脜+�~���9l�b�=[`��eg[�;��pՊJ{��~F~$
��]U~w��,_��r�r��;x����l>u���/�R�=T_s䧣�W>�!w�:�{��9L\p�g�X��������Gru�&E[�_�fN��_y�0����x�� Qcr�y�VG1�Z�
�� r߉�f�BV��\��#K
;�N(��kVy} +��R�^D8p�sAW��Z?��=�(YB|��f��3��b-�[�0H�˴-��'[�*j�@:��3
��Bx+,�f����z�\$�K�
��+}��$sn��q$�R����!@eS����<�R�%�����}K��2����[��a �.[��2�%,��v�|T�:O
e>f5������	�����Ai�p� �Z3���Բ�{���WB�-�?�=����`���f�Ԁ�����9��B��m �����>�����X{`�$�#��`ϘyդTz�ۗ�88���Țdv��|���%,I�a�}$E����V���X��\�Z��c����/�_�d�OS�d7�~�B��뀄���6�.{yA��Z,=���!�3LS�E��Ǒ��Dkj�K�m��e�z���7��G�˨�Lv�j��T�rL�_���]^�[���;g�Y������<X�D��{�tk�$�3$�����!Do��"5��r=��D|�ȷ����L�3�"��O�{���P�o�J��;��v�~��rW�z����=��p�[���	�	0��3����Y��E�,��� 'R_���ObG���D����"�1��Ib������7�+h�Ÿs�3�)�l�3F7~���ތ�JT���Q��r�n�'a�ʮ�{������{����ژrH�4������~��Q���v�B�-xE��]�~����j�~+�lX���h�ʵ7��"7���j�@Wf����KW;=��@ȃ[p�<�:��	�ۤw��r��!��`��:�l6?Qo��\P�q%�~�!Y��ŀ�ݗ���3�W����&T�(��F�l�|��g�'m(����g�`��V���Y���OJ^�Gƀ�PI�/GK@س��  ���s��.̾3<�\�b�f�7l�ErΚ-`GW˟��brh�9l]YI���s�h����j~�ȃ��";�~��h�6?�A�F�=����bJ�V$��A�k�:�� ��zz ުcG��_��|9��?[wl�ze�m�\�f�	WpgA���!�ic#e�<p]���?�3��~齩GMT/Œw��`�ι4z�Yu!�b���wbWԩ:�R�N����S�.��L�W�q�RED��+�D���#����Z� ��N�s�)���h�´4�:��ĶC9%�����8?��QT�@C+l�`����W�7<�+#y�����]���O�V�+6���t-�Z��׏D��_��%)�U����O"ܛ�(,b��ͫ������DU�	+7a%���)S�h��#)jѦ����O��l<���c?����bd[y���!��/�����M辬�J$_��j�s�TYWг)�"���M$�Ԛ������o��v��,��>��E�j�X2��.�I,x��3�:f|�m�,���x�|1_��Y���k�]���0m���k��j_���Ä�S�bsӇ�� Ɖ��Dq�Q
��;G{��y�<�*��V"���3�B��_�A���D�gԱB(|��6}5��0��<�Hl��%���W��Ȩ�x�>��|+{��ݕ6Ы�F/X�/��4f�x4t�����F����O՝ӡ_ص)s�3����P�_���ԝڕq�W��H�rr���|�&�����%���A~�ip�g�
h�f�B���q�8��0j}etT�e��s��+�4lpӀ��z�k$�CKG�#�Grx��R�G���:�l�5Q�ΰ���ޙf��T��w���wIf�ϴ(�b#.�E.�ү䈒�-�)o��;c5��YB�d���h��Jy�HT�	��o��7�FO�xVq��S#7i6.2��<{3���w�Ԧ�W�{�.Ơ��I���E�|u�|�x3g�F%�8L^u@4İ�8v����6C�#�`��@#�+%�/�e��CK�?(�"��(Q�w]�+�Z).��i�T���.������9)�	E��� �ڡ�%���_��E��1*X���M?if;�v?U��F���~�0`�\o44����aѢ��@���Ľ�v��4�-����(��:��8��N�(E�E�J��he�x;I�zLGI����w�:p�Q�5D��g��-��,�A/o)�M�&��o����6?,��H�7Z�]I�wgTr7ݪ��kF�@���H;��r_�}�Lv��3̓ŝJ�d�x�e����z,=�� �V������ /<�Bz���Ҍt)Sq����Wzh�D��	��Uz@�:��_����/�_�w5z��"��j=�7���%�a'=�;�$��Îߚ�8�j��<<��ay;�΀v��L=�
�p���^M��{/�o�6���1{}3n�������%���7�ܨl�ܞ)��f�z-k0�JT�p��Dѝ�{���ue��ȵW��G�ު�ĥ�N���TL��	��4Q1���+u��*mQ�w��v����HN!
{T���Rpt�b9[��X�n��Ȼ@�pԨn���X��l���)�x������yӠvh8�e��$�s�9�0�ܾ�DM�宅5A��0���c/�$�E��Ww�~7�'%�-Kx�Y�&�8}��*�Z^:0�RΠ÷������54	F0�	��O��M�v�o��KΫ�#�h�].�h��p2�8���O���OVK�n��P�U��yh2w7�����˪����7g]�l��׍�9=m�#���0?^�{��˿�6
t��~�1@<W��^��Z��h8��uy�o��{v�d��g���4��/��QV�iZX�7�d/*1�q���@��ڻM����tZ���ĵ��I�(�$�h�2�R��0�,�7�`0��[F\�QH�(4�aw��m���b���̹_(7�S	��-R��J[g�rW��������ED���k�������nc�C�+j���'��}�G� -VsN���q�c���W��3�-�7�����Ge�'j��]l7�<�q��ԽR��b[	���@�:�$�8/��Tb~��:}���R �s=p��?5D����L�te*/�B�A*#)��/�;t�KV��_="-71W��6V���ڕ�vB#vy��%����#�m]�)W�����i(�'n��@�H龍�������GE\]u����'��p;����~��+�"���<���p���!8�4�N ��8t�k	�����@H@"�>��v��tY3�/�i/~��Cp��=�7 d��{�iů~(oB����������E=���#���W:��D� o���0�(��-�E�I�0��aE58�#,�F�2�X�0��ʭ���1T���m�:݂����D�R��u��y"*:�4�A�wj�#'-�g�zWI	�A&�2�pQ=@C'�ҡ�([��nw=Mg�E�78�a�V��(p�D������V��~�!��|̶�K:>]zh6�mb�
8mt,��ɠ��9����[ �,0��dN)>YT٣&0��9출	���{�dd�7����ϼ�|���u�}|���,Z,����A!c>_͗�P�����¸���[�nU�������ʏYV���(~wB(���7��Z����y�E1Q(�׻��(�:��b}#�G�����,��]=� �W���:>=j������)��[fӾ#��÷��������΄���tQ�Gu�%,A�^�E��4�UEU��l�����Bn�$�� �p��#W��"�&�tr�~q�32�j]��qI�,��Q<q��v))�\�Dn"̔��V��l6+�*i�V^�0��x�2�����	ń����&R��ߥ1G'�iٰ�+�c0#�v� ٽ�B��/�'��wQ�.N^0�Az@z����A�d7Qz�ܳ���i��a��d]GZ��7��W'�Y=�CHk9�>{��"=ωN�O��'\�e�k����W6&<�Jҷ��e/�����¸���j�p��4�̣���-ĺL�
��"_�K������;��m��"��2�a衤!��q�f�(E.&��zG�bf&�]pj$�h���t���<}�+�n�My�Q'�L�w2h����9zށl�L��#�O�~Tmi}�$�}_���<-h8����F!Ȯcҩ5�w@{�1�:��$)�qU aw[
|�E�{jЍ��~�BťQc��i�?��	�M􊚣}׬�`�0H�� NS{4��O �WW�o��s��9KJUr�߇7��5L0���Ǩ�i����<^C�������1�2g)$��oV�&���qM�c����RӨ��E�	ݧZ=I`�?�M벇� gAP�nNE������8JॐC(_�{6�!Y`���ؑ:$��l@	���T.'�d�V����×v5x�쫣��/�;vӮ��%��X�c���YW�yP����5�O��
l��){so# QGc�Y2Zz"�R�>�^��A������fC9�MF��>Y'Z��1{0��	��$q=���k���G".� �m��X2�"}��1�0��Wh���K��xh�9�>���'�������� �Vd&"�Q/	D:�7�������Q#�U���\�5����r�яXR�)F���E��&\k���H��oL�^�ӷ�_������@��LO�	e�*m�n���i/���@V�����33�'����/��OC�`�E�'�E�j��|�m�Cm5G0�r9O����"�i!q�����;DE�'��n��	sc�bSo�*��/�*�Y����!W�'�����3�ɞ����6+*�\ef-�k\�?�xG=��.�!�x�hpΝ!�eT)1c��E%<����x��8����h�@-v��Gc�R}"ㅮ� 5��'�i&�r�G$x#k�=,d�M�(���
����&�%�2�S2�P����uI,bt�}�I������e3�p��?b:�"4
$�	y�Ӝ�WL>4	^���0w�y�K!�[$0ψ�̷�kH�Μ�7�ij��ұ�r{�^��޺�л��3�����+#�m$ux�o��g=�r��"#��jn.�[�L�:���pd�O�_�p���ٹD;Qj .*"��_-m	d�=�8��n[�NH��q'0�~�?�i.x_sD���)��6�n
�M��Db��	XM�>�L^�ZS8b��9HD�N�9�Rq�����x�&�>}�E�a~���'�v����G�)s�L����}�ڮ�bl���<� ��#�G�F!��V��(�M�t$��)�N0U�P�h� ��r���T6����K=��pbL��Pp������e5�D����4'a������K��?A%�$?��קM���3�Hi��rvm;S��OP����Fm�y��ͨ��%X3���JD�D��9�`���_��O��+�%���y<�t��B��*�&�u?�:23]�ī��!Y�6���v=����������ŉ�iv�U�~-ֱ�Pc����]:=�#;��@�D>����LW֥���RL�;�����CQ��o�0LѼ	���nL�Ku����DE$?�(��\��D���Γ������+��'a�-�.��ƿ̻�?77�.Qzy��%jU�<�-P`K���1���2a-�'Gh��P��Rw���b����B[�)C@A����̐��G-�S��&��W�J�89�������w����/���Ę�&����s/>�_")����<���a�̞`��}c6���/e�P�d������-�yC˰0����>rW:׫Ԯ=����h�HK�B�(a#3�k�I�&���6�$�D�.��Bxw̼ƒkŠ�twY�7����k��G�Z7x���%�|�������v)I_���KX���=u�:��T�E��˝g-�Ѱ�`0�д��������(���V���Q�H��ۃ������)��X��u�44�������y8�w7�75Q�t�g�[Akt,@zɀܑ3��&��r�۩��ӡ�ť��1�q���r��)��ǆ��cə�jbA��T+Jhi��u���P��j�4=l,օk)ݪ#��
S�t��SJ[]p �ֳ<k�dbs�B����p#��H��dN�fQ������'`���K&"��.>��F�������vJ��+��(;���
a��;����j|�;��Nl6)9=^E���@{L#�W5�A� �%�t�	�-������W\,�|��c�1O�U�AuE���ØD'�8Ke<�Е�(����`稂�6\_�&E�W(���l�\�ތ?���T�}����[:?`�1���<w�=K+����cL�u�7�#����g�>Ξ?��w��1����t��Z��z�N���4����`)E�/��!Y[��T:�[�EMnD~�I'Ik��/��p�Z�IQn%�p��v�%%�e�F��5�R%eՋ]�)�*N�Į�>@���J���d�Y� �&k%r`z�&SN�f1mR֮���0������d��MoeɆ�:������L�of��2&���F�h�]� Fp=31L"L��A�Sߐk��������7��[�%��X�+Z���0Τ����	�A�X��A���{���l�[6iH�2$FwY�C�=噇'�{�\���0m����6]Z
��Jo~x2f^�8o�$��R+h�F�>M2��+�4�����4@X?у�dhz���_9H��GR��c��������M#Z}<	�lEb��{�,�?�x��O4� �M��R�4�j�:���_�}���V�[���b�/�x̻��9p���t	��hc6lhf��qY̽�h��LO�$U�ʥ6��4�TZxq�:Aϊ[D���)�l�y�5� m�%�e,6����T���(�=��[��&ZrH��݊h�W`h_�r��X�UMp��(#%�$�=��$�!!6NEq�1��D����L���:��{�0h���ِ����o����^��,�}�(e���r� �uk� ��r��ӧ��#��)~�`���V�2M��w�7R~/䉞��4��Օ�A�+�ke�?B�}4��x�3��~4ϨI� ķΪ���t
ܫ����o2�^�w�y�2�W9�b�婤<�hG�X�ʯ�y��H��F�y ��u?����+9`�5����T�y(1�^�Q�q�x�?z���5�J!0�쥌�^��ߦ�$�"�w4s�o@S�*
W/ls���	ao��|Y,�b$-'�k	|U��_m������'��k�UW��D���k�óB�5	������4
ڣ������m%��,��D�f^oB8�87�l�����x��w{K��=�>'&���w��a��xRp��C�I�.�;O�DM/����>!e�,t�[��n�1>�Q�ε/������g	|��V�F)\�]��c:ʮ{ڟ��ޥ�5��0����O�q���aE���j.�/�aO��EqQ��3q&<�����n��9�c`�z��B(�c���gH�eķ�H��L��~*�ھ�.����+ (H*�m����1ZB����3��s�!~���0mV�ϟACT%�F�1�B��vw&���deea��k[��Ͽ:wo/B����+��fk�Sه�������x[Ѕ��B�XP
�~��AfX��-��������D���r���'(�i
X�rL�qH�;���a��G(q���by��ȹ}%%��ÓI��z��1N��Zl��S�K~�q��;��~�"gp-u4����#��҃5���a�w��,mQg�W�ۮ��f�A�:��6�Zw�0M� 2�������23��J�� �~�\��}E*�]��6:QQgF�x�PC^�A�;{.���kբF�SЙ�/�VC{�x]�<����퇘Ww��%����|ͳ혏�t�.�ZE�D�z���z���
�����v�����KUhb��f9��߳jB�X�V�錪�Q��O��7W/�U0L�?�m`�野�i"�id��ue�1%0ډU���0��O��Hf[|�x���"���
/@�Oc�T���F�7Xk�ҠO�����:���Pی���O�ӊ�g�����֨�P8��,Bd*��oc�]��*uEO���DP��y��S�n53��oZðV	.��yf��7�����V�� %rd�$�l�cإa|cX�X��ҿ�~-�r��eht^���ȸ�)r[��X�.�0�a,����A�Lދth5;�� P�����,��B6�w{7��p���n���1���F�I�; M�µ|<^���cO��*s0U�$L'W�BE�n-#��Lc#!��/�E}O�1� |)�5�>���Q���&��S<��h��%��gP�����p�[S�D.�KI���G'+�4��1�t ���$�r��	h�b&à�L�b�
�r%��c*�����D$2p:8j*<` }��[�������ʾ�ch��2Һ�{\�q<�`Ĳüx�qST7̀;؜(�+��^�߉�=���1��Jy���%�)�s��sD�-�R�/�W��rĢ���u�&� �T8U=����?޾�4����K~������H�Y.>����=-op��1X�}h����Ѩ��X��i�]>Ђ�T�WJ�^��@|�� �ir.����^Oa��s���c�2���/t��uj��XJ�=�T����_�/4�qpy�3⶛�}&���ߴF�b���8��ԍđY�6�ȼM[A ���HR*�Rj�Y��g��,�9�����/�$��#�̈́a��򼴉�U��&�1�I󳠗�I]��E�b��"q���^p?��0�h�!|SY�3��kt)C�8�b(�
4%J�j���K��w*��+L��:�Yю����-��pp-hu<�'e�CG����E`�\�������਽�^h�x���Z>�T�}�SE�-�!��@{�q�|U�!��u\��(	���Y���k����'��Ռin��e�p���a��϶yH�kr�����-�H�U�Ls��u�G\�dSf\�E��=,��.���6���ڞ���>��k�ݷI��(� kl��M��y��I���� ���C< �ND ��+0}.��ɄU&s��T�@������:3�FbR��8����a,�c��u��s/P�����o@^s-[$p�|�UىQ�;�p�6X���c͆��U�l�.uT�|$�#�7Ƒ]؊k� ��r�2�bhToQ�/���z� t��d$+�w�>�q��K(hs�HR��>W\��)������A8Q8W�m1� D@��Ç^�����f�gGI���J�4�ᝉ������2d뤸sl�b�:<Ѽ:q}�$�ĎQ5�E���kGU�O��6&���恬6ڍ�I���]��G*G�-�w
kyL"���)&�9�����ʋŭ�(�L�N�!��FhE�f���Y>/YD�;7W�B�O�n��~%��I�ٲ,D��^*<O5D��"�,̺ovU
��@ؿ���fr��3��'�K�N�̒5�8�-���g���^�7�0������4���\�o,=ދ�.
h�8Os�	*�no��V��;��"��t��u�?t�|_��(��Do����U��`\��0�-K���M���1��ճ$��TB�}��=�Y[`{�唃�fرuvi-j��%�����z���o �ķM�y�@��N�zٱg���m���6{',�=��=�}l8:4 ?�掊�*t�|�Y�4��\{6ˣ"������7�f_�&y��>�jgA�u�aj���p��fiݫ��i(0��P�a�٠��0����-�� ��� �!����Z5�[ǖ�V�}޲���عj��D܋��N3��{o]�"��|�����M_l{P��$��W@��8����u[��j���ֆ>��^ߚk����.���Q[��(XH�xi� ����u�]Qd�� 1.yCύo=f&��I�����^R��̓����MQw��������z�WQ2�P�T���ce�p���N�'����,�b�F� ���/Y��j�:#O��$�|�԰6[����M�n���&QJ� Ժ�ѢC
�z�䆬��{���[��%�#�����X�O�C��)\�%�tr�t�^/1[*0�����$"��*R`1vR��ʀ�êqPoz�L��'��lX�W͗�>���	 w!����ƺ�����PZi��LT�'��@���G�tr�X��ח)h|\?�wYpz_�?��t����t�$W�u��V;�\wX]�S�q� �	lB�לa#�ª����E=�O��f����σ�P�*�IG#��_܆?���R�W�)=����j��=ćMݞ��uI���AĂq��dC�T`����P�8֐
�����T�$���^,%=i�s�t�k�
�͙@PK��
���FU:�5O�#لݞ��#ѿ���0KʈW9�k��P���c�e�b�qn��b���`"�5#��c��Y�38��3��kt�V6�1+ ��1^)�g� ��B5?繌�=�r����ŗ��²oF�(�A�z��.�BE��s�<���U�X1�i֩N^���D%r��wn�ءo�r�s0���׉�1��GTAs~�ݤ,�U�Wo
�l��J*�:��;0aV`�|� ܊e����w��pS<B�V�]�e���㵬j�\KW@WǍ��D���E���C�$�����Qw�U1�ǫy�m�fO��q=P�A�'�_����%l��yb�_� �4\b���s1���(:��'=�������?\�z	��7�@.��P(1�*4��p���I���+*I.u�qV,E���!"$��B4�oND�j�Fj��#���Mb�|,��H�/����;�;�;�
��sI�Y�`�ѳ$���/
�|������Mp��O_��C>�@<j�{�➵�5���]������@Ѽ��L�e�k�������s�y@$��3bX	�	Ά�?�%��K�a��8}h0���h�H>�<���U�o2H�n� �]��t�?㢴�9E�6��F���=�L��L�ʜ��d�j��h����Aw�{��F�*K����'3?o"m���`�p�4���S	��)ݫ�C	wv�ɴH�,az����������~��r0�)�#Q�N���N�W�a:N]L�f�����Fq�uЁ'n>�)~�	*��!h���)y�G���{20e���@�w+8��חW���,@�2�|9Sf����%s�� ������s��K`d�/5m�j���h5L!2�G!`���b$>��B��*j�@��"�YHO�~RS���h��Iv�����j�,�� ��_~CCz��jpBˇ���x����Ǣ�K��P�װ�V�ҫ �;6Q��ظ=��AɭU�|��j��������{(�g/o1l[�<�⨬��@p����U	'�ѫ�\�`�-�����]=�-�@*��	�1>⫞�eig4��r���\��F\$�*�p���N�)R06^�T��Ľ(�9�#=�	~����]lW!$݆i!Iz��(5$a�����ɅG���`3�5����bx�sV����@<[S��,�ñnzys�9�Dt_���Hxr+R;�3ԄĪ0o����W�$@��*��C-���9�J��UgsFq�~@s�7�U�I��.��l���%�2#yl�|7|>�k8��\�{��9�N�E}i�{�Y���-R��A��~]Z�V���� ��I�v,�	�}���mE���}e='�<m�A���1�}O߂:̯�s�Yг�7��p��^��Д��	l�8:�Y�����s%��G-�V�VR��^�_@�>�=��Y�/����J�y@���{�V�K5��o��@�&����0x<bv�@v���M0�#�9x<��U�J�*���̐C`�3U�@"�v������Cd�P˟��l��Q�8M" 7~�L�T6����/�m�]J�e=A�!~�j��T�&H7�l�6"p.b�b����k��O��&���ż����#q�I:��D�N��2:�ßw;�pI�/,�/E�FE�࿃����:�R�G�]}b�A������c��) "�(����TR�/^��sS�����Δuw⴮��C��'v��t6�03��������Bk�N]�W�#㺩�N��n!rwC�X��t����K! cM�ɷ�}%�����|7/�ݜ�����A�Bf���i��t�o��L����1c�*ki;�kjp��9U�p.�>���s5�y�r�Y�>:��#�;��r���Ŋ��P�<�$fRڠ��j����P��\|P)A��B<�p�<�����q_>ɏuz�Ƚ�Y����|<�b�����kl�X=@m"�_;L�����u�i�ga+��-ƛJa\qA�̕������Io��{d'�y�����?.�z��h�s�QRȴC��X�##y(�d�AB�O���+)�}��g���<�n��@��]���u�������'H�J��I�W�<���\2h&�*��Pt�����#�Q�3��dNb�͎@�⚰w&-�5�͟�K1��w�����S7�QH,xW��#J���jU�hя� ��!��x�/b�g�",�&��{�ZHn�Bx��x�o�Ӗ�� �
��#{@����7=���L/�/�l����-�o�Fb�lega&J��P�ARۈ*s<I-ѳ�T�xB��-W���M ���LD���!5��sRs��������*yp9�/q}�Z9[:,�����Y;���ԷX\���|M���eO�r�����ߏ9EŨAn���	�$�{%$����M� �Z��]�����8��q�v�읪�@3�p$�{��_�A8�GI�h�{�����P-?l��Jb0��ᡎ�:I炦�Nh,ȭ��FӬ�"[�R޾����Qr�a��"��]Nf���4� �����R`������g�Wa�vr+�X�	� 6�B��]�J�ٞa�,t��ٓ�)6p�u�5ԚG.�L?\P>c�"�M�iGkv9��iL�b���+Ĥk�!B\#�w���u/mJ�_(ʷ��
�<d1�bV8�Fh\\'���~09��Ԧ��n��ZL�X2.����	������:?c�]��v�0��ǰ�(a�� {P{�����̴N.rB�&��8�"���h�(L��l"�_x�[�/z|�������u�|�8c�5���7!_n����dw�������&�8���a�4I0��޵W�6��'�G6zf9����qH��g�9��y�;�s2�<�����$c2���p2�iA=��K��Xw:�Y%�V=94p+q�7u}`ԫ���{s"6�2ӆʆ4��{�׻�n����h=W�͠4A�.}�� Ɣ����Żc���$90-��#]X�C8�^�Q"��_7�S2|���?-�Qݺ��.�n��ml.|��b�ɝ�$��Bp���5�M8�]$@���_ExD7C�ˎ�R����mПw���.��y�����z��o�m����ʔ��e(YY�-��5ǉ��/���V4QY��dZ��A�|�\�hX1@���ۭ5pL�t�y����H�#L�Me��GY7D`�q�$_Dw�e�o
{�y�}a��_��x	�\"B�lFA�£�ex4�l�U�U^�
�RvQ�2�*��:�;b���\)��sڬ��D@u���&���&=D��B�Un$?o��j0���I�f���4c'�Dd�0[�l�א�ס�)A:C';�d������£��v1�)i(��E���t�`��"�E�����z�^MSM+�����?�'�-s�g4�]1��i�u/�=�G��}�v����Z���Kj��eı�?�)�iE�o٭��6�&��	�r ��8�շ��c��H2:-E�����u��[�˓,���zW�aU�0���j�5=�e6�P�H����q�G�F���c.�J��^>S��y��.�[���=D1D5Dۅ�؊���
(h,L�E�i���n�ĝ<j���ɞۗ����N��M�S�� ���OӇ�#(*�*�7QW�7	ufb��c����i�^�����%�L�����[B���k����+�p}¶��{_�c�� �݆�4Y��b�W����#ߔ8۫�1��).�/�{�t���v?4�r��=�����|3������_ke5?H�v�p����6mRw��e%�Z�]r�U>Jxu��rW�9J4�O��c��D��׺(ypFC����ua�^,�߬+�;���C(/I��&�F��� 1�<�y��l^��_�U~�}?���zve�m�4�M�������v	e�
T:2è�	jm�4����/214xN�L�GK�w�|peG?^ˤ��#��0@p6Qd#�����H���+�In��5���痪���Q���+��Y&l=�r����s��it��Ʒ�y�I��F�S`�����c[;Tk�Oȋ֥DU�o�~)�i����wq�F}|/TB[�x�A.D���{}�"e���	�U� �7���R���P��t:<F
���K��C�q���"�����dYbDb�]>��h����ҥ��-��$���Z������!v�fN�g_b�)J[�q,6DL�N&=�`��łGw����-�� ��5�W��ڇ��G���}�Z�yk�wB� ��AV�'GvnO�qZ����E�,�=��)u�:.�s����Ir��M�?��YV������5�3gnT�ދ�c��b��$��iOj~��Z�x���FS>o^��ُ`�b�h�h	��R .���H�%�����;&��-ё��$��?�Q`������z�ݴ�&��yN��Z��(�J�XM�`��1̹"JW���  �O���B�L�Q�7�=���Ou@�Sg�
��\�<w(�L��gu��ѫ��?%A�`>���PN0�{"s��b|^�
�-5�Ej2S�����\��ٓy�S�o�����/���}��5;����%����=cR����>g+�1_�Z�$*�>[������p���`���
d
�6~C� ���C��u�_@{];�H#�ޑy y�8���/*�.��֧q,���8���PWE��	��3��XF�\��	���`�
?ޘ����<��)�a%x� ����JX��\j�I���:[��H�&E��y������*���6�ogo"��]�%8h�ޠO�� 8X���bV��1	��J��9ޓꊊ���R����ޫz�Ky#��I����Ni�G���~���J'�.�9�)~R!A�=%�M&��Z��+�~F���SCa�����o���}�&�LZX��)l��H�P��}߬m3ld͌�}��K:I�������i8!���(��2|�������ȫ�.3�R���k�>;P3x;�S�!�"Ih�~��G�����ϯIk�ܒ�)�1L�,STF�p��m�� �SC�ػ�?A�C�7N����Μw�4.�ʻ9�a�:zqk'l��y:����������PT���������zL�M_����Mȋk3ǂ����-e�V�h^�r�u�=ZTzu�[�p����|��ZR=�6m'd��L��^�,R�6��+ݺA�a0���2<O�����䈒n�Xȹ=���D�(l5S��6,n$�y������f�;�'ê�0���U*�d'��B�W$5:kRߨ���;6��&�o>���hE��f�ǉ=�<����q�Q�|�`N�4�>��P��V�=��9��[� 횪C������F�=!�>�];��b���h�-:j>�X{b4μkȉ�����ԓ:��Q�w/n��OE�l����Qİ�<{�#��_ɿ?q��>2˦�ҫ�@~�M�<��	�3��n|XR�D'����W&
vp972ܘ�bb� �5�2|)X����B��(�Y"~kE׽.@�8���V��Dh\*��������<�� ���1��������2���~[�.nW��i��nȳ��o��h��H
s����޾A{IC��^^t`.1;��,��!��̺�.# ��3��Xd�tD��*�S��V�@3q��Kڈ �o�����/S���m�O:v-�[S���M�@g��\������2[�P�|�c��I����
��-��'-⃉����?f�G�f�=[I_��g��\_K"Z9��W�¸��SB(r���9n�t��=^I5�	(<����2���In��e�/�Q�@�a�G�h��&I���P-��I)!�f��C�BT�
�n~����b�ٲ�$��2.Q}�/!���!�b�������^�n
����k�~f�ut�K�D���*�l��y�����%&tQ��%�R}!f'��
�R
�˾�����5�%�N�X�>M��s����.����s���$��C��[7�ѽ�]��#z|S��_8�wP4�ѐ����eY�Q�����S�O���LA�\�f* ;0��IB�����4ybN��8h��w�縺�|��� �4�q�ok��#��4�m�x\H���d�&p
�K`��A߻b�nЛ���Z��J�#=��	Jz���X��#�$!�� ���QӐt�h�3bNfw�b+�P�S�6w����6y/4ura�yfs���ә�����ʓ�?�GwǶ8��<�Z�@�E$��Cd�l�x��[���?4�~��EB��xd|C��qw21u. QS�è�"��3��<�AO͔Wūe]�,����f�G�kC�J�7�����P�2�aX+x2��~%sS�y���33c�����D~�������w�컊�������;�G #�7JV���b�"*� �S�jڷ��T͑�Z��^g�o���m�u�v���Ql �EV'V]�x�V����Md6�Xz�'�:�>.�اc� U�b�}Z���駂��ff��#>̔�1sU_<�F��<o�N�/�tM�"��u�O�z��*>�}�Ud���A_1wt9n�	����x]ҩ#n-�`귍B0{F�o�r^�&��Dw%�exfY1�0����{8��;uW���o1�VtՆ���X(�o1��=7Я�1��־;�/2�P�E���$A:Wg;+��J�2�＆l(���p�C(0��_�ػtݑ Q��
N������pî��^M?�����I�U�.%�!L���P¤���n���6�"�M����ԞAe�����">y�tc ���L[��RN�N�b0_,�Α7��L� ֟��PFe4V�@T��T�AB[p�HMr����l�}�M�xUV@3i~���9�9L�Q)l�b��P.�����J���lL��0�]~��Ac��:\n,��r?H)y�z��3�۱�d0١�����sӘO���z�yL�� $��7M��s�d�-�W]ĩ1ʾ�[6f �ϦҼv y�"��/���H�`�g]�����u#	0�ֺ��p��(���Vw*�G\�����↙I5������� ��)d���m�ZPq��8�e#�gW�V'�%Ǽ����`_ĭ5��x�	Fއ��{�HRLq����cQJ�� ��ST�,�q:�~�Qg�gm���{/�������,�:W�4{)zi(��4���^
Ai�Z��K�۾���b�rL�m�S�Tb�XKD�3W���l��;�n�b������}rU���h�wW��N	Q"�"}��f+Iu��\;����n������z%s��Lav�ށ�!�a3d(�2t� Z�R���h:&h�KTI~�ŃA h?��C� ��s ��U~�֋@���)A)��#��4Gj���f����Ȧh�f��!m��v��+���͚�	$\w;P� &'�
2����#B�v����]@j��g
uoE�"����8�-�����|}ZEO{���(���%�6O�",fFb�5>��ӡ7I�����`A�	�ުL���$����*�]A��*]��Ã>)�9�ɺZ�5(��j�!�q�B sَ����o�"6��L
~��*6ˣK��z�]w޸�(:��S�j�������	*��}-^s��":`�th��j��w�L2İ�4�^� N:�|ɜ#�u��� �}jŮ�A:��sCd�UX|P������q�-�k��]y2b�Ơ�A|.m805�,�N�:%�]rU29&��|�%\�,�>j�y( 2{�.���կ��S2��@q��mY<[a���VX��Y0r`^6���`?&t+���� ��N	9�]�Z�xb۶M!�5y�c\�!��X�#��QD�M�_[�zΆ�E�,��lym�D��Ҁ�NXOh�����N1�/�t�+
��1H�}�
�m�5'r{lͺ.�/�M?i�O�n;�GL�1|�Sg���yc!B'�:���;u�Y��� �!*K%�x�	D+.l��5�ِ��7�������`�	�Ͼ�k�E?{����k�5��,u,�}4����-��+ͯ���3�+��(��U*ƈ�[��f�?Iކ`��Ii}&<���(�a�2�!�tU��6̐�b��1'8;�;����8]s�Y�9iwr�σ0��~���.�]�5d���=#�Ty�(Y_��TS�5|.E�_�vh�� �r
B\�:�z}XM���||�3H
��V������td4 �R��|�g��d ,��������#oMB�ؤ�C�a�Lz�Ӡx�VB���.�w-ٶ���J���jt1۞lHL��NaW�2��#jH�B5bl�9�#�}_���m�)�����DK�0<�{��v��3:� ��b�	�U�m��Xf�;t:�ER?%>�7/�ɋ�����x�Qܧq ��`54@Z 2�]]�W=�R�4����W�L��)v�\��Ѩ��_��)��x�*2�=�e2r�˂	�aYt��M�P�ª�#2p�$rsZ��J*��T��+�T������04ĭ��)��b�Ԕ+?I�k��O�c\�0D�����U�Ϊ$NɁ���ީѴ-�yD�6�Z�k���4�8.d"�|��^?��NJ1{-����8|�$�mU,K��*����dOYv���������r�fr�T����4A�R��k<A�q��$���ܚI��1�,U cCz:��!kn�v�k,�d8Xi{f_'�U���'� ���!���֜ľ.�I�1���^�p����m��F���3�OJ��7<�Dp�ČC4�[�6�̞��ޑ��t�Wi-f����KίS����ht�nM�0�u�Q{/:�N=��@��P����e8�.���z�|�c?3j��5�� �LG����		^5���7�B��/mr��a�]A%&��]���d���
�R��Zc�}�i�5�`r�l\<Д��X�p���ܒ���bAb���G�3�c6c��羚�ZH%kL�E,� �v*���ά��K��Z`�e���LI�	*\,&�Pe��M�¹��ظ�+2��E7b��$�3gf�I�	81�\۵�j��!�_�,�e���[�У܍�£����t>2Ay�J�q�*N�P�c�m�Z�����-�y���<�9+�)���+����qg���Ɠ������� �����U�M[ɸ�J�{�B[�1T��"Pd��#��ۙ8sSr 1$�C�w�?)H�����_\��*�wm"9@(k0Ȃ˄$B�*��Ɖ��q0�o� |s��f�����'w�9"j<NIV�)aC�3O;�̌�x�O�i$. �����	�q��� kkB�料e��W0;#:Y���a�i�<P%�G��e�)�۩-�Z�0æ>)�%S����XW|��#]Ě|&���[���p�0"�8�)����d_���lӞA����8@ߣ;'+��G�� ��)��m:|�ՊK����tz�w��$��DI�#%q(��'�'"�53;0P�()5�b�)av�����Ij�?u���_�7;�/�.ET��3��+�Z";{v��~�d��K���rWȾ�^ʘj���9��z<v�xU��"�7Gg���,�(��V�{zl�c�F��j�<�hb��>�)8ar�j$os$�h�)Um"g��(3��)oJm�1w�Q�cD�Z�O�Q6�(q ���x	�4�u�V�^�U��j�.U��[�2�P���4�#~,���Ok�覸��(ڔ�x�K��V
�LGu6�)�a���SWNT ����q��i���xc>/p�V5Y�$%�� �K���O&/�p���;��V��$�
�$Mi�0���DAd��@NV���LS4��e�Vd֋��-���\�c(�D
�2p{�k��ls�Ȅ��w8��[1;A�^��W�<i�1�bJn�	-H�_.� f1T4%�K���a"�����#���ڊ�E��}�j ^8����z�)0k����ҧ����p�r;����&����[ũ��{��ۥn8�d=��
��D���:�1_��:���=޾�A�08+�ӈLfI�3w�D^�`O��I�;��[����r�e+ZC�3h�|1C�Y3ƈ`h^W�I�9��EC���}��o��<�[H�������r^vNE:��u�s̡ӻ��^�ߣ���HV p����H �yc���90 �"�6��|��sϣ�^��h^�f��0�New�/�ϲ3
�S(��M>t��ؼ�CC���jg�����̡Y���%2ӟ�>��-k�Pr�q�|�K�ҝ��=ծ���v�%id��[� 8>��戛x	�:��C����bȔ~&o�d6�/��:�/C;o��j���5�u�A�>i�~�PDf����Ź�s	:��'���u�7�	�f��Ij�8,�� |���~��r�6c�����.8SJ]*%J�f}уBh8vE1�F�l���p� �z8�7�;�&�Y��cNn�^�"y��	���R;��C}�4���mہb��zFy
��{��-�;O}�g��uv��q:)�RI�N{egŉb©�nt��eE����U�Q�
��k2p���3�4��2��Ҕ�^e�s(�����;�EY��ô�+m���2t���BE�1��C�?9�@�qkf�k�0V�ċA�J��R�)En "�"�C褏�<�4�� ��L���7����`_j>Ν��<�$n���nl��~_Zz�a�Oa]Xp`Uτ�R,'�t"��v_���K��sJe���+�.RKF�&�yE!�py f^_y����Y~%�fZ�ôa)��A?x�����ҍ�1 �Sm12e��tH��� ^��L�����P�^~"��؂{��:��A$0�{�F�3�3�Kw�O���b��CS����n���U.Q=_k�$�� W5��V�h��J�A�PZ��X�uu2����&����f��9��H,�8�)�c�!bA�\+����Ou#4N��K���U�#^�B/��>�0�K��A�N������\h�F//<�ro�Ԧ`��8�`_Q�	�l�_��c���&��l�8'I���N4d0uA{H%*�B�����{l���sH��1���Gi�T�E��̽� �ohw�����'�����r���W�э���̾��MfMn�~1!|��M!��B�o�u���hׄl��5� *4�|��n�H�}���)�� ��r{�T���RU�}&:pZ��7c!�/�)�Ǧ>�����\���rjܦ�I��J�Y�]����J"�y|�|0��'�0�?�j��,��a;ޯ���w��]�Vi)[-yy�
��c�.9��'{�����ލ*�.�CY�<H8�y�[�O�_]Xv���A�8� ���3NT8�zO�� h��9���>�	����/7�TY�� n� �?�#쫭N����O_��hqV�CǬ;�B.ؒmc�ʽs��,gՀ�v�ҀW�@�n����h5Yf��,M!�v;ZN\��!��+��>|�7@D�.��l�/��	���M*T����n���S���t�zT���D$��A��7���D�RU�"{�١�ɋ�}���'���NȲ�)M9m4ۂPd>�
L�0�F׺=}�w� �Hc8�`�rR�yC�	z��b��`�����1�.�X�$�?԰ f|>ҷ��N�P�Zi�lw��gJ�v�i/Ő�;׆_�cN������yu*�}��X��ވ�vE>ay��K������<�;�`�aP��E��̴��v/Ѷ�(;L=;�x{�d_�u���Y��Uj.H��4{���7".�6��ϩm��n+FR' ��.F6���*'�0�˂�2T��k.t�[�z8|�M����R;�s_�H-_�F��h��2$C��\�^�Z-�b��֥0e�Ei�\��)aA�"���
�ur��aA��	��;BF���g�G�4�/9��+˄'�R�t	�U����c8�MS�k |�)�m�����(�ru@��񣴲����/o��<�ч�EhF�`VZ�{Ql�U��̗��rG��t������A�g ���S!-��B6�xzT`8�I�70��I/��x�	ƴ���icn��kbǱD)(��O L0�X���N�U��ةJ�������/&1jL=䀄����}3�}y���M���_ցe����ۄ@�����
A�5��vC�䘄 {[�p�N�Õ[&�ˠ\�3���v�;Y-Oa�p�(K�&>B06����&ܲ�\w�DLs*�,��X�g &7O ����J��s^��HHX��=J��y��vZښf�X����MJSgz�AL�4&���e����2��/���Q��� ��Q"�AC=�ń�o����
H��^`��;4�]��8@z��M'V�x{�9���d��%�	�����x��g`�'f�_����|=1;���D�ҿa1"�R��𑆚��j�s�o�:�]�0���*����=��yo4�ň���dX��DCG�Y������������W}w��G��_.73�O�y��\89	**J'a��5їe#`�8`|��M54��D%��$�_pا�
<��տF�=�lo��:80S��*��4\�a��ڷ�S���������D�B��,���<oK��_�@��DN�ѐy=}i���|Ĩ�����6_���?m���X����c�@��Z�(��C�l���=N�!�2�Ib�������Xdp[ն�l� ���G��M�����*	$�?���?���Ae�3]�SCʕ���B�S[dN� �7�y�?TBH�1����W��}?�(�a[�i��ηūc�{!9Y�0}�`;YH��+�CI��o��K+q͊隞+��	|�}���|4Q ݑ��NBk�3)��q��-kCF4�J�t<�6S�	v�74��	����&�]��� �/�t�X����%p_-%|̺d֜��$�vs�������T��Ш�$ �hk�ũ���{r�Ed���K�ѷ΄*���v���B�k�L�b����-1r�]- �{x����G�'=�Ve���,�u�����w����Nyh��0.�z݈_�z.����@����}?�\�U����2.k��__�*���gO�]9��FC�"ٽ����T�k<���0<�~lO��> �9�7Ap�p��e5�?Nؐ�\Hs[�l5><7���~W&���Q��m�4�4/ރ��'B��Ro��M��$K{����5S黲}ˈa�`f;R����̦xf`��0L�/ �xc�G�o�!�U�~���R�q��܄oڈ{[�l�('W��N?��~G�����b'�%��H�;��z_��l�Tsrҳ���h��Y���SZ̜#x�)��q�8|Oa[,�c�kL/`�}����($	S��G`� B��
C�
R��(F�y|;����\���k>0N���w��fN¨7�`\²�QH���u���L�m�Y%|�O2�#qR�e6��y�-Tl�6��1Fe�~a,��5�s��%B��ʒ��T?a�ᘭJB7�W�����3dpB;^d��ӏC{��-~��{�1r@�M8�^؍���e��Hd>_KNY<!���sg��G"((I�`�Ck�S�f�ܡp����6�'P�o�A7���{<in2bg��l���=�w5��&W��Y4f�� ����0�"�3�1b)�򮷼>m��=��Î��Y��;����FF�����ӆ��Z�Q�.<�P,��*D��y��~����R�`��̲�B��.��=�	O��όץ�����9�+L��X��r�&J�m�f��)�L_�xrj���U$�;� ��ʫ����r��F�}N$9I��<��h3k��y�S�=?�6��vM�ہ�#�?�I��хႍ�1{I��J���'z~�V��������^��B�����-��A�/ ��>�.�)*�R-E��4��#�6��w9�O'��o�cےG�$�O�L}�bQoI�=n��Tҕv���|��<a8{]T4p��#ΊRK*�y��~��J7+�Ʃod�V��N�Q�޺������WE=##�J���9Y��Am��9�_��!����I��z����k�ID~�����˸���7�M�p�o�WV!T���P�����Zى	$�g�?�c	h>���w{��: �N�����
k���$��'�������Q�� \A@F�	͉8ADis��<��R���苅a=��Pv)�g��p��Z9�<>/ڛ= PfYB9��O�j��LW'�܊��&��Mm�+�4q����~4/�M��oy플R�x��������r���E/0����{�:t�>ҭx��U�����w�ɲC2~�v,gE^�x)v�?�TEG�*���Ĺ���J��쀦����A����Z�� _��v�ϓ�Wmk��1�����2M�$W�M�<Xģc�-D��n��J}��~���J���f%���O0����."bMo�Ow��gG]�n�m����ChKR�b�[*���6�;�9��P���0dܘ�[���SS琐�,�'��#MfT�ל6�Uz^�6G� �X�v!ke����췹px���\�L�|�a�Bm��A��Y':{��9�@��b�`��^f��F��ҙX̀g�M�-clm ��=����9'%O޹vY��ح�i��'%`m��L=.vͻ2��F��&����X��P�.��m�*u��Ffk�&Ciy��c�*�� �_7��؉n��h�k���Q���t�|���=]e�0I�sp_��D�3�����43Y��R�XU*Hf]�(�RvǤ�҈H\�m���p��Ḙ���%�=FxJ�Ui���H��.D5]���mAzq�6�ª$=�N3����sA�8���G�B�4\6�z�T�N�A�AN��q�WV#x��9kC^�K��H�s�M3�7a�2g��1��=	뫳�R��7�Ɇ��n�(ꈕ�E����{�g�7����y�F��L=�v��Mqe�N9G:�_j.Ԧ�R�M¾��wU3�$��q4�b�.���	b%(�R4��/:���Sj��8.#�d�X���U.��r�Ώ���x`��~� ���$����^��B	���kv��A;�S��[��w�@BE�" ��Q�S�9u��Z}�*��͇e�V� D9��G�FqD>n��I�h�Pe���_p�Ù�D*��lo{�7#>ż��<�r�����G�Z��r�ｂ�2p52~��H��uq)���Z�3N����''p���v�10���>�t�i���C������e!I�4��\I�G�sv�j-��C�Q�_WS'��?������8
}"8ˠYn�ޣ=J�A,�;��XS�c�O�nH�P��ws��q�ha��VeͰWɘ1����l��,j�d7>��(���>�&c$�bBf�B��J����/��X|��
�N7,�UXxc�6���sW�SC��'�<����-:.�;�Æ��!���_v�H�M�=B��|�"����ymR;���X��_1�kN�������C�uE�{�XC�B$�G9�ncD4�`�?�%K��wk�߁�f����\n:r������r�d�-=0�z_�Ը	���s �
kz���8�kb�H��P�(V��yc��V��*<	��f��g�0@�?�O�}6\�Xr�<zU�݋�����Ƿ�E�{/S�K��|������-��]t�h��݇4��_�f��x5���a�&ag����Y<�mKѐ������[���,��n�<�M�X��
Ѻb3��S?!�N��ְ�>{8�v��o�6�U2/�&2�Bk-���>�\�u�I=Zlܡf=�^za�rc���XL�3�M��!t!�wg�w����LwcΔ��F�8��?h�-m���y0au[�������NT��Cp�����Yˤh{������6{ʑ�b��W��88BBY�
�7(aoa�ס��0�u��`���ؐ*��_b�?�+%�����׍��`ʎ%��-b�K��G��`����R���D��4(B�- 3@y����;�/�}Gt�
�Zj*Y��|�g��*�X>�4�WvI�ף�$�P�h~şvF%\�@�T���*s�p�e�@:E6������E6_��Zt��O��>��d�lE(�F� a�\�V�%F����\)z'��ۓ�*;:�G��kJ]�����u� j:@�v������jS�̨�je�I�.�0�E�j�'�,�zS�Y�UC�aE��C��X���m6m�b�&OP��&���ۉ^��n{��;�DA�c[�j񕰸˯�f���Ձ���Q�����I���b-�rsLy����Ө���Lx� ��/�&&��.Ѝӥ�0�kbݰ����e���n�đ{��S�_�|Y���}���t�IU���I�d8R�.j���-��J��[��Ή�YJxf;����v3+8���d�cU>���v6���y`��Z��y7J%�
Z�(��w}L(�Y'�t���\$K8;��F����"{���ծ`�Y¾����ӣ�����Ŧ"Q�v �}�?�D8�TBд)yXE����'��8��ިg�]@��?�m���˜����R�_e\|詎�S���q�@M������7���N�(��J	���\��nC�~�����0b���+�|�J�8�2�0d?�j�e$�'�u<��"�C�`����rhgNŠ�R�a�d:�#`f��o,�$�������������X���č_��V�����I�K�%X�����e���E���׵?'� 5N#<;m�7��M��l�Vp�R1�
�X0�LaVs�B�qC�rDp�h?҂�n����O�|��̬�r|�^J^�������s-{}�S_~�s|Eј��޼�#��4OX�,��4�H����E��@~Q���I
�g���:S-��-Kil̀ڡ�В���'Wt����K<�5�Q�[����3��7�M5�}���u!/p_�4��p��L�b3JL�kly�]Re��#�)�8M��p�8�;�MOn�r��Ţ�����h���R�&}�R��i��߶;�v_U�5ؔ)�*�.ʳ�_�����d�|]�}���%}��z�-.���<d;?��bA93����\�H��H��
����t�a��A<��;��{��2{������C6#p;�&��b���!ˣ$���U ��H��5ٛ�1 �N�l��ZL���TfDSH����F���:�(dY�-�C�)f&�+)�'���k��+����&����{�k����mEf_�2i9ۯ�q�"����-6��H��ȬN���P��W��?�W�˒�'��/���!��)��YV��Nr�̉G)QS����ͮA���M�}�-��'6iT�l��$c�΂=jmL}��H�i
��+��wa�b�����b�P
�E�S��)�6� LBv�߁y�����ʂl��Z�T�`��\#�uo����{٩�A�'w�R��ȑ�J�w+u�S��Q�Y��s�ϵ�S�7��G~��3ꨯ)���1A.w~q{k��0ђ�D���6qu�/B���'QiG��3Ӂ[��[�v�d�b�K!\=����D�I"P˂����b"�c�ދN��V�)rSW���0�(ȁD'K���isb�^M�����b�h"7��̆�d�I��9�n��yzm-��R9䶛e���*��뤷b�=Z�?	�u?@	 Ξc��F"�5�M7a\}}��fY�|�k���b��O)���52,���'��v^�R�qO�!s��m^َ�V�AFNWh�>]{B�֜25Kr��ö�w�	�<Ԫ<8�Je�&yb#vyu���2�ޓ�+��q��=��L�P�����$�V���O�!��	K������u�H{/*۷�X�{�uk�|���ъ� ���G>Rԯ穟n��2��F�P3!���{M9�jt��<�<�z�����>�&�riV'7��r�
\)'jQ����0��
h�a����D�:@�.!jsh��_�A��#�x.9L��B�����!Q�|y�y��\�A�e����Z>)�`I�����	M�����	d�n�e���d2@�5VhPE�����J@��T%{���%չP�+�	�$����		]7���n�������]���r��͐x�VCB��rg�o��TG����^�"����.�;��US�a�]�}h��(1�zt�����u]�莴G�HƱA2���L����a�g�PT����o(�)s�Y�~~�X0�����ɷ-�4m�z̓-����"�#���_�I qI��|ӭ��ک��J0y�l��o�6�o:������%�$��R;8�00�#�>���>xҡ;�=�r��������մ�{�7O&�����D[�RN����F�!J\�d�j���㔠^�Q�wm�F�����y-x�@0���P�_�m�u�v�D��R�	�&=sρ'w|9��� \�A��yº6��e�]"��f�F��[5��ΰ���ף}Z��s,��S�ǈ��(��՘���m˻4�M¹%�(� �Rj��ȹʬ>>�x%A�>J6��xc*bi�mI$�pM*Ԩ~���άs8Qe�߻-��d�(.�е�ZG��`D� Oާ���Q�W�T���d kT�"����$���՛t*�g���n���}��͸S&�)κ�}���LBDv9!��'W껬�^��s��(�%⢟�
X������6����K����݇�؍�CZ��fzN������w�;B�C�D��2,�f.q�L�o���Ұh���m�Cjy�d�\���S�0a�ǈ�M��8�D0�H�O,b�I#}�@6�BO}�B-�3�S�4g��뭦�\�'s"A2	M3��1�Y�fқ��x{;8�jZ���z���g�z'y����e���V��i���T��]{�dg��f�0���K�b�a8��fL����Ën}g�Yl��#VAD&���O{eYI�?iW�p�1c���H�k��&UVZ�P?��F �n��I��?�4�-g\DXz��W���m�Z������Յ�u;T��L�+���ʦ�4���g��өB����$��q��O?��3�����4�C�q��*���x�0���~���m�5�Љ_c���EVr(%N�C=��d��5����,l�g�|8��o��3H��N_��_{
|as$�h���(��}D��WWG⤄$f�aj��d��̢Ka5���K��o���*cy�
�Q�8)�.!=�m���B4��ۄ��뻧lGؽ���}uZ��#�m��̥��??#˖	���,�u�T����zN����.��ș������Z���S�[ܶ&5íXټcW�<yajP�"�~�}���u����g-{��D�ފ�]�v�`��d�oa�o����-���,B$�ӡ�n~��\鼡Ԥ��7�#3G�.����i�-�_>x�&�U�Ʃe����N�)���4��-V���̯k�.�.�Wj�-.Z�V$s���"���>��}ܖ�E(���U%�XB��ӈ�O�!qVR�$H�|4�m��/W8�+�<��|]�
��86�v#3��E��ː������7nm&
���l}̹D()��Y�z�"�C�=���p�P���\)�Q�5�d�O�ArR �Z�+歎���D]�6�q�ͥ4���3������XB�z��7�(����e�x^�X��_O�D�z*�����?��VZ, ^l�r\A��+9���6�%��l���@�"��t+�Z�Z�20��J*%0���<�cnF����e�Iqя�N�/�-����݈��NV���g���b�F��:_d{p��I�i�$��I\� ������*���RO<�є"����Y������&{i�
�6J�Do�1s�E�F��� Q~>�� K(�x0�Z��3�H$#j�u+O��%�z�U�\D%;��-'���O�Z�S���+�03�n{[��yYD�è���N��;��C���=�ͱهe�]�2�Ilszs�å��q���+�'���*�K��>��#f���s�w�3B�IN�����=����+0���l��>�}c�Ɣ�����^Bq�q&��s��Y�#���!�Q z�e&ɴlz
ݐ�X�t�w��UZ?���E�$%��ןu��5���">��7 ��#�I�����g�+���+Z�h�n8�e �D\�%�=��WAȑ��?���l����*�aR&$��gr����I,���rո���F����IF�d�983���ӥ} ^���ɲ�����S,> ����~��ݺ3m�`خ(^�9<*KY�-Vƨ�����uN't�\-��?Lu9�w�G-ļ��U�FRk�n��7��`�2�0륨�s�{�$��*p�U6���2���r��/4zc�G��/ļ��&p?�w=�|�Qu��
2�5`V���V: ������<�S�lC.M�&HE�s�]]41�4�jF�wG����"�� "��0{�����Mv���D����i ��7�6�-
�TU�2|�]v��6��h��^���o_��G����L��XK4���»��:7`^�`�n��L�dc|pJ>\���?����!�����ѯ���e^���9�S�ԙM�]9�q��y��>�0M�fƆ�m�k��K7�9[P�Cq{P�$=��B5��ő��:�G��$1'��iA��e�Sq"���]�R������+�\$P}���{��6\�	�D�ԡb�z�*C&�^�)���]+C�WJ���u�h��ۛ�V��	3ZGr&�%����F�\I*X�c^&��A|�x�;��ʝ��L��i��M�5�C)}6��8�� x\�zv<Arg�A霺�aX��d<��	y��2�
���q`STpXJ�����z�<$���Y�E�S�vi�+���|�SeG�5.=uE�i��R�V�Et�@ig��ij�B��3� �Z��,�G3d�I�Ǐ`6*�[�]��X,O�T�T�nM�6.��b7����O�͕f�l�vV0��K��i�a$���D��D�f�wt����;���u4�=���Qp-�p��pn����.;�n5.��JV���r��]�m^�g�y�D'y@bx!M^�t��	]� �^ϴH��9ݩ�L���%R���U꘥['R�N�C�q�M��3s�cj����7���F��FۊrR���;4DM������-�y����2͢:����W�ȷR��R�syB�6mʎL��Y"�,�sfA@��7B�CW���&ێ�J�Ѣ��+�llZ����[�KH�]4����e��7�tl\o��X�fi}[,�Azꀚg��i�)z]7�}?�s;IK@��8���Fy[G� ��˺��:N�������a$���\�㳪ܞ���h�>
'loQ?�
���W�T�P�����I��A=�,���և;V��<��Z�1��U�V�5��"����:W�?*o���+�i�Ú�j�d����ϊ_\�kl2�=yb�DX�߱o~[.��*OA|4�o�uQ�0��V�3��} �Ut�����&��%��8.Մޖ.����?.�J9��9���,̑,�3����*���Ɠ3��G�	}'�ީ����Nr}?�a�
�-���
"(S�
 (���h����	���b��:��:\��V�w�����`#b�l�����m����G���U�4H��ܩVT4�H�B֩v�K�fV��Ɩ|�^��xX5��bb,kc��A^�m\�-e�]ى"
��$1]�3?���~�2��M(l�v�P� MWY��V�=#�$���L�K��m�@�"�@��@�3��YB�\�pV _c����$��ȳ�EzAtJ���eHi*bl����`��,����oAB0F	k��-N�׬���#ׁ�����l��kR`^tL�#4ͭ���7�g�hR��/�!��h`K�ɐ�'>�bٮ���Y*AH���f�&t9� �>$!EPg�ܪ@��J!�S=E�,ݨ��K�g�'����}IJ�6��:*��-�{�º ��XtT[3�����#:�A�Ӥ�����X'�o W�j���n�b&���^9�6b�i
������jW�����O�7�#v���̵6�.���@]���~c���@|I*Ķ�أAPx����e������{M��£<v��_5�CZ#:g��Xf ��qC��x�������u��SLA��J�o���U1����SS�i�v�����4<3i��{&�����|.r�ōX��3H-�pS�>���ݨV#��Lɴ�@Sx�P@տ���)�Ec�o|�&~�K�b��ޒ
i�
ȃL���j����4��,��k�)XJFky����_!Q�%=��s�m�\�Yg��:
+.�Z���_	�Lh���ܮ�9����/S��O�f��Ğ�����R�'�hP��H�@�sB��#�^����X�c���4P���=w�(¹
��ݬMA��[b�i�V��9��ʬɸlP˛R�����3pteY��fF�bz�%\���G؊y�ڱc��ӭ�d����aNɽ�Q�1���A@ԕ�|���GER��a��߉WV׵{w����x]9+~�o��a�\�O"%�j'���+bc�&�<���`�/U��hJ��B~)n�����R�DB|pp���i���W7�=:D��b�V<V�}�3Z�+�*6�y�+EMej4�d#��l+`7sKÍ��j)�t����!��2- ��H��+��NWB��t0���D�RK��e�����]D5� 9�J����!�G��{�y	�h��a�W"у��z�}	���N�hnbC�dL����ph��:pI��QS<M���Z�����z�$��A��z*�~Q�WwB<�����ە����^��e�O9�l�+�8-�{�k��sr�sY嗬��k�������c�
s-a�K�'+F��6=ϝ��z��NY���j���B�4	 �Q�/kh��0'R1Q�7�o�����3��P�<�뷈�o��@8��x���c
�I���@8��ޒf
���da���@m�'��m�	ǃ�A~A�Ңd5?�yow�� Z�.u�O�@�#���O��b���	Wm�r��Ђ�����2��BM��q`5�bx@����Ū^��'��	��YE�s�����u��m�cв�
�o�(�j<F��)W2N��=��ԗˑ��=�����j�"�[��R�<�+gm܏`���Ny���XO�$� �!}e�zs?[�����å���
���#9�^��5gH(+��E�X< d�$�q�ŗ�e�Q�H�)O���Znč�3�R+��9e��Ȅ.k��{Wl/��A��2JԚ��ێ$"�.vo�j{rKA|M�`�\ݥ����z�rP)�痸W������l�D���~�����`aa���h�iL}�����E��+���7�[F��K�����e�u<5�ˆ�����[�EY���k�y[�_��]���n��}�6�3AfYh@˟Y*�αGbj��,��DG����m��"����Զ�|H���]��TM_d�w�����(�EmNE�]���_\�D�D�8)�eh@e��P�R��[S�e�@lQL��!���;=K����PM�\8٨����V�R�	��׮�@��*]���ny�
���c��C�$Z9�E��;�-8,Y�&9���*K��v�E��jB�H�<�v����i_Հw5�~�ޏ�A��;:��3 k�����M����Xu���j1��$��|�T�o���)H�Ӭ�8�6�xm�/Cьz�ܲ���G�8�ؿ�g�n\޳ �S�uX��HKj�ҁ4����/���:�YO����C�m�7�<g�m�ĭ�+1�P7D:>�o2��ʹ=$�./p��`�=�e�� ��X��AC�V2 ���QN�gF�Y2i�=�iI^Nr�9�I��|��?�s `jʞ	�hHV���}��R��0�8� �2�Q�z�Q�Ou�I���jt۔��:]�{1ӀB�b��r�1i'���o�Z��d1����`��x{��S�*��w��)��M&����D�`9�Zw�C��m/���҈I��!!J]�G1cf�磻�����MTVnE�KC.��^V�Pj�9U;F!Gڽ�_��={#�	�0�*Ĺ&���M+ʴ�g.a �DP�����ٗ1��>M��
�  �Sx�V?i\Vp���H�`�������{p<�g�L�����u߂s-���@j"׬��kA�pa+�~��i����F*ϒjT]��W-'�
���_)�B���)3�{+���"�����1d�rd�Xa����5����E2�4 ��"쑦��%���w��v'P,�f��:�lD��%�n,@��-3�6,״0AN+�C��6�"�_K{Ji1�+��#�%���9���7�=SP���.(FR�'\��0��J�潱�V��Z-���%h+���L-x9��*�����인%����/�ڨem
<�>�x��_���9H}{�����CT`�I�,: Ҧ������wl�
��W�,��5%Ll�#E�P�|,��+ y���� �|u5S��t@_W���D�/�+x��2n�4�ɐ��'�̠����͜���AcY��_ m��z>�b��}����~x�I���ɅR�8�]ެN�]��������8�8�}C�=������{040��~���rh"tK@)zw��hL_2K�g�zˏ���cR#6d��vB:�_�&p��B
�+S8����`����:�*_���������q��u��~�آE;���W�3�1��Ѳ(f�K6��Ԁo�}�R��>(��]n	�Iŕ�)���$3�5W��R��z�{p��̈́�%�7�Z����C�z+��R��N%E���&a p��M�U�%��4�R�WE3G}��*����;^���۶����m�����83��>�S�-4�2⻟���@���c�Ǧ
�(��"��@OCd!��\a�0�����(���Y6�v:�����餸�P<ǆLun������ڌ\y��'uP��@F}���	㩳���|:ן�{�!�C� Iw��d�)��	d����ܧ��s��{4̼���|�bD�t�e��q,nd�S]k�8_�2]���ke.��+a�*�Z�x��͡�7^imǸY@��Ps*v�r���� d)�|Q�>X�����
#�HI��I0�ŕ09r��~���H��K���qQ�J48�S��獫Ʊz56)�5ͪ��|n��4?<Ԏ�����U%O���N�-H�4��嗡��1���J��jTǏ�2ic�����e�Ԉw���nl���G7���^�����BR���WG'
p�}9%M8��X��e��_��3ި��$b�t(����ƫR�Ζ�:�>�d�2Ln]�Uب*�D���zƨ@�Jd*q�W[Q���k�Ar�k���6�+�~���g}XG����7�v�[���3o	˄������2�#^���5.?A��"�%?)�w,���?���$0�R��@�7s���P�@���zo�m�H�m� �#��d���nU8��?��=[��AW�M��y؃9+���ƶ������i��x�|��<J��7s�u�Y��&��w:��yf8{���8�S�b�l�����Z�K�qN��)g^�y��}����H�m��\K��3#C�O�_��M ��:d_�3g��o��M�E�c8����7l4�H>�ݼ֓B���y�!�\Ƨ9���a��M>�Ϸ-��=�mR9�Y���7�s�k�Y�W�U-���ŧ<�|��W�節C޾���T��r��%+/R�7���8gC47B8����2�D���"�U�v%`�V2��j$��7��QѰ8�-��	r��u�	�6A�QL4r�Q~��� ~q����^�aF�*�2��ƥ�����K�}{؂�ō��-孥�%�뎌[Fu�fr7Њ��"��
)1�D&�M5�F����.y:�g�n3�#>.(|�[��`����y�6���Kb�r0}7������ox^�E���L��U�5^l}��u���Q{�,�s��!�IM���f��k�71�U]�����Ė�@�W��F�a��^�Z��w� �GJ��W���(%���71�#έ�B�����CHLb�"9�tWq�uQE��{�<��# �}�q���s�L�� Xq8F�3�I��X�$8ބ:��|�r@�i�����o`�o��x��df�2�﫶Y��H�VZp�;��F4mB壽?�Z�[�i����tV���w9����lc���1J�,^ sڇ�/�c>�_��)X���l"��F�0�����t�*�üD:,� �ɮR�1�����}�z�Qѱ�#,����eC���6���yy�E��~�h" ��W��^��Rלr��5z�3&�{cWSp:�-����I���.1<Ryqe�l�|Q^ �t���|���j����p��wbeqAb'Zko:? �pT�>oBy��ផv;ch��r��E�!�ԒT��q^��6Ykx�n�c;��<�SN�
d	ւ��"��d��{�fw7�$W�# U)��0������J�ո���
U���;۳��#�^4z8�E��,�����~�αr��d�e�!�ëR4�x?�; k�����j{���;9S&��KZ��`3��S<�A�J�� #�x�Cr<g��K�1�,�)!w��{����,�7S??�
kkOb��(	��	��Xmk�/ļ�(��m$ժt���h4t	��;솗��Τ.W�O8D��&�s�t��:ꂁnĺ��8
+5(�q�y,�v����'�2�uvCsR;m�ё��&ߛS������qL[b�<:�YV3��tF��NQ��/
��Q���ҿgӏJ�hT}�pe�M�_i�k��B̻Bd���ܠ()_nϤҼ�=~~fZ��!>UU&�ׁڈ��{��"���6�ߘ�X����qI�=�	K�}����&���z2����b\�e[�˨P��X�(�,�ci���w�����8a�;io���p���Z|�UH���$�~��׷���k?ZC
�����C:��(�+�q��l�9ɚM�����MO�9��F���(N�'J���;wl,˒;�t�E�2���4�wi��L�T�Tc�XLJ��#X�k8F1&	�@ܟG��s{�
k��@�sjI5<����զU��AX�u[�@����bU�Op�@�(��E�;?�pO�/��Ӟy�)�o�R�' �I&)����o]��
�[	q�"Ԯ�[���c�r]�>�����V� �b������_Э��g���Y��P��9��ND�n�ഀ:|^f�:r�J��|Nۗ��r�:1ٴFʋg�ʟ��3�\;+�DZT\��ψN�:�[�i�3�c�*c(� �x;��n��φ��L��q�����1���+W��amY���>"	i`W��th�86<��M��L���t�|�U�X�mD)��QF��Ǣ��[��
n�� |5٤�Pu�M@Q���1�������ߕ�(<Z�y���K�a{}Cbs��e�p��	�F�hG� U�
%@~t�1�_���(�1��	��Ť�Jʹ�5zQ�Liέ����=1�X`L�����lY��Q��O�S
Q@���m���Z����My��)�~�Y4K�9\��Q�X�2������l:-!��_Q8��=|$��[���0��)m�V%����H�}|��8��m��߁��2`+�}g��cԫ6�KLyT��q�o��v��e�W_(?��e�	����C���,1�P��+� (Uy�/��g}�O�Wྀ��9TN�ނ��`MLN�y�$^�����<[yio�| �䐳Yc�D�~�f1��)9�4+ g��3Q��%�&/^9sf��w깠��˽K� ��@��LF.��/�{�7��X�a[B�/UrT-#o&!����x���>��MI�Im�6��WK��� �}V'��cc��?�����o[ڥ:�����!'�Zv]���#Kr�̓�+k	�*�]Lj�,��Z�&�#IS�U������^���Q7/��I��Ck#L:s3{FO�B���[�*�����`@�x��n��X�lΜ�/��"�N�>pj��r:k�If��H�4�@��+�qrܸ�����#L���4~�tV��eI��M��0���[ t�X��/^l��������g�!�܆��}]�8��q���2j!F��)��US�����8 W/��:�3]斘��o�8���r�� L���nti��"qK7���M�^Q�wAQ�ؘ`�sV[�M�l�ޅ���O굏נ�/�H�u�h�rL ���aWz��:^(��
�5rԻ}j}��}�ͫ7��4��r��u����1	�L"H* ���!�sh���h5T7���l����(�D��Hm��'r��kf$'�A��hG�8ʬcuvF#��N5y��l�;��X��E��|@9���(�u��WaP�T���r����t�M��N'Ĩ�4���vs�M;hA�t��8xs�ٜe�V������}oi3�	����D���s�y���w�+���ZZ�F��C��������L Xx�A_����B��4��n0��I5�.��o=�k	�i�;��~�B��_j�@�rn5{������"rF�l3���N��`Cv����j3�T�4D�z�:�#��#`�E2r]�-�CD�¨3�0W�	(����r�A�,�f�[-�.qŚ����v�w2J}��}����W��:$MC�yƐ�X�=aL�H:�hm���IGcs�{��p���Nh;r)L(^��D����b�,��Ҫ��2��lQb����e�/!�O(id+i���.r�_�F�sLT.�<E�˾^��!w>U�Z�b9�O-�d�΢2��v�AG�q�g�<*\C��B``��x�Tǀ��	�v��PA=Ī��^(��Xz�e�ғ���A��������R�Ѱ��M�NL�ÊK��Y�	7TI}�݄��~�F1A{�#5F�j���n���,� GQ�����!�$c���M����~^��>�������1���������/�_���Rq$_��@}2z�K0OxR`����/BG4�a�
5��Z�3՘U������ҙn�g�W���@V������Z;�6�N�}��G����B�� �U^�7�K�';cN���iI�LE�[�k��R���}1W���j4�!��s5��K�a�L��|�)��9���׬���8��<
%�����>Y�pC�wr�rc!��_�$�'�fT�s�OG��F�H���_�:5A�n�p���?`Y��vJ�L�R>w�^"��ܫ������hr��gQe}ۤ�L��R��>��g�a���F��4w�
S_���~�ܗ�������	�-�?ÁD-�a+8��Z�L�ҟYf�`0�<p}.1IR�JYI��Ձ�StL�!�®�i���+��/�M������>(d��I�9�&ěNb��A�P�^��c��,m��:���P:F�EFx3Dg7X/ge*son7���S���3��[�=^��e>����9�}�2�k�U;?)�����
�g��ɶ�e
W̸
m�S��nd3D"���ɾrټ�T�`��0��X�<E|�f�)�E�T8�u���9�Bxf�n��VяJ�{��#߾����M�_-4 ��)^"�qb����l�_EpUo��K�E1I�����$�ta��U�n2a��������e�j|��K�@�hĻ8��x���FAN�(R�Ǒ{-���K�tq��� E(�%I{Q
n[�j����[J�=k'$E��k ��KʛN�O鸖�~	!��&��8��F��/�L��!�:w�^����3��z��9C�ohh�$���]1��7�Yz�s�mN�L���{J���d0]Z5��D�\�j�iW? �J���7y��P��>K��k�<3q�R�����֭E�	����;O�A	���pk�``�p����ҵT���}6T�e�V�vS��B��� ۣM�m�R�����y�c����J	�"�3#5�[$h�Y��7��2d�AՓ���'��M�3}u���R�7��Ԕ��,~��䆞���b+�+�Jk���߮套����&BE_sMl�>��N�h����[f�L�g�R�<�h{�փc������p/�#)���l�)�W���zY���w����~J�1aIV	�M�n��[�ң�y�ek���-eX��J�I)_p�c��A+��5�g�1x�qh��X�K�0#�Q���ֳ�s��v����E�;�읝��lz��j�D�8P/��S����s�z��̬X��%�}ٽ,�B v��	�E��cNIzټE�X5MM��T9���"Z�h�S%�t��<�`v�$�����_IZ�;GU��ћ��3���C5@U$���4'?Ў�DW�2z�ܜ�_�H{ߓޞ�~��1;]�J<�ɵ1�e����M��WAR>⹢|4�Ձd�;� ��L���;�]�! ZJt��q����Y����bɅqR��Ż��=�c�"�qL"�1iy����[�R@C��-��]o�@�r�<Ӑ��u/9�~�ʵͩ�7a�T7e�a������l��KW-�@�|Z⣧���c����Azc���w�	#{׸��k"?�xe�a�A���J%z�n�T,�\B��	=�V+��Z|kAs(%�Ո��<ūu���e���!�#R�xb����h2������A�R]�=`U�	�ڒ�C���b]���<0bC��=A�E�tV5�Å�+���Z�|*��rp�9�1��*H)q�b�jI(�lP�y�;!����~]q��'�Ȓ�����+���8mʤ�^�N�W+�Z����]K�/����z��ѿ��D��CMm�$��Dݘ�Ֆ�͝��r����?46�E�4�7���R=�
	��(o�ڰw�	'���22C-W��5_l~��>��]�S�dh�{�t~"��3��N��F�IKA�~W��=M����6n��dˍ� �3̜3:�^Y��X�+}�C���?:�G���<z�j|ݐl����Dw>�_�gw���?��O��l�p�]S�>�w����O+b���(q�ʏ���V*��+Vr�ɠ�������.�:z�
B	Z%��۴�>�� -�EH?��0`�Q�"�r��j���w�ϋ���{ը��bw�bs�fQ<��Va�(@$��ġ��-7wm�z�
��n��XX�?�;�)jS ~��p����'8�L�$�J̛yI�����DW�>�s�"��Tqו�$���j+P��o�T��GN%n,��4�RD��@<[� �Be� ���z�ii[yESX��w&�x��� 
;�1����(���p��|�0Q��u�O���O���������?��!��|i�3*'z���z�6���$;gol ^GR�L�.�6.��v�a�[x��,�r��<ʨ} w�:v�Ij{��3Q,�NX��J!�|�Q�x�N�>�{
Z}?�$�iNB�g�16����܅3�8�`x����j�~![/)~5��l{z%n��;D�h�Z���ӑ����G�@vjt��;��F�Z��!�&djX���Jl�1znd"�5R�3.�s4\������qѩ���h��?zJ% U.,E1H�ѝ@�T�n�$o�D&�UN�B:�$�p�ө�4�(`�6���}�
����k����_�^�߫� �޳�V��M���P��ᄥ�2��M�����4o�s���QH�ŝזk��\bC�)@�auK����i4�ЈpJ�g��^���j�3������pY|,�,L��Bq--B��~�wF��9/ހ �<������aH���nO���~]XZct��ѵP���8V��8G�q����g�O��ᅮ ��K��2��Hn����@v �Q�B@Ǎ�{_^��^e��ߝ����ݝ��AWc@^�b^}M�-qФ�|v �����k�Y�PG0�����C#��7�`X��?��R���#�p)�	*���gbV�%&*����
��o��uxB���H��KK�MYv�^I;L��T�s,����,d
x[�H�&��7}!b'��W
R`���.�/£;)�zy��q)�?�	!?Z�A7��|c�uJ�K)W�JCU�Rf�1	-��W�O����hB��s.8A*[��)U� �=�\�<�j#��H��{��_Y5��k9V<�Ĉ��C�-f�@ m�)��ek�^��_ͺN3�U�ji��b�ȸ}�كx���'H�ֆx֒�����R��X�������Z������szs�����^�c�7�5{�qc���u���	��R9j�)!N䶷˖��ʲ* �k��k���|,��!-a���tCx{Unw�W9E��a���\�b�#�fdT�;�L��ehP\�y�jS���$�!�_���L����_���Zz����� R9���ݹ��e��yh�s�9��S���Q�4�����wͬ�nז����}xZ��}R~�~7R,m���+���f�Ϙ�	�@v�P	D�J��[�x�(?11(u��u	�w�w5F�TFT��j]c0��o)�%A�{���o�F�[)�lo�����R�l%��.<�g�3��>E���w�K<���K��ݎL��S�T�k�ym��i<�j:��!���L�oQ$A�2�Q�[Xt��dS9}�����b�>����#��#Þ#�����M��Ҷ�'غ�c;�־ל�$k;����
,�۠<��a�oǃ6����"��jh����~Z|��LM�0�6��߽»G��|l��<r7v��B��#�'��v�$�Zy=�y��Т���;C�MM����^��L�e{w#�����l��-AC���d�,^x"NF�����E2�Ģ@�dء>R�c��e�	�a\o��Hس�D�����0S��;M|��΂MuL�q�2�S�vH�_��v����`��r�='�6���iXr�.�'<�hK������]�N�$���s+�� �픺4g_<�ݰڦj���w�ڋ�M_ ���I�^�����?m��R��Y��g 0k�����F }!mI&C'�Dy��Dk���[اHE�����x���L��|�yO4�,���	���>(�����w�Lڮ��S�Y��JGq�La����|�o�EQpqA�&!Ȓx�$K�� ȸ֑A����a
�\�%~�w�@���&v���: �2�[�S�����SW��C;> ����bg��9p45>�<E�XV"�Y�J�B3y�J�z���=��Q��g]F��L�N�,�@��' ʀ�6�i"�B`H���s����J"��sBF��9G��On�"4�x��E�h���6]�M�� ����k�ȇF�R�M���ϩ^����TO�>p�	ޕ��"

���I�3cf������0�����)��P�O���c����%�Iv`�X�ŕ㎸^8y:��w�=5L>�;��D�YH��Z{��sR[����;�%y��שӍ������a)P6L�\ң�C旣ǁ�N|�D�$��"Ϯ ӊ@�sn?@����یL�z�$t��CG�Y���Z�ຨ�+k�)�)b%%����Sg�PL�j�;e�������&!��`+� �����f]$M��]T�/,������Qƅ"�m�rAs1e=>Q�Ё��2/lN��O���p���-�&�;��ھ�-7��Y����� a�6��"�&؜oDjH��cޕ>tQ�b���&���mH�Kg�Lh�Qۣ%�͖��xS�A�5�̚w��g�{��t��8�՚�	��=�+)M�av&��51���qK�j{��
��%�TU*���k��"2�*+�0"��������;�
���N����<��7"k|��E8cp;�H�BF��n��pq�+?#�gt9C�1~�[�:���"r�7��3�0A��ml���B������0����2���Lw���y\�w��R~�!�<�u�b
��|X';{���)UE��-�	C�(,��u�[s@����<�Je��:���ٴ�.��c����(� ��Xd�������?�̆���0c�y�d���~��;Ǳ޲t�O�l`��]����T�O}���&d"�W2�]���4��/�T�Z�ݠ�dq�z�?:�P=�J,a tt�t�� ���QG��C8��
ߵ�u�∬��U�
PoI�Lu��$���Y�i芬���	�p!����eJm�\,�����T_����+fT��H�(�I��SF�_�/n;��tԎ��;�"M��`�G��K|_�g����-~X�cD�|��4*\%BnWmWs�.0QR�g����3etFV�苀�vY�T�����+TG�h=y��2��ϗ��'�`�~��j��1H�M(�TnjzB1�@T�eJ5�3��k T�i����p?p��1�H�]i�B ���+�О-���E�A�U�n5��i'�_�Oe��X�]����K������N;�e5�?�IR�����Xۭ�?�/Dn#6���-��^��P�ׯ�-���"��Pé��h�u߃շuN$��N��4�w �?:�s,=-��p
 �O�`N�p��pp�1���O� &:j;����'�j-��Z�y?�NE�Y��޻�Lo�Џ�<g�ƍ1=�:s�_�:��Tr4�@����_+%H �|���G&a��/�~׽��\~Vq�f�_`��~����:F}\�@e�զ-�I�1�bz�\\Lȱ�Wj��Q�14j�;Z���`����T)�3�Ή'��%��d+a��f3QQ�o��B���v]/�E�7{�ɫ���������٦�!G|m��)�1�	�_�@PB��"���l�����Vh̎~h�K,p�8�����χ�,�s�q�t�Ļ��*ʅ��Q�o)x�]��.��E�7$J���u}���=�$sc�S.l%R7ȍG�v���2��.�;�䟺�o�-�}�v�g^[�*y�]c������$��LG�k��E7k8Ͱ��V��Zy�,UX	M]O9R��v�eKAG���&���s�o6pI������K8�	"���`'�&#�=�a�o2��ٴ�Vdt#Ҝ�bU���1*�	~|D)$o��vH*0S���]�,����HVm1��W�p��Uw).nX���_ZU��I���~i���!��o�hb��oa�q�PD�|����	}���O��u���eD�@븪��`U_Ĉ\��j��J�?%�����	��ѱ�Ӭ�B���v��I&b=jdǚ���02t	��i�4���%�_L[}��Kh�e������"�Lz"�f�����;X�SA���[y��(E�K����
���3wge�_���	�F�X���w�>��1n{�r���7璕
�H�0�ᇠ77��)o�� W���.����uV��2Ӷrh��!����l]) �qg.W�t!Ä���������Jw5aK��7���!lS�&��ʼ;�t�XFB��ݪ�[Sc�s l@�]���Ξ����P5M���?��L��)B%G[�F~g'�ǍS�x��o�ǫڃB��0���,�8�����*��� ۼ^Vbp���i��KӔ�ۜO�D\����韅Iϵ+���a���	M�xnl�[�ir62�V,M��M!��1�	�8�S�5�3��mJ/H��~�zT���f��[�}!�������g������l��腣�����:�֎D��0w�@+��[ʯ��L;��p��7��k1�e27�83*c�5�$�V�����x' S���T$�! ��nIy^+��9�sq��޿����?�r��M�\*��j˕6{M�����W_t9E��ݐ�R.��86���4��O�9Π�;��y�6��e��'�A��E�j��X�ܙ�<�₁��Ra��Ϊ[�~+�g�\}N�^��JI3���������L��Ƿb�A}�q�d�];�p�6���BZ8�͌��J�n%t��9!�%u@��%՞Q�t�e�ԝ}m��;�t3=4�JY*�>������N������=�kˣ�D�#�'Li{� S�!��P������x'��5�Ռ�A�G��������;���T� Bj��Q�i����1��?�d�$�iJ~FJQ��;鞈�W���4<>�&VNv�6�mZ&��ȆF#��ᶭ YՋck���Q���-��8̢S��~�
o�[�094�ą�Kuh5�Nc;Lp�x�Cw����z騒�T$�UX�{&��1�l�h�:��k8�L
�xK�� DX��$�({o��eFæz�a��L�u9g8�Ddd����U��C����J�0���Ř�����{Xf !d���%�
 ��=KMo�;��x�ޓ�i��]���F�r�j>��6�Px׍����Ҝ*��u���3K��e�cejK�"��������{�Z��]���F+R�/A�=D�ܺط^Rp��z_�9�?�E�J~��s|�|߹/�t����ĄɊ� �(2=��~3�����T�72\���=N�{�]r/�)G���+ɔ֍jQ��t���wAnD�o)&X���)ڶ�]���Qn�`!�iC�~�c����4���#�5��{h���d�}����S�c�Mu��:C�8�����_P�������[L�zQe^~����xy�c�xx �`.����'��>EYب�2�e���u�q���7~ý����?�D[��U�d��ʙ��AIm�o]�{޼�ܟ����>�
$�,-+J=<͂%}Lt��2i8�@�Y/�᭥�/�������ͺ���ʺ�!�(�/��am�6ؼ��]� ��-��)�о�bʞ�����w/�j��a��B.D�doVK�+E�\��V��"-�˧45��UFG�t��%�o���Gg?�o����Li��L�	6QuC���xZ�|�	ؘt��Ţ[�5����,�qc�[D�~�����
�m���z�z�9k��̸�K{a.%y�����Q�����{�P&�P�5����k����I�Xع�B��"��Y�ۣ���4�=�X`�<�V1��ûpb���Ą���jh��8�:F�b7�����ٲ�Ժ׾S���B�d�\�m��~��s9x!瞆-���˳R�O���'�h�;��W��ٝ���Z��V�Q�����޺hm�F�c.rۦ$G.F2ގ4�E�#��\�<�10r=^ �p(����73�qQ���U�&$zV���Hu/l��b�7W��{�Bxoe)x�5MO�:RV��SŜ~�^�%�����ˑ��b��􍉃�
��;��zs##Z-�i�\��4��_Tl$Ev\�e��5����5�!��0�/��ńy~��p�hW�É\���|�r8�okA�=��#qK1n�p�$~@���1�8eC��b) !��U�-k(U�F�Rx�aSi;D(
��&ҿ!�Z5����� ��rTW��Kz�T�oӡ�i�ǆ�->?:����J�;���|[�g+��&i� ��n�n
�_=�C�S�ؠ�7$��u1�a� ޚ�pf�nE��zl�P���q֋��{��aU1�uC��A}�~8��H�z�F��UΚ��D�Ηj.E�(<=X@��i����|�K�X���l�o�bF2_���`2�Cn�&s���j���6Hco9����N�9B�?��Kd��6�����>}�ZI�"��q�Dj�z�S1�5��$t=H�������^34����}V+,�u߬�1�����)y��#�YԊǽ�� �����s����\=�Ǌ��q�˔�ԛQv�}�W�-�{?��S��nq��zqz���>���=-�����W����*ahVൔ�]�3L�6gq�-ޭ	���|қ'��Zwφ6�އ[��%G/��3��:����i3f��͡�<1�>	qvV�ݜ1��,$��7:�獰b�Z��L�_�$�:�}�
��>t����Sg�muJ�$��YQ���G�� |(���5͗�/e�U�|�;�x�˘mJ%mX��y�v��=�� �q��y�ON�W"wb�w�6��E�[��M���: 7+�n�I�<�Ji�õ@���Y�"�!��!�����B�|Zm^c�e�P���M��Lĭ-M~�W��T�1�����6�SN&�,��i��
�"463Ʌ��|����	?$��[���J7��3s�Z�����''�f.7�K���a���:H;�di0P�j�\뾭�HKEA��� sJ��_rՂ�&���)=Avl-6~��T���z�.Mpa����iuאn�v�QD�]]��dXJ @ov�6��K�9�y{��N�X�T,�OȚU� ���NX��� ��E����t!>����^o�X���#:�
/F�yr���Y�d����f��[o)��ϖ֭_��|�c���/_x�}�A�E��Ah�=�~7������@){9&�� ,�d-���|�;��_�L�q�y�#6e�����s[�����R�^1������Gƀ��j���q��ם\��Ր�U��H��c���<����|��=n8�b�"�K� ?��bn����V>-]��t���7�#�>�-޲:�h-Yab��?f3ZN��^���⭕����.�h�hh�U
{��磸#�a�ݴ�K�PB(q��y�����g�}�:KX�)�6`s���wB�I�f~��˻�Q�a�*��qL�j�X�8�J|�~��2|XtP<evR��I<�J8=�.v�O)<w�ϴs̊a�|m-Y8�s_�N�W��������Ǵ�[:�7/Μ@�8�@1l�:N�"v�����VD���?��Ǚ�����$�ɐ'�+Ǌ����d�Y\�"}`K�=Ь��5&=��d���z	�|kz�)�ŏ(O�YV�/�LU*�\5�4p'�o���`�-���-mJ��_�;x�NEx�*[N�d��T#��Ӥ,{~C���ҿ��N�
B��[��=��G�>e����no1�����Ņ��*y�8f�T���2��-]��J�qD[����t/��'V|}MM�g��WSI��]�2)���d�cʒ(����-�9��.V��a�!�&�z��1���S�l~��$bC$0� �}%IE�??4���(j�y�@����!��$<	fd{
�L,�6��
!4����o���M�L�^VO�GG�^�r��I�
��=��M��,<�w�mC{`o�$����X#A�&o�4O$Y��ڕ�&���"�eJ�R��o�.�Q>L��
�'��wg���`�"�3vB�N�~�I�c��x��SV�����W���_D�O0�/���4�Z�m^j?�����m�-6��)�F�C�A%U����o���3���L#�%���IM�}J�d\�kN��'�:$�?�Y���fT6�\"1n{�5]/Ǝ(��^H5;f�Z���_M�>���WM�Q���'��I�O��sD���t�Ç#s~���q�ķ�ݜO�,h��Z�bx�,!z��K����N�'.���D1��H�U��](��!?4�[�mN[/q���sں�Oo�b�����n�<�e��oÅ�(��+k������R$NL;��Iݡ7�/i)�Y_
!@���=���\�a F����#oh&(o��N����W�=��z{�?@����0�UR[S[aB�1A������GcQ'�_�'������獱��i�wrt��n���m���[�����p8`	�
����T����s�3��J��u���1ӛӔ�X	VHp�9��M?=6�bGاWp�b����]�v�(��Q�#_�P��K��*�
JHu7Z�G�Jp!�t)[_=݅��N.�4-�vwVZ1/3?Z��Km+?�N> 7f�m�&��:{��H7v!�i/�F��I�s!4o����c �{����������D��n,6� JB���� c[��q�rr��"���]HSGct���M���-T\|޸Sf��+pe]�v��*��u�)��O����0"���MqKw��e�A�/�������3��}�����3��JH���-0>,BK��Ċ˳m��dհf��EmA����M0G�@�\�	��;�ߖ��)/��� W̗�)���ibެ����=���XNn�������^11Y��`����@-�'���ƫA6��/��B?|&&��A���t�+Sp!�M���d��ܘ���&�+�xY��#���Ԇ�T_ʎ�O��@�l�B��'"�:��pH,��4\���f)%�Fz� �:F�v�xy��'Ƹ�Co��9?P)f2Z?X���z�˝���$��3Of�f����D`h�v���r��o� ���1n��׌IVak�����F�=�������
��T���n��� ���A%aW��ʋ)�y�
�GߙU�B(�C5�[�]�bc�T�GSN����
�牕d����=yZ��	2S([.U]w�&�4��OcEQ���9�č�ɵ���2�Oa�,T�O��j��θ���f�u�J���L��-G�Q�_9��HSZk����@i �PAyM�D������_cD��ʵ�7ܓ�RG�Ơi�5wl��P���jMf���߫I�+�m���R?��&��dj�F��Y�i~�*d\�+<���w���sF���>�C��MIhI�D�z<zR?������W_���(Hʴ�B�:��u�tl�'�Z靯�z��1_l�8�\&uL�T��췎��+1��FK����+�/q�L���">U��*��ҹ o��O��/��ך����J�@���,m�w�C	_�������U���$���Aâ�����꾬��[�o�2>�n��<�x���-ݑM56�ۦ�:�l[�eq�߬����Z�����X�ZOj]������qe8=@|/��G�͌g��ac�������W�?�Q������F}]�?�09p��Sҝ<�03�
OQ�V\����2<���4 ���b��Wᢓp�O�$��v�3l�
f�>��E_�~����S�:�QȆ�*�w@3����7s*��J��T�ݤ6���ɏM�{oh���˥A�����]}b��SK�Q�.L�լMf&�m��)V?=��R����KU�v�wz`��5@(�s&����{�!y��M�Tq�p%f�����f%�*�I��
��hvMՕ	��R��h����do�UQv��#���-�^m#8�U/=�,��ט��3�?A;�t7�v^5�]!l,�m6%f�)1�'U.�Q��k�i����'0�{���L��O�ǁ�VT].6�Y����H��W�;J!�@M�>�85��z��C�^���H���r�ve.��o3)��~�9L{nu�e6��$�4G���1�$6f8����h�iW�r�nV���}�Zv|7��VV�7UJ��~����Pm���Vރ�Cm�M}��X2ѭD��g�CH��.j�9���p
qea��Ky�� L f�?�a�+���)`5dw�׼y�t�B�|�N�;�_;��������"O���R~L�R�2�zOIf����m�С�*����Q~�����F�?
�mU��lu����E?m�1�푦%�R"�*�(^��\�׬3r���.�q� �эpHW*�ڤ�pd�U%#�+���t:d'}A�t�gh4$�ٙe���1�M?�����D]îjL��Чa/�c�-�*�=��Nt�jq�	��d�P	����T�~�V�g]�m�D�&���:�bG0M�����4�Z�� @������G�t�@a�'L�<�gE�@k^������P�^������M�4.<yܷ������X�3��< ؑ�\�p�������F��R
�X�x�"�zu�f����#��Fd�<	W�����;�ϯ�y�ȻI��l�$�eO�{��JD�jm"=�A�ClQ�#+³n83.��H��<>!x5*.�L.�*����)JJ>g�32/�!f!� ����O�f��O��
��[�d�^�k����[��p���9��t+RO�ܤg�[�m�j�H�	��{(�b�����ˤDSo�j�^�W������m��_H�&D  e�AXj���ם���\t����(���=EA�qH�@A*L��Y�q��"i�����������C0���|T�PQg�琪tBo�+��g�EB������Bi�yv�����	慣���GĖη)��F��f���dϻ0��H�I(�SGp��q��(�E״��H�r^�g����z����W���b�U��f��[lI�x�̧�O����~T���vv� >�D�q��$���o8�������9�������2+��Tұ񪿼�i�H�=�u�'�.
��D�O�Qk���<��IO����ˉ��D��2Q^H�@�T
�!����=�P���:Q�1�#?-t7���/��1'2���
1���Kbڦ0h�����eMȝX����8��- �t͒Jm� ��_r��~b~�'�X�M�/�:o�Ȥ"��ŗĊ+
�D&��6�^�q,h+��U�F�n��Lc�u@�q��!��Q�'����ޮ��SR\��q[��U���v4�ps�y��Bo͚٧G��B�naV@pA�PR��TL�UR`w�ø�v��X�tk��;Ǹn���$<Z]���T�cAc�:J�q-:B�� PlZs��8����B��~��>4�4�`s��e�)(N�Ț�lN�Q]��)`�Ūu�oGcy5�G	�f�}{��v��;gj����P� �(ƈ`9�y�W5��9�HK���a����]�(L��b�󊕣�e�C~0݆�x�4��j!d%��Ae�}x�%�vF.-Z2<���Ҥ�&T-?��D}ro,���>��Y�Ե�J�9{Å:��_�7�J�Nw_��&�n����,'�B��1(;3b�<흕깫QJg,6�8��.֏�w�ÉP��y��>� �cj��|�7�&_W=}V�����"֒ht�ۓ���HH;le�������X�=��?5�j�o9� ��ڦssAI�͇	re)����ײ(ፓ�@$2n�8�r�U���4=�%� R��� .��w�H��ӒH&=H�����T8h~n�?���ݡ�;ҏ���d.�Pͤ���*]���9�j��V��$Y��p"�"����H�A� �{�����̴�%e:�ࢃ�{���_�"ē�x_�ݨl�R�H�Kvܤ�Hwi��3��=�fm����#sw��XB$A,~�Ӄ��,[�c�GEg;�@:�I�4+�ネ�V��֤LeY'���t�S�-b�Or�Z]o��q�ۦ#C�W;X
���7�9䉇a���!���c��;���g��a1�"K�-~����I=4�r���c�� }�w2��X����:�M¡�#̡�m�R�X��U�����Q\����(����r��5��)���0/��5]nۖ~>쒒��Y�ŷ�ä����Mߧ�w�+���_2�F�\���3���A�Yf�ֶe�A�D�ɥ�B����@a����SZ��c��ꭇ�.}\C<!���g"~i(����2A�b����$N*Ѵ�f7߀Qh�+���56��z@ ֞�[�?�dK۹�ctѽ��ve�p�"E~�+f�a��%j�������/2���a���7��L/=oH�Wӎ��Q�sQ;2��LG[Y��U��}N�ƞ�'%�j�cN�����b����мu8�*��IC�C��� W�$eBp��q�;���({���N��'�v�y��m{�=�t� �?l�`�]ḯ����������������c���!��:#�Y�6t��}9Ԁ5u����������'��nfh.'�P1	8��҃�6jD"�ހ�ZI<\s�zs�֑�'�����/�g{�M�R�W��曊'��ȋMO0�Ϩ�.�.D̉�bf���j
g�|���B�RDl����z��A�
�=o�!h`x�:! 26��J���@�����`�S�*��0kK�s�7w�O��=wO�]ㅱSAb�V��n�Q��ĵKC�x��b� �Ġ�����`���#�R��4=W�����!hh �	��/~K`��T9c=��ր�;l%!ʄ1�O�:w���o�����ʏ���Ѽ��^#F��ƈU���꒕xOb��Fc�p��|7j�6?��)TY?����kZ^E�5�8�U�޽ޣ*1��ն�-	%�ױ��,�D႙+�e��-���]�$~.�gv6z��d[eG9�`��#��N�vNw0�V]�N$����(y�w_�&���JZ�j)�u2�!�X�k ��n��,P�j���gU�ŰTz
#$O	&o�mv�/Im�cA*v�ʸ��t�v�yB���u�VysLj���'��2 r=���(,��A}a�s��M/G��-z���Y�Vdv�WhN.��Nr�{M��.zzv���އi.}��R��9���d
�)K`��k�����J��i��Y�j�#�m�p�]�8ҹC�
,E�J�)�|}O�
�o���%��η��B�e0o���l��}�&,߯��c��o)���̈���l�[�����W
0Ґŭ4�^�(un����ʐ<":�O�mO��Z�'�@�4��H����i�.�F��ONl}�;��G�$g��,�1`�6��ܐֽ޺e�5:��պ� )�l�[�/"p�vL��	�lm�r����p�b [�}��R��:���BA��Y���d�;�`P�?�����<ț�bf����)��MGՁt���"Kk�3�d����uු�)C��aԜp>�x-kTԠG4����~������ܲ�\s[����64:�c�釆AM8Q)B�#�F�6r_�Ѻ)~ī�ӧ ���Zçz��u&���KV��� Qwt@�;ׁD���n�&M� aїh������)8�^e�1�0��R�A:�� L`(��b���UeL#~���s��w_$�$؀�tO�y��W���iB=\��}���9��f�iin��cgތ�0e	�f|1�w�2/�������s�䞐��poq�n�b�����;]RF����#�#V�y�}�#��_��D�~Ҋ�_�S4Cg��z
�$Rn�+S6�G�����6�����*���\��ն����7+���}l�V@�t ����4�k_�yV���=LS�zdDeB�Z�c`!�薽��;Uo����g20���f�<���?�x�a�=��>H3�Wګav'6���0U���y�y�y 0�7��T4��x�u���a2�Rl�a�yla|�jHŖ�6�e��3ժ�l;�^w����^#��s����e�R��6d5L�
��W+M��kZf�.�}P��)L���΂VA��,�~��Ժ��������a�BL����K�Y�y+�9<��P�e�gmM*�pT��e@UAF��a)��c�V|p�6���s�IoRj��̩K�.6S��d��pWGZ}ė�ۍ���D�G	k$�7:��T��K�lE����Mq�UG-z��_8�ͦ8����6�����d���Y���d'��!K �q�+����rE4E�{���b��^�J�0~˟�cOL����X֚�Qݧ�^\�����8��  ��i
�<�+�k�ӕ���f�o�B�=E�h���
+�,Nb�9���SZ�qp��F*��V�Ӊ���C����=��!�5�M|�ۆ˓Y.�ٵ�\��[��S$��}ˆ���4C�oX�	��1-.��n���x�>�|�^���	ʑ�>a �94G�_zz�DT��
��3a����1�~Yo0��l��W(�����U�шꃣ}[��eο�J�L�j���چ��#��v&��7���@)�G��jת��f�'�*�^k�Fd�QI��N�����c��v@p�dJ���z��N�V�Š�ݧ(.b�A.c�YݶGi 58|o���Fp�F�~��J�Y�E��t]�J�q7�LV�u=!���Bh�FEj'�B��K\+N	A"7������n��r�3./��{���je�y��WC�n2�������|s/�4�R�VM�"rr<��j갵"i���߀r+}���!�A���-�g!�Ŝq�)ag�[��_+�\��J�.	�N�T���³ �l�yt���v����� 4���P!�v�B��I?j�wo�1��db|A4r����Ĳ"~���D��rY�a�����9�\X�:W-��РK�>��l5�v4X�G�5֎�(�� kf�+�P$	�O��5��b�<mt���J����ݫ�5����K�mK��.�����*`�Fq&���M�QV��ٱ�]Qt���*O�}Ny�=j@9S� ܯ.�di �HN�""cP�;���ʾ�4�%����E�ld3���^MM�}�aHt�8���'���4ƌv�#3p�d�<{�8�S���e66��Hf�W6Y�n���ccz���l��T��[��6O�j0�9�:C�T�+pC�[�!
���a�3��0+����NH�����g��#�����g��`��֣���}�����nN&s_U�|�¤H��x�N��� uBQ�V�190@��??���8��4�Q�NveF"�ԦlRb�����b����9�g�["��\�c��}��?�Y��@O��8�ڦں�_�}�蠡�X�`��/��c���9������ܙP��-l�d�W��𯲫�d�('�Ip�Z�n�C��F"2���(��v�-��;{�xnK�:66�����1<��KOQe�J�bd�Vw�m�=�t���A���{�f��Ԍ�[m�C1y_�tE���]�i�H�r��c�t��tnfF���ZFC�$��D8x	j��V��F4S^����΄��Q�ٵ�+�~H(�+>����ԈW��$�xݜ�(R�P7#ک��Vf-��gb��	�>s�[��WN�.R�I���/��u����ǌ͖J��Z�x��.�ץ��e�cѲf{�GmF+ӍN'�Y/y�) �#v u39i�yX�$��3�e̼OwH~@@���xu�B�c8�Ա���Η�BFlg�¬l)~2��3Z���o����!�x���V�_S*78�L,�O"�c��f��-�ĥ��qRܤ��5u���e��Ox��vJ]�L��?�'���1�5�#���U��"����;�ȵ�F���#ϔ:B괚D����6�;��/�=;�]<
�s|�Rn]~�;�6���v���PC�_��(��+��B����g�>���bb�څާv�6U���Y�+��6��q�\K�9���mwP�,g����IF�A�ك}nDj�[�f�l'����L�o�$�2��Y%'��s<��Z���QW`��^
���Bj�/qZ�t�`.A;2,�:4��2��Z���� �ev5�2����T�E8�8�݂��(��6��mE*�v��9����;�-	YQo��LG�p���Uhp��|F0��ǰc�;;��S��$I�
o���C�|�V�՟* u���l�1k��3�k��C�ZZ�Xc��z���.�q�
���ld�5�z�˙J�ӝ$EK!)BkвW��V�	#�񌼸8�b,-�^�^&�L���n���`1���[�o=Cx�Q�݁��1dw�&���Ϣ����]8��eJX~q°2�����F�ELP�����<�Pѥǩ���X���[z��ih�]�Q]��Uy^\��{��L����^�3h����2��S���%Bm<���l��2/�iA�:8�V��i���� ��G��Q�)���n[�)�[6፟�\��-��R�a3�3���?d�`����qfsp�KGc�_
Es�m^�$�W�SC��yA=����<1:�ْi\_ޠ���&��.ׯ�x��;8���x.f(eo�j����ɚ,9�D� �/��δa�q�k^������@���H�)q�B�,���G��L|oe���던U�v��(*� ���Y[ ��O�M�pQ���o��=PT'����2}�I���CɑW��N��3�Əj$����û�wU 7m��/RV" �ES�JN>j��O�<�C�U��\�a�Q�V2���R�}V���W40�k�p2h˘�މd+ꏶv��gEy~ܝr��i5���jA�
�R�@�
�c�h���$.�^鬑
��pBӽX2`Jư�|���X𼓪�k�}�V�4MH�.wXϲ�W���L̆�PlY��3���hEjz�q��GH���,3����b��lu�ʘ櫷j��s�`s�/�����T�֔,�Z����������k��LS}f����ؗ��z2��1B�a�ƃ.|9�`�u�,)F�EӮ�|o�RpJ�n�Ū��'��.���f���!�a�6!�T�9�q&E9�0�Ǚ�b�id���V��kR�v���pD�I)3�_s�Jq!di�%�H�d��Ժ��m_"��E�+���d^����X��Ԟ$�>�g��>u�dN���E$�J�3����	O���Ձ�E%TÜ�V��)��%ê>�����?��]��fE�m��6�L�t�6h���+�:�����[�����I��~��J~�h��:���=��:M'���)Is�s�j�Iaz���`���Q��9�	ҘcO3�>�h!�1�+L0�Q�}�n!�ԩO@��F:�A+��¿O�	 ��F9���{�0��+C/Ч�������Q�T	ȶ��Z���@�؆�4���
w�����Z�a��n40�mgx 0�srS���@�)�$i\`��n��Y ;E�������[�d'5�$��Vʐ����}��*p?2��#�v��,�Ұ%f�A�_��H,�	��QA)'�Ý����E	[�d��X���m���Sշ�v�i�ϪCԝP��m�Z)�c��>/D���IY�Q�����I�r'f�J����5�T���-��څ��n� ݜ+*��|u)yW{eyqw8cb=s!8�,#���c����c�ԩ^��I�RK4���<��ceK�����g΅�C	��2o�;�����c��T;+�$1�mv�w����M5�O5WСHmV] �:<��ɳ����W&g�5i��|֋��FsўG�2��7~4�\�f�.�n>���I�g����*�����hV���ts|�1��}�kݑ<S���B�؎� ��"���
�C���+*0;���u� *^k܂�6�����֥b�� ��d���;�� Le�p�"�!�<P)���b�%���K%�v�-+�5� h��yx0:�<�SA�������EQ�$�}2V�i��V���-j*�A����}gJ%0��Q6rSb��8��ĵ%���3�LhB��I���,�ܵ�V-�[�,���WT!����r�Q���U*�(m��Fc�IN.���a_�<��o0z}�Edv���|@�P4|��.W���
+E)
����8�{��zgDv(��L��*�%_nf&5\��=���Ձ�D��ɜ'��	Lچ+�P�EG&��J�"6~x�1Cd���w��IN����?6�������xʧ�0�G��7�'T\+��{��K�Fn�t6�)+5fk�4�G�K0��ʕm~t��9� �i�	/(�Xy��e9�k��?E@"�\6���>����`��'hY&=Q1ZfysFq~��������`�.|"��#�L�+A��N���>`">HL1�8�t_!/�fB����KS'q�/K.�oK)F�G��M�n`�.:�Vih��Z��m�`��.x��x�W��k�;������,�&ӧ4�!����<�2�Y��ږ8���2@�(����ى �Y�1�gvb�:>	� I0�nl�x��.~23nDb�JW��An�M�-\V�F��k��>W���nA�*Fڙ ��1����$㟬J_q��a
T�_�H��WH7� ��N�w#��&��︾�3
��q3s�:VZ��Kh��� �L�L.��/)6p�+�;7+��t��lKV�����ᄚ�'[)7�$�l�Ho�u��d��O$�rZ����1Z�K��H���w�џMmE��į��Rʹah�\;¤徳M��U��M�$���'�ԙRp9��o�IqT�|V_�����N��Hl����J�+m�*��s8\-]F%��ف�01U_�u���H��V4��Ѝ3ϸ��������VQ�8!�8u�b�K�1�r���b�k���\ni��s�@b��,7w�#=���|Q�դM�� �6h.�Ԛv |Sz� ֬+`/ڿ�V�pt�e3"���lq��yiͣA�р!l��ʬ��~��z�dP�@���n�tB�R#P��D�h�
iN"�x�>�'�R�~Y2l
7��g�������y���\ٲ����2���/������<��q�B���Z�	�,�?��(X��Ia��F�m9�mX���~�G@�LT�K������&\b#v-
1@#;yFp)�ʗ�uR7(�U6Gq;��Oj�u0y�T��|l8'������M`�麃����9��