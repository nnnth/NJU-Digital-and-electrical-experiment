��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����v�c�{)
��G#�����]�*�b�~��X&й��%�֌��J���N��<1��B"L}D��+�Ci������ P�ɨ����~m�Lp2��}�Q���ɳ�\�x��n�::�gZ�d���#ށT��T�YDrBB�8b$���V�R���VE�֕@�h�����?lR^�SG;����'h�=n��pz�>~D�j�c���m���|�u�n�/�<��]����A�7^j�Q~��C��ҟri<�H?z��0�,���C �]�[�Q�zgY�俈xWs�j����x��88���$����wփ`u���f׌i!!�8�V���N �`��<���d�h�S11L�Jʖ�Ydv� �����I�=���(�B������vλ�/�0�Z�d��������U/�l1-i�Rt�ߎ땎CN���l�o��Ӥ�w��P�fIȹ)�U�U%hL,ym��\�ZC�.�YRqc@Ã\���g1:k���U�2��RSe��e_�)�ȝ<C1�s�6�[bm�p����B�e/`�O���=�=�Of���i/c�<��_.�}�ދ�SK=O0����]><�/�E�ݛ��O�`�?����f�9ðE̨/f},�72���jLD���Em�w�A�ܒx
�@j�/&}�z�V���R�
�Ϣ�B�X�q:S�h-?"������r9�X�D[ʦ���@bb�1�o�n3GLa�c���R�����v�����0�,LRڛ�Qyl,��!���Х���0�o0A��x.��H:�4ƈ��#^mh'S1)Ie�{�S4�7�e�PO~ =�r��j����N v0�%} ��05>���~����ݖ�� ɭ���2���I�&!�ry��/�W��kN:bKu<G��{����}g��Eվ/ٓ�/>i��T�a�`d�[+u���0��lJ��	Aޠ�
&�����]��inK��73����g+��H1��;S�_(<z<D;��y �GGeK⟠;����/f
OA!��e[X�EP����3:b�' ��Vq��j�h�y�J�}3<��¬فw}swP7��4�U��D�sS(�x����M)*)i��.�8f悟�䎩���O+P	64��MǊ9�͂�Xƣc���1YM;;Y������.=�C��26E���j��ħl���L_�`�B���)i�n�:Q� ��v"~+Y�r��y��鰿޵����]���;	��<f(���`]��O�<ߩ^�����жһ�妧3��rJ�*�ܦ�03�����4�����}y=�|�� ���05��cdR���i�?'���Rط��ͻ:3VO�����4�N���9'������W���'��٭��wDL���@���^�g�OjzG��O��m|�X�ai���d�hp/d\6eԋR� �.��S�j��j�"k������QK%���4����l,+�(�Ƌ�g�(�r4�UA���DBW�?� �S�ا�޳s�q�9�;�vO�S�?��fF���	��C�'A2���N�ffz�`1��R?��p��IՑr��Ӂ�� �?lf�5>�H�X�eV�A®6�1��O��d4��ܟ�-�oI��'���Ӧj#:<_��|��&lo�h+�8Q��*�8�Dj��q$>`\	��	T4�˂��P�Ʃ�?�^J�o�GSII��U��hޜ�<��gUb�o��s|��x˽�P 	i�^U!�9�W^�{R���/��t�.9%�F�Q��Q03��q�!����a�i���E���U�qv����/"+\��5M�G��w�Х�>c6����B�P���
��'-&?��,@�:=Ҁo�mS�˳��Tn�TmV�3��`�R��:։�]ag�N�~Z��2W��U�@�=����,1s�A���6���a���Y�{��U��4�$���M������3�d�ːҘW�!�'ObbJWvxq�t�8���X�lL��:΃���4+�"�x�	Eȍ��j}b�`�!�|�)��X%�A��#���ȥv쾈p%����D0#p����Q��P�4�>�_<�����V�9j������VL"���/\f�����X�fƋ�X�>������~�z�-k����Y4ܮ�y��*p����U��sT�H��>l�i7()�7��嫂o�nZnV\
}��o���̫�>^
r8lh��u��V���8�h���B�I��^��������w�Yg������9m�D�p�U����J"��	���9�f�g;k��s\'���Mq~͘���c&RQ�a�?�� �K��	�J	���p��QMP�p+pJ8^��Ov����f顚�8�A�*�v
��6#U��|\C��z���0�A{^0��+�*;Ģ �D���L���Z�������6-��ˬ��G�u�,����B�`���q��Zp����d�SS���*�oaܪл_�����:D�{g��'~}C��`�����F?�T�f���@e`��X�N1]K��<N�m�e���h��z��ZF�}�-�'k'_	�p�`�z��?�H�DM;�����=���J�Ԃ�i�Ab)�����ȉ�@��9���k-04IK]��^Z!�G.��U�ԍ�`���N���u�h�̴�)�P\C�C[�mV(��e�n"&Z.@����a�ү�oZ��ʳ�s�����m��P���8y�0ýU�%�2�=/
S����� �%�k�:�˄���F]�@M��w�2PΏ���73�W�6 �7�s!���>�(��X�}��-k7�����6y��!�iG�,�U��q쏎f~���23>^��z���@F��Ps�s's�Xe���!n}aI��v9��n��E�m����dԈB���z�T"�2��A+4��Z����9���P��Ik�8g��I�$���v+�X@��2�7��IB}G	)g�e?�X�qX�G
,;���U�w�'(�y�`��������{��^�s;h����h���{E����g�v��Qrhzb��,�mg�챋m��Fs���~�gM�V�Ǜ�ku&��rx�Þ3P�s\�*(F2s���D��ph�v����dq��&�SۋPt�J�(�� 	1���g�:`�X;���;&�0�8�p���D�w����P�+4����մYzL��[;��,����C��b ��ԫ�!��L*�����z.��R�<-�y�N���*5�^�2;��
��yJc��ς��TO?0/4��~�QT�%�����0뉤B�'���������^G���2�F/�|3cD)��r������憑=R�M�:K�w��ڏ�S�u����(`td'�Wl��~gf�O�GB�[r�܋-���$*yb93F��)�r��Q��-�h :�P�n$\����p��gB���`a������5�c��/�(	�B�~� ��Ź''��F�s�]GՌ�B���(�Pp�磗����,�Ƴ��P���_�J��5��5�r�,4�$�S�=�	�3�6*5�����]�����N$�Ú=��n��0N=� ��\�Q�v yǆ�kx�����q�Z������-O��*]F8Q�0�#�����N=��l�H��jUb ����!�I�Е�����g����u�NDv�8f0{벧�������8)��r��3L��,��.M��u*9��ۈK�JD�F�S�}�wiqw�.�SЫ�ƉSz3�/��W= b5�&���������Y��Mv�Ц�oR�b���
��#4��Q�$���j��>ŏ���p�h[DX�r�S��qU�kT�{ojVڙ¦A.��A����_�������X�R�Q/O祔��mȵ�/_l���Ie��&ϵȜ�ѴR`i}W�dyrC$�>f���zc���]VA��w��^ �7w�K1��
a=���,�]h�f���f��gl�ğ@[�)f��;]�禛�W�<��9�lp�����r���o2o�7��3�g��!?D~%+�y�)�s�Ԅs���Hk����O"
j��欰T�GNG��j8`���	�dS�1K�(�rL$X�8;�>�C�|H����诼_*�f���KT�ϻ�.�E��f�52a��=�V�b}���l ̦D�htq�z�w�V��n���V��Q �.<�?I0�-� �><ٕk�:Y�[����2�l���+��E]�S��L�h���������oq\�̈6��Qr���[�S�@ǿ�a��.�&`?��eKarf�Ҩ�6}\�ݐ�"/�t���H�߀MK���~Z��\��'�Zᝈ<���K��&��Ry�Ny{pb�{|c��ίl��¼��m7���f�
�k��@a�>��T���|t�i��n�Ը���d�f��_<)���_&Eb��r�0u���9���I ;@F�HsRO�7D�?�<s��'ty����r˕fb�Zu�+݋x�V�p�hz�ry乍���S^
����ZwJt}�(v�^�z�=�|-2H��	�]���>���/l��	�?�m2V:)��'���L�j�J�2w�p:��ܯ(����K�m��TmR�bLɈ��F��܆Ux\~�"C�nd��0��+�J�ehQ���0ʈ�K��R�%��1>*�*1s8�<UE�a�ZA����i^q1��{8q�ъ?�u�E���I���u5����x�t�$ܺps���m�P���I2�&֊LdB�G��_�廂B��<�âb�~f�f��B �O3y�g����T�[���h�������6� _�D�`X�IsZ�\��d,KXp� �c&b�(��#��j��e�̮#[%4�Q
\�b�2�ha<�`)]���c����(a	w J��#Q��'�nyZo�<�F�OQ_�O8��]?4�C}��f"Lk@+5iؓ#��f= ��O� ��Ux}�򖔞u����{����/髠@�e|��
�ܩ ����#�J�x���l7�	_n��OM��b�E9H��S� c��18���,�;��sb��)� �e����.濕��&��R��A�}�� ��
9��l m�N-8��R�G��q�x�W�=	�-4��^ݒ�-��*i��c�H;1��7@Xg����ހBA$$=��u�F@�c���^��|�,�L��.��C�`+ilO)�rs�.�[�E"��
z��R=zCO�;�;}h�ذ0�<�k�3]��7���2B�3o�L�:+��zI<"}��W�;>��rx�CF�2����WfB�eҗ��v���\�7)N2>?���%�@�}��a'���M$��yq4r),���!���rxf�nEV>4h'��32I�J:�g�b:����Թd����,���2�t��zh�k���'�q�JKT��d��?=R�������B�=Rh~���Ā�xM�����b�������
+�^��׋�p�-Ń��	�)����ҿ�ZwV��:�V�eb�aLW�*��a,1��uX�iY3Cmb�	'�l�v���,�hy�^�t�4Q"��
a�\��+c���|V �_���b�R�����ֲ��q�I��D��R�0���l���6�ڪy,��魝�~R��K���`Ȉ��XFE�5��W��#�S	�O~�ƩK+����Mxe��a��ee�%��W�"1�.�@+�)}���b�������cw�,�tyep�/�T�u��y��<t�6���LHo)��S�k_��Կ����7��a���̼V҆i�paF��6f}��jn?Ǔ�)ޅu���#��,�ÓaĴi6��>��" cw���H��D�ˮ��\_?�&Sq~Ȅv�H?/|s�y�aG�|��0z���A��4�T;��oCĻ^�&��@�MoR���PpVw.,��I���G�^�)������(z����ٓ*�*GM	W�8�a�1���=@I���d/�f�\�6�A�.���=�6��}��wF��,d��}��ʾGc
iZ9C(�����e~YY0us��]W]G:����J�-��m���,�$WBt�d���p�)�~s��1%L�R���x^X�ڸ�<�D�gL�K0�amG �J<�*7"V�������j�%
e9:�Ǖ�t/OI�n�wn.��m�D���8���OX�ExPh�&=��@����[���틔5���ng���B��@�-��������@�h�Ìg���kZa��48S"� +�&w|�Z,v��ж&/�t�ly�¢�DRa^xZ���3��2PQ� .-��8�VU4�yڈ�l�%#����|;�<�Zk���B��L�3W9�@���sa�Z�>��n�>&&�r�e\EuUza`�L�;�Cp>�cO��ĭ1�����wl]G�@O��:��f<�I�O�o�V���#�;*�s^G�Sm<�`�w��x��c��S{庸NF�s�,P�Dt�$-��x��	��Qc��n�fbwO�r��ी�p?y��?���+���8A3�Tcq,p����pNx|� ό)eh�OGN�l"���9CQ�YR S�O[��%�1d���\(#3�F�U�$PI��D|M�R�Cmʜ�I?�4��OP���$�	��a����(S�٣���'i~�ZKu΋&���C:Uf��O�i8>����������.��u��
��^��YjNȊ��2� ��<��2 ����p^�'����t��f����R��%�w�3��u�b�6�����0�1���Ŝz�vZ{V��b�(R\�M���.B��P�HR
���ٵ�����S�g��vA��f�?����,�v�ʜ��d��p�aUj�li��q+���I������[~����֯.�U�'�=�D�8�Y�V��њ�IߞF�#�﹕n��� ��#�gV��_DT�l_-���#��B��<�{J�s�����ge��ȕ�c�m�>9ʈ3*�k2ӥ�Z����b^jZ��{`���ʪ�0��) �#�)��o+{����3aQCm������0�<���`R!���P�^��8���R�n!-X�6�x��ɭÒ���v�II��\O .�C�bB��K<��D$����KW�S�a���:��� gYF�2 ���,�>a~�ف���d߬_W�k��� 6�fo{6�c����c+q��J���;hiFS}V+ v ���T�ԽAX�����{�?�8��vK�'�,��c$c;�u�i�)9-���m�X��d�}�O�Zv!�U�n[��4�m��{�'�+;�M��T}m�e�ۡ]�~:d̮Ի��d\����r9�:�> �$���&Za�8���(2��n�A�/N_Ri�ڸ�bݞ�K���>���!��5��4k	��;�Y_���v��X����Y�M�Cp0 L�U� �Lg����y�@�Z/�os��[�#s�ڹy*�\�HB��>�!}i�~�e��w)�ErcҔv��0-�P����v��˧�G���[��^[�:eFnWQ���{�>�˾ͳ�.��o��7jWS:M�'3]�5�]s�k���+;��}h�L�њ\�'�'P�r
q���ۯ7�`��̓&'���KP�t$,F�h$L����{��g��l�GU�R'����6dP�N�⹔�倱%����ʷ�bXDzps�(��39-i�ٌYB���(F� 8P�c�ۓ]VU�K&^U��@;j��V��Z����ɮ?Q*]��U_s�<�R�Y������Ɖ#�ok��@Tz����M�u��;p�Wf�3�)×����?#wNF� H9�(�7є�%#'nw e�6i���@D<�($e�č�Mf�ы�P �A�+������h����c�I�X���ro��|n�y�*��כ���ɢ�����*ZNv�H�M�nGem	���֘���8�4�GaK|��U.�@��+v�c;����V:MH/Sl�e�Ȗis���8M�#@�\�R5*۞��&%�{���C����y*��29

ç] ��tH���Jv��{0֡��ֲD!O�G�XG�k�鿚9���c�M�F��%�Y�;|'m�BAN�B���E9~s��(��y�{��da��T��r������x�p����1l��=��G�J�p�ڢ�"�-����mO=<g"O~sT�T9�<�����7E���8����7mW�RZ
\�Vu����Ûꞷ$�á9t��+Z?O�F� ���a����~�}���Po�"T��B%������lDw��i}b���q��"���}5ꆻ>˹��|?��G�cxV�[�ߌ����G�D�Ka튮5M���EnR�#P��������c�>��~_A�\�T�71x���6�����w���95$�В*�=�W۔-����z��x.a�<ó�J�dP�rO�G��-�o�G3�Q�V%&x��ۏ����_F���EE���+�ȚB���@��uyD;������dp�-�8LȐ�f9�B��#��\�E^u���߃��I���2R�%����=l!�4L&��R5tc��|��"2Za���ĭ$9�M`\����H�"T��U��-�k:IUģ�GC�Ix-d�`V�,*T�DiWtp^�/�3�'4S��2^Y�²is�p�������y�B���]�ŕ�W�����]#/���O�����"����߷�8V$@z���KK�g�y"μz&�Q�o�ń^�g��ZZ��5�f��e�# �'//Y�.������m��c���׍���M^.�?���wz�,�\Ŝ�v~�dJ�l�^ݶe^�=My�U@�X���8�k�V�U|$����F�@͎q��ܺ��&��&©�1B��l�ĥ|�Q���u��w^�w#动_S�ozɸW�a2�� N�b��m���Y�<��¹j��+2�@�C#p$K�M��?p#����m L�72PM,�Hi������f�V��G���8H�G�ǖg�Y)��Tr&�K+Y"�J�B�9�{*�ɣ�˷��[�$�5�j5�>�w�4]|V�6w�����Z�!���R-�����W�;L2*Y/a��|h�e�������e��I��� J{َ,��>
��=YzA����п�N2�;�X���Mأt�X��PZ?Q\�D�o����o�ȄA�UH��4żŵ�w���E�A~�v�q)�j�M�C��6s3^��]��SD����ʒX� ��`��|*��o������b�M���t������=��P�G8U{td�����P�.�h���<QLc�:��n>2�k(Ά�&|?� �C�s�����|~Xp��&bo�қ`^ܬ�ճO��s�_0�>����d�/��"�$�����>'GOX�o�:�#�T,:z��qN��>�YD��4# <��(E�q� ���T5���YUn���P�Y���;GZ�JK��R�s�$g�k7����!�-����$�R�@[R��ҳ�3{�I�t���O���q��h���a!+���,C��k/U`S^�W�=]ܶ汹i�&��'�o�g}U�7Bm�O	n� �@�w�THd�1�������v`7._Ohj���w9F� ��r=���ἣFWN����,19��� ���f�NkM?�M��=��me�m���~��������������j @aw�}��2������G��a$�ad�7b}�j]T?5��z�m<���-��b~-v\lz�?]K���)+��;2?��zCZa���2�'�d7��#�%�&C�;��d��I�����ܨq�gl0�����VRi�b3~��Ri��9ρ' �R��My�U��y�T�7��3H��u2�+l������޹)?c��;(���������ړ�|�>�����h�$�签���)z\NT��<�ҀjS�x�xt�e���1���ٍK���]��"˩��X�7�'�;�5��(���{�[�5�4�����&�
v�s���6*����T~@ِ���s��-}ic������}�6�(Fp�]����/{���:�e�y'�" 'K#�%�N�q�~C�,��=YLy�w3��}EX���(p�4�j�o$�GԈj2�ks��3T��c���9�O�+G6Y��Յb�
{���uzw��(a
���7��]ǩ�k^d$\
**-b����4)	t�T_Bi�5�cP�B�o2A_�F;��9#tH��~򽀹i�����i�zgJxe��,�;���`�T�:{*iO	Kb�@JHO?#�K��?i��������!�`7�3��a
�6��~���+�U6Y?U����k�Z�G�@O����YA�~�*+
}NL<=0x0�ZFJ�S
�g���	%�&�ʑ��O���e!Y�k�SI�JN��u ����K� ���yܖP�V"wpEΒ���G�u�0���? �<��72^�Op�Ѣ�u���,�	^!�]�3R��2&=(v]�}�D�x|A"���X��"�-?��S��G����h����#��\��Z�T@D@p>��c�
��n�{:=��v�-2�b��9�%`6OC�hF���ӝK*9vV�INR8KZ��^Q찟�z�,����~�� 4�<i��"���h�����#���gÞRA��� :o	��7����*!�	8cM�I��U5�V)�0���)�e��	�Eb�h�u�M�5F�� �P�l����*��ӄ2�� 7�>��� �J�n�
�b��qn�f����Ök�Զ��k��-�v�^.No�8�s���ߊ7d���B1NME�cW��
��7�ћ5Z����]p{JQ��������5��5���X-IpXͻY ٥���	�&�r��̀ �3"䞮R�D]Y#0`GL����VXU�@��� �վ��O��,p�8�St�OF�7��sa��38,�������B|��[E]�?�*�22`X߯FO x2G�<��߹+��尲�ٽ[��z�8A9*������:ɇT�pVKP	����тg��D==���9�QE<٣��=��]d�`��.�3"�x*ªMD`�Ȑ5-M὎{�|@�wݦ���}6X��"�A�?�ʹ���2��oȸ�4�U)��)^���A
�]�]�e{J?>Le�G���CU����J��0H&���Q��g�(N�܎� ���?���ӹ_�vΜ!�ElB�:�#�_O�����J�-Y��&�J<Z4j���o6t�>D���"p��r$�0 w�h�R�����"%�kD���%���t�7���IK��qz������r�����D�|�0�U��6?��S&t�e2�`�����&5I�`��A�^C��2 s������ ��Uo���Z�\����`��;W4��_�n$��H����
\���=��M����wr���O�}=��v�[<�y	-�D�j���:*=[r�D�E�����QԴΙ� >�������%Ʉ�@Wb�C�L�ד�N�g��/\����q��M��]z��
i���O��?:�U�. 6��.
p�e�:������(�a��cp�/,l|�9�-<�s�|��1{b�]'I���)Ve�tH\uƋsKl}�ذƨ�A;)��o�#[����asG|�r��4\�VJ)��;�'��HSg䶰J�:�t�m��?ȭq,�q�Q.I��n6rO�R��,_ZB��Q����k��$�zy*A;6���K����ޒ��v�]�ے���Ǻ�����y��67+7�Iv+�,�q��X4�5걢�>8���v�F��n�q�;İ_	7�&��sYq�z�.�����>�/�b���FF|��j!��h �{����q�[x��Ms�L~@�aX�F���N]�I�E��U��m��T%��o����Y�G���A��%e1Q�20S�Q ���;�,K�'�������3X���!�!�@~�{��:p�W������\��k��{�"��ZL��,L���61e���u4~��+jtEp5��i�b;I�Fsvap�"���n�(�+�� [/x��#����bq9#���x���u��i���'v�Vbd�H�B�r)���P|�	��<TR �d("N�Y�R����V���ϼf��Խ`)�`sb��|T>q�Z֪ёX�<�r�.k'��ݔd�����sK�)�-��(w\�VC�姺Y�J�b��/�G�e�f:ʔ�\e.0����9�bd ��c��k^i���D��7.�U˙��L��rJp[����6ю9 ����e�;�]�_Go����&��������1�?�X�c�+@jѡ�D�v��&d���t�`'�!-��$�p>,��x��xZ����������D��(=�4Q�I9{��<��5����'>��+nD"�e�l�j3q�>�6 2s<=�`��y;�#� K�	�;�	���Gsd���ѓ'�KUA�7e7���$�\�n&wp�|e!-TB'�c�Ϻ�Ɇ�0���k����%��	VO4Ԍ�Z^ͷ�ő(��g�� ٯ�/��U!5yE��I"���8��	��LP�E;]��/x�*����Q�|��JL�V��;����!�Y�I4�X���Lbno���|W����FEx
���P.�|���H'���(�:��"�[60��-��t�TLw��אD�x� ̐d��ͲδA�g��>��3�1O~�`-ͳ`��o�]yFxy1YɡߪR̗		����8��	,��A)?W5�U��=�(A2b��oF3Qk��Y&�-�F��s�%� 2�ͪ=2#*j�\�`l��!��x�k��V!Dg]艜�U�����Qol�ۗ�E�1]��u��c��V��!H���t-�k5n�qؼ���ӐN>Za�Iv�a��>Tn�D�<���۱�0�q�ˁ���'ğ����������?�^�Ϻ�/�!��Ԋ�ELގ��k���O��`�V�-�����
[��D��s�H"0��tAX�t��vm4�� '�B�����ȻHd�m����#)n�Wݮ��F�~�"No�)�r��R�
���t�*Y�S3� �A�G2K��Mp�j��x��{��JG+oYw��J���Z�� ���o ��0�U�c�l"�{߶�i{��-d
K����]����ǔ��D��u�wu���KJs�mQ��͉S��	'�i���$�^�F���.��\!�qX�f�߯WU�i6��3���s
ܮ}_�էs_I�"�������J���x����ư��p�w��R\�ѐ5F_�&)���/�|��?T��J�Dc߇,v�GO��.`j�B$K[��D��w�Ɔ,	��G-Y��3����׼�Kh[�v��8}�E�.#���v��ex�t�Ǵ���&��dֿ�N��ڷY��qU�d��r�a�2���l�߿�i/���El�\�:�rUdk�2:�:�,�'P�%s� ��L�++}%�y`��j!�
�Ě���AE�Jyq��D�af76���Z+��}�ٿZ�-u�D *�#{&H��:�<gq�F�����K� N�]e���G�{C[�4�z]�n	��=�Y�#�!��S�g$P�G=� ���^��\N��X�.>�;�3)�9�'�DK�a���a��8�#�^.y:[�̓]#�~8��SfO^�]�����ڥ�p��3��M�4�r<���5��'�Z@g.��0AY�ڠ��v�	v�Y�V�&z�z��u��J/W��� ���Y�`z�սr�/۾�3]��9�WC�;�u=*E��`_5���.,sι3�x˯0f��5V���dEL:�ϝB|�jzJG�O�:f���G.��O��g�s<���ݞ����P����ݐ�����$��x��U����HqC�[��	�@��Pu�)�Ҧh��RkK��d�6�s¨���mާIƱ.!ۨ��d�vN��
1��]�La>+�pn,Q"$��q�$�6�ZA�.w#7��4�v��(� S�����H}w��A��g���40�+��8[�j���+��ur�PJ3�����MR�>��d> 
m������=��Z"�*��n�n��x��!{�EM���l
���K��*�X�)[JK�}����
n�e=7-�Z�����Fj��R-D�J��`���>�ӿ"u�D������O]��]���34�67^Ev��U��N��-��G3�ժ\fq�$��;,S4dUo�|�b�	v��#�;�S!Yf��P�6�,M�̦�.U� G|U����&�Ǽ��F�|>�;�t��ߥ��)�BV�A$Z��K�`�
G��B�	�2d��"������N�ȀW�������r���	_��-9ӼP<{B�%ɛ����6��� .�+�@�4>Ӥ�E�=�ƌ�6�4苰]�:	����G�r)�`ԪH�;�[�����Ì�h*�T�����}&�m'��1�3��^�Jt��V�7CdЩf�q��TbU@�][GM�
S�p�Lhk��B��9�~y+������S �t.�`؝��r*����a��āXY8i�*�����%�7l���%��f�x�ؙD�+V?ֻɔs R0�nª�L��́����tz�U�؁#OK���e����v(Цh�n���`_Z@�g�5鳹"��p�O��T&�? ��#3D|�N}v+OB�H��&��)W�O~�|ǒX>�4�Wz�q���>Ҿ�O�_y?*�+F�:����TfPϓ:�ybM�󏜃%�3��}"q%�L\��3��ӈ�*�_�T��IP��+����?k]��T�[�9�]>�k��b�𱂊��fZV���,�C�'���:�p��A�J����N��m�@ǂ��\�^� ��>Yz~�QuPUĉng����L����} ̊y��}�j��_�D�SvUe�{�5ȃ�
@&���C~zn��Z���pWZ�����;��b���Z�8��j��k��*9��q�D"�'��3?�03��H7~Rt�ʘl�
O�x��BN��� �0!��4�/_J؆rY1%�/���2�q�3� �i@eg�91��/=��dx)}�"��;?�X�0]Xb���ܧ	��|�iA9�H���kN��G�gҫ�k�ᒕ��b
.7Ro���6[c���#G>������[W��|҆�.��{~+2�ў����aע�w=��;�e@��1y�����]��Z&�XI�hy�#-�#�����}�kk�}v�oi����$u��`����������Z]40�-���%cL��<5�(p}6\���<T�3�c��mX�Ѽ��e|:9S߁�6����\"^aH�հ�������_�g��O͋�yQ�mkc8d��?�2m����L1�U+�)H���˯�5sS�~�9� Ŵ:ؕ��.5�Z[�8�PGC�@:b�wHS��U�R�_y�
SS�-�d�R'�.��2��BZ�N^}�D2�v��\�g\�{C�sU��O)'Ǚ=B�������B��R#ǜ?l�B�����;B�|�xs�K��I��ѵ���T���U_"��eVW�"��ug7��߉E�_e�%��z��P�=��k\��]��S�|���*�ۋ�C�=��Ѣ��< Pr�I��w��fu�x9b�B���w��4q򐉤��{7H��6�;k���S��Z�`����	۫0�O�\���G��9��?^�TepG�Q��W:t�ō�KX�G@�!>i8����I�B�Y9�'��̊Jʮ�����X���؞*NA�uOOZz	��xF��]P4��ϩx�j��M��+��Y]���|�2cs����r�)�e���qۨ*��\��.�c�PCr�d)M�3x��x=:_�ұ:n�@O�І� M���2+x0�?��Z�j���6;�����=�S�@��԰eH�!����݆��M��U������E���}:K�\(��@L~����vQ�:���֟���	��τI�?Fҙ��/����(����3��K=�n�>wbs$�j�D���)�>���C�6i!�<��6�%��T�&���	\k&�Ƅ0�Md����5���ȼw���ۙ��4
�5#�D�E���C7���/��ܗ�z+�K�\r�||��d]����2�C�\l�����;Y� [�j�ws�vX �0o�E��>ѵZ�?,��+t��C���i��u2<K��6��q��j8�%.�F�z�(�oǴ��+��jF|���Ҏn��{�WO��>���P6�T9y��Y��޵���pF*�cڲ��'�,�:�ܞ��!� �e�Xu�f¦��\�V�kX I|��^$��x7�/��ꊯ��BL�#�5wd�x�`�`"NEf�����V� :n��I���ޤ��b�Q���N��f�b�E\Hu��#��� ��Gí�B��I���7@��Z;8��2rF�����d�~�����c}2��g[�㤷�\]]��Y�Ü҂ħ�U��C��r�#����}s0'�.!�Ԫ�iu9TE��L�.2O��q�8N�^���z�"�S�"�2�m,e5"q��3���1Eե�9���
�+5)͆�F�a�lP�L�4=Dæ�Bg7NO�8�Aa#K	,�����*���c77����%�]-h������W�M���ٻx�G>�,�ɒ��/���|,�:uer�K\�r�4|���OEs�w2z`��s��h�+GY&�sA��iT΃�t5F?T����B�),������y��9�� ����˱ ���?sjމ"�&.Q��Z���$X�eBǵXG��:����?���""�3������+�ˠF�{|0mF�ŝ�}�=s ʇ���'[��Tj�+�$`O��/�;��Zƃ�ۏڳ�/ k��1dC� <���T�R� =N��%���A�R�č���0I8/2�`��M�����,,R��`Kf0�y?#x��/%���B���������Эh��';��;���"es���E�Dzz#���c�ѿba4�����K4\�͍�,C�'0gz�\�i��Hk9��,� Fc��T/B��o����{}���Ɇ�H	����>���y r�k��|���ִ���J��&�6�%��W�/M\��Ne�`�ا��i��T-ܹ��@'˓������w�Z+r˽��pdr��r�O���x�76s'C6���C��_�{�X�O�GƮ�K��K��(iN\5 ��F���4U�f�bh}E)���yN����/��u C�;��Q�:��[��B��=�?cϜL������{�O�"�C�JD��8�L	/�~
u��h�R��p�#Q��C<���<�9�Зz�N��c������x4m���O�`kBѻ������o25��A��Ō˝Q����WE�R<��U�֩�邰'�&����rm��SR���
��'�'�^���%'m�ŧw��9�*�f��%n�X2R��Q"�R ��^*�����*~�]¨�D~"���G=Q�m~`�.
�|�O �ΡA�Xޣ��i�0��Rن]~����g��,���a���ЧWzC��5a�#�����Y�!H���7GR���h?�rWKӂk�Ub���T�;yfu�8�<V�Lz�wR�,(���±�ēW��RN���	�2�,ߜf�x��\Sbb���.ӺQ<��i?��ϖ0�)$>�K�]�^S7ؙ�z~�A}-R�H�/�_&��p"�V��Ӊ�xؓ"/�T�.�;�.�i��T��6��]B/�ٰ��-��Ѥ�x��/�@�ԁ!���>�e9��ZK�g'~Q�TC�e��"�E�܂+etM��^���}�;*T�؉E'k�ŧ{�ϓ^�B`
Y;����CX*t�'�F��t���&�?�?��^���6�#Ey���Ck�����J�M��9d�wm�9MFb��������c4n=�~z�������Uk����7h.2�ז�xBz����we���G܇.?\����ࢁ�;�kS��+���G���Pl&SV���'�x�0B Rz5��v�V���ɦ�6V,e��>��&K��%T�rߔ�0)N��+����ψ��樾o'�<Bi!6N2��"|؁��X�}�%n���gZ���#�;F���4��vT����I`W)�|J��2�Y����Dp��#�Dĕ>쿻'�F���б+����<W4Q\�e�'�{� ���_�{y�Q���O�EM�%h���^#�^m.��R|z��R\���Ǚd�p�>�. ֹ4�v}/��8��!6�����M֥|zy�w�$(�چ�$ay��vH�G��[���}�AWo4��]��'�� b6d��6���6�jZƫ��z�o�3���E.���GC�K�%�u,�8�&�ƫ?�i|ko>V�K�|������^H�����i�8W����<���,������ol�H������5��إ���aA ��u>����P�n~!���6+z|�^xn�����H8����Q��a�
Np|Q'��_+f����i*����M���Bo�aP-�3��>	`�60�+# v$�JGg=�|Ϙ���|�O�H��H�J���J1l3���(�8_���oo��إ�`OYЭ��o��`6y5&6^����nB�Z$ D�@gn�S�h�M�`U���Ɩ=p�!�~�����;��pQ���c*�)1�nAZK�g���J������i׏��2-�@�Xva}�W�ŖC�H�j`���4��2��$U�>{5D�ɻG4MF��<�HJ3��H��R�P������*��Rޅ�V���z�Q�1��:���4>;�������H��d>u���hu��|��l���3K�2歷�&�m���¦!����E
S�|�.>Q��9HG.�;,�>p�n�(Ti���!�h̆n~�_"b���rl�	�������R���t[L8A��\��0P�I���!N��Yv٤��_���5tIw��S})㐣x}Ҵ3o�g���}��#����g��`�����������M��Zկ��=Ť��Mp�}DC6��;0S@��@I�rJ��Cf�ovF���\���5c���E9��WGYu8ks�; ��'��X
��ॽ9�5e{u�� NOemk1��<\��V7񸏉v��xs�;�E������s� �FC`� ^��x]Y�e�Y&N�`�P3j.3�;���z��KO�n_ҦB�qΒ��m�"����̗P����M/��!��qm&��h�]��z �F�����)�^ф�)"�O[[�������a `�[Af�^�����������/�G\y[6K������Kf����S041�l�p�$�+3y�8�CԊ�$�
������U��G�p���sN&h,������|Yi����Z:G;��bP^� N�Ā\ɀ&��q��V�&SQ%M��_Ǟ����,�>�y��:���!�H
�j��WVh�Q��W�����ſ�Z߃ �"=	�)�׭/��V�Ӿ��."�8�����l���%"�$���;�*�fM�na�涥~1� ���Ўcu�+��/[L ��y��j�}ЫC��.q}��cfj`��+����P���Q�d:_~�r,�@�5� E���Ŏ�.\��(=�I+�Q���D\���!��ϖ��T���Q�h������!����7�a��_ĀiF�D��l�F�-�L�\���A�,����R��^�[��_���K߁��]n��%[̙:��ѭ���!��*s�nw��Uq����p		�7���i�~^���*]�Q�Ӎ�*�#/V�ˀԶ'�_��Q��c&B���G��P�9�r�p!}�Z]{�]�{�p!��x|�$��O����6���t�;]U�RA�����ʊj��GD3dx���o���{��+m�F�i��.�jeX�M�;�! � %E�؁cݟ�S]�;�C���Fi�|D �*�˩:��pL�M1���grm�&���]ӤIQL���\Ű���v��qt�g0s�M�-���DR(����n6!Z\F&�P��j�oGj0ɛeB
��6�	{r��.��8դ��|&�>���	��f�=�[ND{�B#�8�ed+$�ܶ��Y�-ȅK�ꁊ�F!4�X�y�,x�P�}>�2�}���y��C��c��i�wa���q��F����L���5;X�qC
V� �B�V��osnZ{(�hxFav��NN\�Km�F)B��T�����0N�A�J�^еnQr��Â�H1;�6'�U%�l���;�#��z̮ʝ!�P�%1��L���>��<��m�5|�r�y�AU�W�?}��H�Oq��jbc6S(�z5�"��"ؽ���t�}�r������mU�U����"�X2�.������K��~�μ��(&�D���}��v�R<���c�~��U�Z�����r6�l��9^T��[��� f3K(�,���1���e��g0�Z���0��:�Б�u��	�$�Eŵ�b��O+5��|�����3��I��1l��-(���7q<�L._�[���F<=oC_,�S���˛e��A�U3�����#D�|��m M&5��,YQܰl�-�Ћ�{-��{́�R�iژ��Ӣ�#��FW(�mLpHK������G�=�UQO1`�5	r�O������ط�������	������H��-��(wg�� ��=⯚���r����ZA���Y��H����'��bZP����3���H�kq��V��zv���'ĮR
ez':K-CNW���������f����wYXu%{��
G9 f��MV����Z�:G�r�|KM�����K�8���OHy�vJ�8�\�`J�Q-��̜��;�\�P�d�s	 ����Iٗf����qI�b���0:n�B�T�j����yp.l�ڰ������)&e�Ū�x?0�D}�'�>�2e��=2����1o��dW�a�ფ��^P'QW��P��oP����@��2�T"���]daUQ�5q!�W�XK~���j��< �F�'���T2<��q;��H����`v���q��F�y���x��tX�>�t"3C�w�f��ZQ�Qo���f��PcP/*�0��j~{�&���e��m�6��JLTG�N��0K�����pˑr����k�R��wT�%u�����lN�a�t�t�g��zH����jn.���G�h�y�"���~"�гVRV�Y#��S�Ƭ�����=�׶�$���R�lf�����$�>�M��=pL-���uK] [����N��쌪WXY�!@g�Ŵ{ׇ.�	��k�0�����4t��H�-!�k/2W+4�P%0�Hcq�SAi�H��*c6K<M����<3Z�f*=0�k�-9�?gj����5t���:y��ʆ�
�[o$��hSJ1�F�-1w�� ��wI�����b�%[W��sY��>����$Y��Y3�U�P�!�ܯ�2��rK�d��W�\��Z�iG��#����r�H��Y�^��-�|1t�W^�'MQ�������N���5~�F[weV"\���s�(Nb�T9�����Ga�G<�a\�kq��F5j��4�mg��W]��0��*�����e@�v=@�Gx�&4ꄁO'|�����LM��2��ǎ�1x��=���ܚsĮ�P��~+@߸�헠xۛg��"T3�Z*fc}ޚK�BP�
�Q<�l.}�g%]�}��W���v$��z��7b*�݉YFl�<n��4S��ֈ��z�c#��	؂V���4�G��h^g��d����W5qj_�	pY�@�3�	�%�[O�[�o[a�vw,��o�����f�(��W��^�N����ہk�$h�6��}�>�F|z~B������y���Mg%�0�]��1�b� ����<�������[��a	2���:���?l�U��p��V
�������6�)a��!ާ�(�S���bk��	�>�Ƙ˵7���XH�T��Kނ��3�T���@
�!�UtRDֽ���U!%���4APr���;H��z�pz�`�(��^��mʞD���M��f���p�x���{V��5�)��|=���a6�BOB����d�������2���#0Aj����ٳ��MG���r�T���px"D�O'y�AH��쥲���)���f����T��j��T\���*i<&�u�<������ɳ�"3\�ɐ	yƎ�:��Ie��x(,��׳I�?�y�"pbJt~/S_͇VWsH���'����(�|��,� ���+�y8B�i��F���� �v�Gz��]Q�N ���U!Ui�� q-a�>:�?PN�"=P|諟�C�[�}�V�I<^��w����B��@���b�H�
L������ �=�� �~��'��%֏�ݨ��`W���8�F�c$��!ω��:
_�+k���N�.<�����|�V���P�O�o\�(�����]�m�@J��5���rf�����KΏ`٢w���6��t�r��iɬ,^���	�	�����������V����4��,��Ɋ)t�D�ci����'��0);;q�}*[�-S��K8q��(�59Q�<��J~Iʌ1�$�հB륽	t�����Ҧ���9�^!)�LI�T���j<T��,�<&�*��)�X�>�|
��v8�nt�h� �����_���[M(�^��mw>rAl�v���;z���_��֌�:4��y�8�7�
��	Vfx^_�]{Vہ/�`r��?HC��?Y))��]�����W�gp�=zs�PHi]�A�n(x�M_$�ʎ&�ӗ}��Z�j�
`J0^�ɶ��5�z����A���\��T��ǿQ�t�J]��J�_U��Z淓���_�8��i�Y�DvfF��LC�W�W�eN��I ��wFO��� ���rʭ��Rݧv��`E����n�5E ���G�kM��Z>ܛ˾lm-�u������W��9�]��&���m�L`h�#�,?H��fg����K�!��?n��(ھ.��@Aˮf(��f�i���*1!ad	$����{){��a�!�n�x��=�N�
j�|lO��Mٌ��Ȣ�n��������䦹���B��]�Dl��R�7[q@t�f�^�������`�2?,6 e�~Z� �����ho����(_ ����K��#_�y]�/;�4N����)ߞ_��⇄��|���O��%;R�L� ��k��E�5Ӗ�Iz�~�]���`ױɿ�0����`$��
�V���D���>
-J^rOJ�0\F���ͻVl�9�f<��s}W�P5SG"����߄ M�J��$��_Zp�C�Ӯq�$C����1�y�\D��j�O�<?��non�/�.t��:ֶh��l�������*��o��o�����bˍf����]�Yϥt ��B%2�v�z�ɋ�v����A�Ʌ4DJ&��?ԉ��F8*���ZL7�H�Sh���%-1"�%t�屋�R��{?�%��	�(@�������o����}:ÿ��%��F���V���n�t5M!�p��C��O�S@5�����:��#��L��L�ږa�٥�R�*�"�Z?��$���V��`��� �e��&�}O�q�b:�`��m�@��M:�k�t�m�$�"7�pnd��Ԭ�Hi��L�Cp��8&��G��W.{)�gqk����/ df���.���܈�!m�a
�J�}��Vr*e�9;����9�H��z%R[���쭯Vt �i���2�@�ߦ�)����F�p&+xRN9����� �C`�_wڶ����3!�%4�)]6e�.t'�@_vf�T����^�8���u�\򩞥'��A�N'�L#���'~��H��̻�_�a�H:`�P�r��X��UY�����:�ʇ�i�?5(Z��i &Whvv*ַDP-R���ivB���Nd�`���;�x�띆��A%���a�cZ	w`����Q�x���yY��Z|R��FS��Ɩ9>��Z�F{�=�{�C�{��[~ܗʖb<@)nj8���R(��2�F�VN��5�;lS��0|��y����Hk���Y��
����<������!�U�Yc8�YW~a�5�S0��f��H�/�S��A�_ȵ�!zn��p��k!���1��y_9�8m���|> ߆<�ʷRR4�H�,I��R�I\V�y�cs^�R``���9��u��N�?!A|J9Ԟ��z8����o�o{�|y=�Ϭ���(��N��6����c�3�(�S	]�.K�x����_�X�N��lJ�-�LhN+}�{���e�K�a�Tg�*$�*e PB:j7�2��媊)���O�bkfl�$�.����u�J�r��S0K�y<'�?#{�b'{s�⺤"���V���oU��,��< ��[g��Ol�:vO�A�&�_�L�{�.�a� w�gy���7|`
�4`�?�]���@��hȔ2�������N�l*��lY�
~.
�%C~ �uѼl�}��I�nbQ�$�eϠ�.�'���ʢjdq3)�������cDF��(6̒�%B.�mRc�/eV���v|&0M<<BՌ�t��=�L/���*#նN[ �����O�@������i��n�����7G��P��A?+=!F�ׯ�=���W�#�Ɔ�w�Z��ɾ, ;G��mqk؝XJ�試��٥C��=�?9�է�l���
�?�j+��Bk�Fy_YF\��B���ϖ	�(�<�%��Mx@�zL�(|!}f��!3�C��m���x��������F����x��V�@mz��w���Xdo�b?�l}G�֋�:�����\�iy�W�����?�ջ�`�z����I�آ��%��}�Q��.�oE;X�Wh�30ϩ	C�>s�����C%�p���#Y&[���UeLm��$�}�M�����S-���Z��(����N�
_F��g�S�� ���.ԕ�~WI��������x5��b�{��ҟ��^�iڴ+e��ZS�5����vj��+�+������,Ç5��{�������X��c{��}m3)%m�k��E�د�U�������V���Z�/>�<t����~Z9�;��s6#{u��@
7�C���d)HE���"� �0��|��D�ݽZ\�[R�|VK�����>g�z��ِ�4j��UO��,u�����6 rކn-NB����j�� ��_?�ez��bRi��ǲ>��Yu8�=�n(̱���0����U�A�A�_	h��$���Q�G��zT2�Ok\��`ȭhý�e�1&��Nb瑛�\��K�,މ�hK[���K�e	��p�7�
�	�`b�xW���cFC�4�U#�V�����V�����ǁ��4+j� egMK��Z�;X�G������5>U
�����M[��x����ȀzX�(�i���B�u?B���'֧P�]y�{c3[��S3Kjz{x�e�>��] � z�Xi�d\���S�r:+X�f�A�
��X�{��Ц�N1>)׆�t��� ����ID�_O��b�wt�w��P�gzr�I�7`��p��x[�M�C�=t��S?�<�͕��R��z�-~d9�1hK������~��k�Q�������sR?�X�2�c�u[ouS�T��� 2�H�I��,/�(��/^��ͨߕ:�j�3�-�Nm�Kj '���=P�R"�KG�W�K��O�h�]6� �Vk���oy�*x�R)��8)a���n� ��J�`!�i�,���2�=��>%
�'_\2��KUz�N�t�o����gb��c+��|4!~�,������؟�l�t�^ϵqĵ�d��k
��+ ��~�f�{��g��ɭ�Lؕ����-�.Qm�v��j�<�u%�5#,��(�ܑ�Q�A�eV�$��U@�|��DX6���&{H�;�'ظ�0N���U����1KV�j�~��t�����ᜠ��Mm���M�r��+R��q1��"�n��Lp�"�(��L#%�I����� �����"D�|RlGi�A�Q�˞(*�?��r���`����.}^�������x"+mXP-�C��ST� zINb����8�_�y�m����؀t���Z!j��'�Z��������nQ���I=e�����fI&cqi}q�E�k�՗��s2�?L�ր�\�\���4l�gY�+:eq8��'>���������j��;�v�V�7��GѤ�>�<[�͸�cQmNl����:��x�c)!g�I��p��c��e^t8���4�g�w�߫U�c.�=WV2MZ0q/.��6��w%p�~,J8�]��鬘�b#o%PbJI��ٸ����z?zL��cц�S�KQ,_���/�J�x�q����@�?0p�Q~�q(�l{���Nx������E�=+��Y��M�Hj-;��mgZb��k���@{'X���W�藍�DV ̷�-#kS��M ��Ǒ�#T����k��a��{W�a��gH�j����ן=��E���a��"��O�&¡�d��T�n�^���n���<���\HЖ/y�=F�U�2�^B�O4��Ϧ)�-3I2����y �KȀ	;��)���`������s
��Nk7��a2���a�?EGF�X]}�OW���-zEis�EM����Sស/%��f�	5�\�0PY�%�{��,"ߟ��A���[���k�|V��j	bJɿ���zw��hSߺ�g�,�����k�;)��T _U�.הZ�xѮ��"�B���>�+�K�������'�D'sv��0Sz{%d�w�-[�3���ݤ�͡&\6�0p������ʶ��,lk������Vj|�,�I�_�I�[i��Tct�Z��P4�)N��Be��~�#�D���EM�)��jaj��n�
y�՝�ԫ����k���<g�X�gC�y����Tx'�Z���t4�l���hT����>���zvUy��*�l�&[��4�;��ɞ�@�����[�j_�%�TY���OY��H���\0�;���#�4���[��z9��A�fՇ�-�svx����fk��/'��%�D��3�vܩ��I+	��ŘW�s�
z�Ei�����c�-4�gyd��
�Ise��hzJxG|�
>�BT�����K�
<2	"�yz�hKDN,�$N8�9�pF��û0��mZ�p��b�f�b�N<�?dh��a�������������p,�U&�^�8�^��~*f
-J/�P�j+�~,0245�.�Fјj:�(;%#����yzdQ�͊&��D̞~�K	ٯ���`r����!�e#�c�T���o�x�YVy? 9QQ�P7�KfzH�&߃��9�}w��^�m��zʾzz*�T�����wO�^��λ��B6X�wذ
=F���$���AU<@�?^)D�:C°45z3����.��a��y����������'j��S��=��?��A�$�Tn��A��Reh��ؖ-����
�l6{�m����㎎>��+�Ne��<s�ųـ�$���N��E�� '��T$ހ_�|�Ԛ��s�oS��7Y�����p�.ϑ�-�,�&W��%b" �k�]�d���E��$�<��`�z��>�R��v����������F�5E5v��@O��=
�	���'��ZE�����
;��a�>s(f�P9#���.|Eɺ1����m�q����_Z �F9)j�����ͮb�0�59�����E�t�KM8�"�m$x<ȏ�7HS��e�΢�"�lc%$��)��;1w�R���%�M
S�Z?|n����/�����۹\��7�}1{B:A,�	������C��⤼~���%�zu�A|Ӣ�����ú�ˉ�bc��=���6��(���4Z�A#w��ܦ�7.r�U���sQ:{�Jl�f�- ���e+~k8<�U?0����2��ҜoŮp����q�~^]�_w���R���9'^��K`%�S������m�i�����98?"a	����O�u�I�cY��v5"��i�`�qf���p�ү����(wcL.����vOE+?�Z3�ߑ9�2�r� @|�8�9�`��qiԘ�V���kb�x�/���R�pۜ��Т[C|ےr�8�l�B��R
ib,RP9�����.:�HL+�����M�|��"�?��c�MSr�J�h]P�E�}�`(Q1=|oY�N	���C{S�=v2g�"��L���ݭ��/�d��hI�ׅ�Ơf�2���es(���8?/#1e���,���'j�.`�~�\i1p[��T��X��p���.��aO�і~W�MM/�}H{�����i-�0��v|����(�3��U��R6Wk}!_Em�6��B�Ed�:���WF�88�������h t)����̩��o-��� #l�������p�6���r{��+>�^22r�I�����['�',5��s�L��P�/���
2	
s:����E�L��{y��"���F/Wz����6ȚM�)1�s��O̶n.D�I��p{W�r���"MY˯r,�{���9?z*{�Q�QH�B�,�Z�kϪ����/1g�;�}1�@z���&�*���\�)�>5�p�+���_�8�_Ǌ��)�����\�E�u��*p[l�Q�T_!�ؾ2�!�P|�q���
���Ì�����(����m���Mo5�D���c%ʠ��D���w�Y����m����̂��z_����q%%�z���T����O��_��l���0�J�Pڶ�e;��a4E8����'�M�#��&�}�,�YqH�N��&����8�+����r��zV��pf;��k��F���E��5���B�+6��o�j���&q��!��YQss��r���i�Oj�z\x�U��I�r~�ǯO�0~����3Ê�� � � �	H��hpK��%����1�uᣫ�o�;��<H8�G�|�p9��iL�.g����P>��i�ڪ`����/i*� ������H�+����]P!�k�6G�]�'"t�SX�<�4�������3��3d}�D��AtxО����BV�1�%(^%���kT&Vm舘{y��q(O��Sj�����xP+a����k_����4�$��|
�C�A�|*�N���8𛛞t���}�$ǎ���X%Q��3SF�5]z�B�i%l�)+����̏�j7[�V�ŧ�M~�uL�75�m��	�~1F��&W�����h���}�Ѯ��d+�G�����*�n�G����bD�n1��M�ͦ��(��������+̽'&��YF
2�sUng?`$��\������.�����ax\0;> 3�6�C�Y�A(��]��+���M�S���yY۵�q\H��EBF�r}f��ɝK�
-��a��#��^�n�a'dOM׻@���՘;;��Ecc��hgo��pl,��OA�`h�h����3y�Mx�w�,V*%�5f6�L&�p_20����ɋ�\H���R�&#p���W&�l������y��o�]Ĵ�~�Yn�/�{����^�G�ȋ��	����F*>�wV���.z߷�6��"]=Fz�;>8�bd��־�����T6�=\��iU"��)�m�����	km9�nF��e9 zC���������V��wf�
�Q�>,�^����ꁟ��)���l]���O2g=��;"�<�K��t�q�uR��y���Zk�AKHR'������#��V:�{�w�H��-�\�~~��c�K?�T`����A��b�Dz�h>�����b����Lդ`�k�BW�Xi�,1����g��o��,��Xm4wҘ�y�������aK�F�vu���)��}��"�g�߂����g�{�㢷���)���G;��(/Q]iZ���K���s�.>b�t&6�V���MB�y���ax�1���bef��W����7�]��Ph�Ո�72�|n�N�,n�?�L�{�H�zh��ܟ}��%e�{�9+�B9q�B@Ƕ�T�a%�9��=d֏��J���k4��};���3��	1��UBt=��}Qj�y�?���y��֖�x��˲oi�Ü��;���o���`'u����-���I��f��Վ�q���u M�=S�-��]�"pf��V %�����Ia�����n���xOď�$��p�Rd�� �ohT��ՠ**������M�Î|���-�T�/���a���Ղ��xUL��eĹ��j�|5���5�p�5L�e�Y1�G��.~v����~d���i�T��h��uٲ �����p�]�WQ_�����;��&n�rV�:�|�&��o��D�4Wfï�v�)�mǃ�
CC�U���n�����@��ևQ��ݴ �u.�y8�六����_Xy��N���S��ʂ���r
?����Z��72�*\���ܘ��u�X ��ִ�$���M��(< -,Q#B�h!������e	�[Q�#U��e��ӊ��b�]��x׊�x�G��f���D�۞O��Q��0����p�z�B�� �ޥ�«��ܓ�{����/o�J�|RF�~��L�N�&X�h��¸s.c���}�]ܓ�0Y����R_(L�ߒ\6հ����S/	~s�$3$�F�-������4��mZmDXod��<d,x3�~��<�:v*�l)�n����f?��qfRcN��Vl	'$K���V�p�ܞ-��moM�/Px?�٠�q���z]�0��K���.�O5s��̓f6�)�-@��k--|ٕ�(�y�`�*^���ĥnA�8j��!�L@���J��T)�Z�	^��#J���cE��O7$���&,'�*0s��f��z3�)��y>I�p3`	k����~�5�z� I��2u�����6���:�Sp ;��Y��S9^�goƒSXY�wz��h��.� �|���|��� ��E�gk��4�)�:���~bly�5oF���y_�DZ�� .�+�ɳE�5��hvN�?�Ӯm�C�W�(�G���2��2a�Y�K흼O�?��jFJ�GOG0΁u��e�����q�؎�2s�:@1.�*���%]L����I9�\G�H�Ivo f�al�(;[:�$�<��y�A�G�@=�f�4z4y�$��ꔺ+B� �䭂��ƃƫҘ���Y��C����D,�La�QE�)_=�&ƃ�/��V:.�۵!֏®b��H!>��`5ԫ�kz�� ц-$�j�FA/�@x�jM0�&6�\#�<��*?�4�-|.��db?��jYI�J�q�"t,knm����8z������Md<ȥ����p�4y����e�+A�3�TW��!�{�7����ܦ�^[��0�{'��^[�x5�x���ԋ�&��������1�i����vA!�#޴���J9K'�9���a��I�S��&I����r�;5�^J_l;�Q�F	�jO��}�0U��Mg��;��@��Lh�j��-)����J��P�]��wy#�^\�,ܦ��7$ŉC���1��!����ET����'B2�z���5m�'2�|�W��h0�m��6t#fjs��*.q˛��ZΊ�ڙ��ث���l}܈�u��u���1_T�.{�ΪUA=��w� �)erbۨ��5邖L�F�8$���=s�ט�S�v࣏�A�gX�AG�	d �&~�\[����5D�3/B��] {8#}�D��	 �� �݇΋�����3x��c��1���,ו��s_��hN\���e<��>d�-���9D\�2�b�MK�*���3�`RV3�Hh0�Jt��8�؎���	"y���^�7�s.�9VD�w�X�o3���%H vˮ>쉏8:+�_����3m>�i�qh=	��.X�\�F�f�+�!�/�=����]��\��T�����`Зl��c*=�4&hyw Y�A��Y��2*���J d�&^��4:�u�(���v������V¦���Z���Uq�
�_����)��4<��ACU�*|���Y,R|&fU~(Zbg2�8�FA5{+`D,m<a� H.j����	>X.X�Wn�p�-������B����FY?����x*G� ���4�G���Ģĕ��2'>�o]g#˹2g�Y�&u�RuMв�#�����ҵʿ5��DO��v��Ib|��N�V�,� ��d�S���������+
>���ؚ�CuR^���R�'�_�2�v%��Mv`�N�pƈ�1��D̇U��Ni����jjR���i������:�x�N!���(��Oze����-t��u�qG���["L8�;r�clwe��	��3�j���cRse����s�[�K���Rg�s%������u�2o)�ry��Td�G$��^��%��$�e��O�F�Q*���S�x��z5E���q%�ѲC��S��+�;���Z�.t���
�	�2S���:�>n���u��n�\ck���!fBV�t�;f�ou��޿�!s��8%M<߯��i��A�&lD黤S$��M����65U����#=�?��*�wz��p$l���Ż:K�k��/����	�ngT֭+�� �8Q�\��a�%y�&�Q>:?B١�X}�b�QI��FU�"嬈�85������TE����ؗ[XA:fPmeB����K�NC�^�]R�����)�$�m�9�3���T�:=�3�����ߋ���hX�� �������YCҔuX��n��	阅�0h!��Cu�ND�a�����������!;�Jo���t�j	���q ZM}��_O?�f�=�tp��15�ʥ� T�2ב�kb��]���<�;F�����\����;���m�q`�ZU���)d+�[�Մ��wǑ/��F�U�8H��
#b�nu&�x2�P~ߠ��t�%�u�?͵P���^pfs�/��<5�<ʦ��F��!F�x�5Htօ�l��"M)�nmĈ&�4꓌����:Ο��d7�C�}p|@F�S*|Y^0��l��&��5���,G��q��s�Xe�.���]�ʲ��)�5���@�:���_��]բ��Yo |���tQE���Թ ��=��v"�4}�K�@P'�x4 e�Z�q�}\��l݀LyL�E�!c�Na���)-Y����xe�A��]�Cn�Ѐ��pf������~�l�1cGs��U�;�X�a��
cӊ���A���&��w���	9�NF,�|Ypt�bU	~n�y(l��n��<��2x2��ٷ�!��n�����}Bp��{�ѯ��~	��;(V���)��yș
�:�\bW�͈���g�ȡ�4��GT��� ܅nj�w�r�_�x�7� �}!(��d��NW��DE�<���l�'Izh&e(c�V�|XE�z,���I4t�
���J��S �Ɗ�p�<�'��V�u��B)�b3��bM}b�~C�Q�v��},eHIѐ��B��rJ�y�����P��r��m���| �#y��^�ÔN7����n����<Mr֐I����e[�l.`���MTa�F���aGEޱ������՛�Ǐ{��ђ<�w�Oon),��4ܕ����`| �iI���W���D�<BA�v��1�kmGl��}�Y�E:���0��;����P����mv�QJMQ��f2��F��d��*\�8�.S>�u����b`���A�V�Շ�Y T�'�d=�w
*�`�7Q ��kvɹ�����B:��3�p�?
{Tk���]�� �;�wU"ɓ�8�g3+Y�Y�4��0�DY�=5�]H⁤.�	H���	:�Ļn�x�J��RU,��stN����C?���(��?b��1�Dk?����J��?�m��;FwM�
��
(�~ι���_�;����R�PE�x��v��v���$o����孻;����>8n5SR�e&Zzn�5�S���/�J\�:�3W��IV~�����
�K��H��:ʴ4����8�MN+AD�䏼����tK�r?�1?�������Ș�	����QrH7�pGN7�������rWnl~m��Ӆ\VN{} ������Ỹ��W�Y�s@�0�7q�R�������,>S=�r��t�bY���)�S{�ּ7C�8��h��Tύ���+ռ����ecX�N��h
��`�;�����?:���cW��g���
y��U�a!�\!6*�� �
 ���A�l�V�U�v{�r�:m�,(���#��C	T��`��M!TY�^+_�e����L[4��( ���cԚv,��ؖ߹���c5��(�ً
-k���ڏ����ÿ�eo�ș�"!2�J�~=5N;��c����ǵP|�UHܭE;�B}�q��D�ڹ�ا����T�(	g8��<�CTQނ��}�)�49Q^/L^Jp�b8��"C֕r评ߣ�����X�촐p���5�
ӧ�h��v��y��j���s�h�uf�4���de�P�߷��=S�	]��O�u�aCA�}���F��̔�������/*+L�%x�u
W��c���k�M�Ke��zc�jIw`C�:k��[�pg�$̨Y����IoTn=E��e_����`��c�lK�ޫo�%z�Ù 0��dw;?0��C##�{�`ɧw� �m����lK�;}g�m[[iar��cŮ�FA��t�r�3��v��~�w-�ۄ����zcM�@t_��T�~M��r7:Ur�h��w=�Ytu�;~[����O����&��� �����]x[����u��2kߞ���7���%�f_)�BF5�|-�De���"�-}�d��Ep��>1��C������ɻA5��t�.i<)��`�NU���0j�H4r�^��S�Ɵ��{�+06�7	�!N_�$4Ǒ��s�
M�
��ON�98Ɍ`KR�m�(��i�R#���D������k�̸�{[s+��-%.$�I���3��41LA�9�XG��O���A��{��bj3ySI=՜Z{I]�K�P��9�D�ե�Z�X���������Lh�CA�DK�0Y j��4'{�,�]�q���=1�z�&Mf1�.e�"/��i������\���;�qa
Q|���ίC�������7ȏ�?`]���.�[U�;E#�"��7D���w��:��l��R�D�tF	�1����y�^�{�;�!�*�1�I�#�@���N��G�@����ZӛQV�������;���eJ��i8���Q�#]�"|��䐑�ґ�@�{����ǥ�X��õ��gD���le�㥿�c��D���|t�	B��ZD�58����{u�>#m{�R�I)�OgPvX��$]`y���N��5D-:��m��2W�.,���Äy���]���8���������Oā��6�57X��Yѕ̕U%�c]n����v��*�EQ�@�'���[W�)���O��2��J蓘�Av�[�Y�[WuT�s�������R�;��p�V����rU�!c��?�d)`�ǆY��Q�����)?Q	`Q�,�zn·�Z+�M{`������2R�!	���x���x�h���M0qBzW�6��S�����^+ ����/wĶ�F�$ty
���)�=� �$��s���q,US�D�<�~*�P���{����j��(��8C�V�T{@�BQ���]�J�l`>����`�-#O��ϋU�'��@i7h�X΁M��%ݞ`,���o�'aM�z�f2��`rU�}�XJ�}$�n:^�dV��#���OY&8�R(��1���Ҽ���R+J��{ofWoq���Z�����S4ԙf��6#y�\^C����}�k���i^���B�j����1iK80*�⎫=9b���y��"	"��O�
�m`�j�&%s]
�G���H�D#��9��y1�5 ��\o;�D�k��_�Q)���]%,P������g�
���U���Ѥ;Z8��-�N���m=Bl�N�JA��W�U閎��0�3�	1�\tyѯ�#����5"�t�k<��Gq��3	 ����W��FL�N)������a��L��v��g4j�4Pϵ	ޅ�F�_��E�R�;�	�ZR��xT�~#���L����{g{�q�q���/�O˄����窬U�j��ּw� ��v���QUɭ���" �gz�^O�ὓ�5`F�PG�!&�[���$q0@�P��M�jDKխ�0d{l)&8�Ao��G/�v��w���ݲ�MHڔ������J��/�k_-%g�FI8�uic��ώ�j�,��dڠ��r��FN�Bwe~����e^���%�����`���Ɛ�i�ש��tp]o��N����4⽟�;a���&��1o�>_1z����}{������g"�dz�э?c*l\���A6�b�mX�ђ��љBDW�1�n#�����r���Q�Ä�E��5�^u�o$�x��̥DA?��h"��=G��7:#�d%[
��0rp��6�"�)\BԞM�մ�]�1���*� L��<�䠳�ѿA���shb:�џ��?5.I��B�*����B+K��R��8�\`L�=M9��:A����/Be�xM4l�6`W�ED0+�~=M4�R�=�����n{���6�༎����A���5;������Q�:�>�[_�D_�#�������MgMy��ܭF��\!�i9~u��ӓ�.IL1ɒd�ꉋ�b%ᑜӡ��W��P�ײȼW.�'֎T�<KCa����=b�2q��l��i]�w�C�y�y!����um΂���1�҇F�w�MĦ��;X�@#sbКd�
Y�t��A�y�.�r�up����DH���Fr��s���`�)i�2q�`���^�S[����\4C&"Զ�M���w#=i�o}������/�ξ+�1dv} �CV�P��/�>��~Q����RB���'%��1�a��
��˗'�IMM���8���:6��~��"��ax~	f���E)ɳ7e��X���r5���e��OU%S������9��4 iS�Q=�j� �r�kҳ��P�4����b�[C0���g�����[@�@�����v��o��,^'�)�m<k��*�W~��|r�� '�*��4���� e8�� �?a=�NLҊ��`�R�������|�$��@�x�vy!\F�V҉�OZv4�tc��_�W�JGg����f�� �i7�}��J�c[�+A�5'hf�x@�4����	vC==��������X�ݩU����9�8��u9 M��~t�2�%[L5���C��k̇$u��	�>�	#���o>�?5]���1F�����$!�����6��䫨�|we?X�yR�0�AM�3�	�Y�uĎBG���[�^
t�܉]�����2k�ִ����@�8���b|�g��AT/���j��k�4�(�@�*_��|зUU\��4��KB��c�J�+�Yf��:�_��rj"����lnގ�=��%�,Evc�I�#��O�}�E�܈�� [�D����Ve�?��Ԋ93�K���2����FA���j�����T�����.Ev�ˏ����{�|���l�S�^�U����H�����u z��U(}h��t�5Y�Ҁ�B˧}�)���d��F�[cJ	m����ks=��rk�t�`5-sP:$���)2�L'�j�؃s�4����/^���L�V��M���v�7�\�p*u�!��ٳ/9�̢G���}/}��yAŦHP�n�MȠ��'�\�����O��{{�9��3���/����Erɠ�|V2u��?��ec�c��Q7`T�o8��=��FXqЩQ� ���eJ��$�Z��Xu,ˏ�z\h�t�<�?e��U\��jkN/W:��"��ؘ��6Cү�exӪàv$k^�c_�үRe"�o�C��_U�6��C�ɽT�#/����qg�Υ�*VBv;9��2q�k,&��~a� ҽ8�a��s��'��0�	��8K:����&<���k\�����:�!�aN�8�&^����Ώ�����=�6�!P�\9���W�ݾ�9�K����u_��=<���������P8�ܔ�*
`�:��}0i)��p���w���G$�j��k���d1!�,B+��mc!Ok�
�4���H;�a=b<lҨ�_��Q^IM����ǎ	Fd9(���ADB_���l�Q=�G����`��Jx�����1�w������8���o�%,|�a1��Z�2�9��-.�6J>�pxsH�s�Ƕ:$�@6���ebd�wA�mV�:���uk�〬������f?0 9L>
��{��vr�����[[J��tK�`[SQ�nK�F��Ž�5t��鮪��n�~3��&�S^؏����
K���q �8�xT�b��!�N�ȼ���%MV�Lt�!��c�#�(��L�=�G�����'�ـ������l5,�����d2"$m��K>�:�8��2(��~Q��~�r�o�m,7�ȹ��['��NP.�����Hɠ���>����ԵK��:�>*sYհ���A����p�k�n�՚�j[���\� ��=� ��  l�(
n���JK5Cw	���3�7��}^��W&mH��&��E��#1�z���ZN���O����Y���
����qU�P�ĸ�:C������[,6��`��+�c 8���D[b��q�dy��ed��7
��1O[���9��l�[@�7�]
���[���Q��|�ܺ���3�Z�����_)�Y(Ӛ�?��&9�?���:݆�?Mv��+l���C��Zc��I�2{3NH��yk��I�^�,�	�`�W�sw�Օ�{!�,V��YM����IUW4V#�UF@�d��+�����w2�y�b�m�L'���/�q+��ĝuV�52�� ��{���m��H��gȋ�8�Z?C��8V�p6���O�2`�o���y��UO�/ĚӖjTT���oo��1`�:���H;���$�IM��d��2�G`ZQ���s�;.�p"�l/	�{6W��T*����Pf΃�)�|ˤ9h�:��󗊧���`�����
"�1��/Y��Z�g-�$I�k���ԝ�:˼ =�Z�V��|�I�$�M�d����a�S�J  �Q<v3Yُ]J�h�?�hߡR]I�Y��J0��v��k}:�N~zS��}\
�Ȅ4YD�gm�	q<g�p�g�=k6Cȵ ��U����_��E�I��C���B.8�/���mh���i����Z�a�_�
�-�����ƪ��g�,'q�R��YK�ca�x9
3�/C�	��L��A)�P���~fm�[pO0l�?��7��1mWN`���)9e��;��������Z��q��x �*�З�%x%80SS����'Gu9[4x-$�=�Ā['�������jK☰ֽ��}��7X�10H��X)�sU�����gAT�>����D��E:�#�����k+���P�q�Y��ǿ&��E�1�o�+==������3�Rw��ڹ����}xY��͕7"���e�{�[�)�B���.&-ѱ�&ùc Z~i�,{P�W:R���6�S��=~���� .��{�y��,�0�5%˗�����X!`1�#c��k�Z��?�������_�P�8{P�r�rj�׀��5�~sq���z�T�Y̋���e6c�xz$Eҏr,� U��7YrP��+�3��W�������&ܸ�*� ��椊�=>]lVM~��yg�V������TήFs�-�r��E�>Ǎڍ�M�,t8�Z�`��gо bI��a^�����*eu}���.G��4�H��0���NU��0�� <�>[}��Uӓ���6U��;����+���U6{.�"��vߔH`m-�������:3���˙IG�|[N
���ԕ���s������}x�e ����dϘpyl4}u����9��x������t?q����V>�T��
��]_�⢞��ٶ���+�H�-EG+��e�1"��*��b�+qm��S�4��f�~��=l^�������b��~��j��n�5OSW��8�lk�NR�_�\6+h��"�+?z�[N��+��9_
Z���_o��n�5W�as;�����;~�̣��𒤩{�o��9N�<�Q��!����Rs�����R�XM~�1��b���9��Ti�'w�MH��cm;��n��\p�%�"//lR}0=k^h,��^Hu��l�[���d�&R��Ѹ+�<��^PB�$E��#���F&�'إ0?0Lyd��Sd����Zai��c�ϭ�8�I�p	���Ԍ�M v�����f]ݏ��]�Ƞ�0�ٚ��
�; !4g2^?����h�w �����eS�I2b�0$b
�����}�J�e�u2ww|�7^����[q��~කSR ����)��c�o�;y������;�7��p���c�a��3+�w��L��In�a�rbTVq���U�*IS�d��g��JBf�)��k�d�Sư� ���k�(�����Ⱦ,�?�R�(l,u�q�����\���
v_����؂E
Mnh�OO��^1Ep�S�%�^�C�ԗ��<b�cy��.��F��2+�J;׊4��H��Wuv=HZ��q�"���X:o1�pPWH����j�/B���̯m'�CY�tg���eLO'(��X�2�_�r�����)�e�"I�s�ue��2�+qO0Y��:ZQ�4�s�,��U2MӁ���&�ϔPr�= �I�"ቜ�yBR���*ԙ9z�� �����eU�u�{�/
�UB�J��9M86i[�~`T���uzӥ[O����:f&UM�9ٚ��(%� �TƄ�(�����V���fQp��0�9T6�p�}0�H=�4����f�7�	��f:dD��1�����I��2�����p^���K)�I2�\]�?��b=Qdb9��h#�n��CT��\y�G���X����Z�OM!�$	-�v:֝2��T(=�I�3�>��?o�OKm�{����<C"�U/.=-�ûeB�-j嘢h'��!p8kU"����ze6�ߕ�HHP(��?4�cK�A I�<~��	�_u�	��?�r�S�*��rY�����X�)�d��F՚��K"Z��
6���5����@|@��1��/�l�t�Aa���A� ���5�0�c��/����"p��5�5�!f�"��6H3ӖVE���&��
�Y��C^F3/���L_oX�o����mM��}���@��\U��L�g�7���j���_���;c}�l+���Eħ�Ծl��X$��&���8�_�Ʃ ��ZJ��O��*ϱ1�Kf���f�;#��1�i�aS���L�BQc=�<y�̕�Ρ��04scݒ����T�MU���<jW�ط|o��/X!G���r]�#5�!Y ?����e�ZZv�!Oz�GJ�ネ�z�+AΙE�Gz	+̬�@���}�����籐��㈶
�2�E�A����Ҿ�Yj_"[qV���g��;���M;����y2�H�{�_�u��Hn���z��d?�N-��
ч���)�G@�0��5j�{��ǉg"��2��߮p[p|�6ȉ�HRj�-�R��_���gs�� ���ꢁ�x�/�C`d�N~�92&��F��ll�}���K5I�퓞û��pMЄG�ȓ�Ip�xz�"I�S���Z@��=E��FQ����L.����֙W��*Z$ɸ]v����!��ʦ�H]�ׅ�^N�Ul�/��s�F��&��=��o�_��>��Q�<�'��P�i+Ⓩ��W#�[L!�L~{��� V}X���.�� @i��n���E�o¿"R �Jvu3'T����p�c��c����d��sZ�ZA=$��L��h�9J,4��z�{eA��È�/�����F@�ǽ��\�$���e !����S�J���l�D�ط��0:��po��G��� n��{10a�6d�X!��xx[W3���YΓ7�[ޏ����E��c�sC��)�`Q�'�L���9T�
/�8'�
n���L�M��5���i��������5����K����P2�̬�ۃh7>3�	ݼf��3 �����m��r�:@�D��Xu�wN��4�dv%m��k�^��m>�} ��A�̓*�*��a���/P�\^blB���W}��.�*V���`#��B�9{�uЖ�� 
ߚ�̑Wo� "S.=]TiX��jm3�U"*�]l�v�~֋��Q�8� K�Λ�R�e#�n y;C+����y��S-\Ӟ4��g��8n��(7+GTOgF�.�@����!��� w�h�|4����