��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��X[&-����v|��y������S(�o�o�r�y�����l	��x7	}8؞��ZBg:��RX�]�+�2"�쐉@.��o���kH��h@��'␨�����$k}����\�K��O�n� W�t��J6�i������|;i��@D�>.vܸU0RA�I���Vh��et������u�IOu9������3�'��&b���|R�Tw�?R���JR�,K��8i{ѵ���T@p7�RH�ڙh��NZ��7��H�&@�6��߈;� gS�1,%Y�K �C�@���!]vo�����1���rH�5 �G}D���5W��@�4�d�6$�����.�렏�l�	{e�!uk�������0�u�������Vd�Uy*[�7:(�0��B���.˂VqDigQ�x�����.S >��V�IL��� H#�2]�gnA��ǉT`4`�o�}�*�aܢ4��z�C��Г)αQ���	I��>��v�b%�x���d�����{�ym�6���2�X�F�~qn�t�G���ʷH�)k�U:��Ugi�0F[K?��<փng�g�'�XQz��$�C;�<щ{O��)�ٿqh�ds�����@�!q⻃�����e�g��-{����n��%����2�g|��S��gmn��qr���`/��Rc+?7�6�I���A,�)��!���IR�i�bb0Or6��5�ɣ�:y��foC�����0r]�d{�I�u�P��#�SC�҉��cN�&�`#�Y�҂55��C�*zvO䪊]ڭf,U�ifD�rP�`��}��9g�Ǹ�I��[h�����I��C��L�2��l�$b�4,VF�9��/1Q+�x�'�݈=}j_������֓�M��(��BЁ�A�B�J41��A�]�n=���5���pk����]�ؖ��9�_�K�d�>Z1k_�#�&́�~+9�je���
�-�G����=�ny�:��Q� ��8�����[̩��)J���nN#u��b'�=�\��εd���r�h�p���LN�r�ൔH������0�Įr[[-k]jͨ�w�ɪ��"���{#��o��1i���]���|�h+�Z�Oz܌6!� �z$�>�w.���ćY�����j���&��oVr񨗂�r��*��?�;l��Msk�!���=�����s\�0�4��h�$rqEˑ��>�䴝���=F�����D���&�pi�U-B+\�4�/-Ue6�����YD^�Y/}9dR/.��z�����Ir;�UۼwX5��3[Z��u�&�ً�k�!�Ǣ��O:����xA��@)7�[�	���!��ol�+� ��)[���V��2�tn��q��\�6Έ̿�U��a����l�� l��j � ��kt���Ak{�N	�!z���-+K[6����\�v��kk)+k4 *E��]0j��/<��0��J oVI���;�|Ħ	�%��B
�'G�4OS��9d��;�����7���1L ����n��Щ^�� �L�q���"I�m�Ae!�Ĕ�7ȋ��j~���N]Y-L=� ���TPY*Y�jȥv Ե3$�ψ�CE�)�6>�҅�~� ��f����R>��EO�ϊ��$̦ �h��F�l �g� ��@SVu� �sv;�<y���	��˂�����xڳ�[�mo������w�?�r��!�i>����]��DYBAɞ���>�������iJW���GYW0��Ʀ/�"$aK�a��\oޥ�{�z�w���1ievP,eD��*�~PB�71FS�@Fs9�mBX&=��<�$+�oa�����*o�9����O����^!,�n��3�[^q�N��X�L����̱-�>���:YT{�.V��A��Yj̧6j!�Í�x��� B��وZ
�CNΏs���ԭ�ܜ����Hץ�'�.&� ����E8�POgDy�\b���ãY�˘H}�i�g���>M���J{��U�LA2��#
��^ߐ��&��
�(�����)?�� �(ecUj�u*W�=z>dS3���~8�;xhs�̿���^���������K�HC9����<b?�}�z���v���#�*މ����+؈���1�磤�q��Ѐ���LKM�\�k�T#�t�,�)�aT~���'	@o�5�m>8 `cP ڥ��S;ByZK���T;�A5X�B�Ij�ͭ�z���av��7x�1U?e�;p��CM�1g�p8c�m;�V��^����Qy�՞�uc��Ľ�J�UlV͘�1^~<:�sU�Z�a�S�j1̔b�Qv�X���a�|%�E� ��,�O��h�k�l�����%k��=�{�j��oo��O���a�eE�A�E"0� ���!�����1��8�12�C��'��73O���4��&KK� ��C1*a�3zDՅ�X=��r!�"=KoPo�UE���h���7A����L��-rC3힍�û�`��!$qlx�+�|��Hw�&��X�9�����%�J��V�H�Ե����@��u��G �gτ
�>�t��C+؂��^Q�����%��x�5������=��=-�|U\qw-ou]���Z�jv���*��I�U^��#�Y����l�z�F����������|�דq��O��UQ�	��+�l~ZZ�)"嘀��E������ۓ��$���r����sa�*�9--�Y�@��k��*�.�#��r��y�äZ�v��d8X��8U<1�a1���K����Չy���qi?�e(s�vr����+�_��`��3;rUmq=2̽bq�j�l�a(��o���@[�>�ijJ<�d���#�z5����8� _���xt�kL[|\C]<(i;X��m�^�P��m�A{?�7V8�Nөh |F%��Q�����Hp��D&D�ii�����j�G�M�,z5E!r�Hpݖ�)o�w��_-Y�U��ѣ���!���^��Cw,��kMpӎR¼��(���`��Lk����g�+AB���֢4�3�A�b�:�䪢.�,_S�ٻ���9`�|��\bq.6?�<�� ������B�~�c���?<��w<&�T�,;�!�^&��q�A�: �Pɭ��wp�1b�w�@B6�~(��)�8�[��#	�"��--4ߨRS6ǃ�h'��I/���5E�	HB�UF�%�fc�R� �0��zU�Z<)�'��'?)PZ)��shHE�T�(\�-U� *N�-(��M]�9� e�@�ܰ]�פnQ4&��\�OT�j�3K�.�y_zR8���FA'0<w�mz?���j���	`aD�Ӿ>�c�ޯa�Y�uojW1�;> �Ԉ��X���i��ؽ��d��/�bu���G� �����X3m�
"�,���k��~ӹZ�v���>WL6-=d�p��<P1ӯz.Yܮ��;@��0�h����J"lA*�-P��lא9���`�$9@��G�W��;.MLٍ.�[�Ws�����HH~氋�?)�e�&��c�*#s_tY��Uj�,q���S#�
z��\ETvP��MlP1�^�����SR�'k���v�K�1FY����RȤ���b�8bB��/���,w��$^����TU��tB]�콆�EG~�K���P9}�B��K�٬��\����v�RN��I�NҘbYPq�	u�=�y��A��j�+��c�o�~���vl6X�GW�����~�5����t��{��H��HN1�C9�/57#c�m&��l��j�E�R|�=  E�H��ЅIe��:��p��I&��N�r@@���<�C�8i쪱,1@-��ʛ��^���ݝ�y/ס�_�.�U2M�3�3�X���j5�7����=US��^��ؠ�1��g����T���(�"�R׋�r��'Z&��1�#ؕX<���2#K*��6����ݗ`_'��P�U���$������I�ʺ�q�"�̪ߠ!���ꀞ62�20mNbrݙ	u[
7�z5½-bT���寇�5dD� ݹ�u\սn��g��d�?5=a��w�[ٯ�QpxvOz:����[�ng|�l\�0�_@/6M	��|��'�,� (g56�Ȭ�Z�@N<̠�Wk��@(����ÿ��0ґ�0��@=��e��;��;.6����-Ie
@�3�C�Jqʩ��� ��'��1a�ag2�F9�(���E?�ĥ�h�$���f��5C�t��<ko�j�)��}�����3l���/����(�7+�����C�C��,�e�AS�笟�"�J{F�]�o�Q�N�J�i�V�J��Z��25�zi��7��C��Xr#$�B0����Ģw���
�������;��Np�Z�J�?���c�P����T./��(���a�k󓙢�rIl"��#��TNL3��t<��wy��l�����e���aS����� ���0E����n�2�8XW�rk3�^�1���W#��5x$;vg��K	oD�ؿ	�^��0�c�I���`<�Iv�jЦvв$y���.�/1u0�����l��,�+���0�m���&�H3V2��DH5�����L�A�DD�r?L2ˏ��L�lu�[s���fJ?N8G�{��Ű?P˘&4]7��-κu��Sh-�G2X�b����4�C��Ou��s;�M!>/xG һaqs�S�h�C
�8�����BJa���`r&8�i��J��#T}#��Hon�dW<|���έs\m���cU�^��>��>Qh^d��P(R�(�������͎J�����K�M@�դL��V �0��7  �-n�S��[���zi�G;�V����4�����tQ(��p�g�'��Iӥ�4q���"�l�Io�	��`���ʍ��z)"c*��U��#0fV�f�,��e��[��c2�n��Η��*0�k����:a�,)���0;�-:��J�R����� �RKq���	�J����fTL�u��̅��ͅ��$��N�g�5�m/<����B���I��8n�����a��B��/oGPd�]�빩H�wz#*wSf���A�:@˱�S,�pm��e�y�"b�f@��']����Z���VB�^0�_6�ju��
�	ފ�9g\;��A~7r�V��Vݑ��pЋ�T���'������yf��ʗX�cx'n��N�o3��:�N�����-j��`23�Ș�牘�V�2Y��jpq��q���4�aA�#�e�� ڒ.'׃�i�m��2���68q�aK*3��Z�l-Z�:�fcp�C�01:�ſ�B�	j�'��u9��ka9-������S�e����c`I��!y0����23�K4%=�mH�1�"�)~ ��@���齢��>�'h�o�DE��Vwq�k���� 0n��O���t�P�(.���@��k#��[�b ?�pw����;�*C^=VaA����\h�?�/夽U~�0%*��i����BQ4���HU�	�� �e�Ga�� ���*;��j#����H��،�5\w�!I'/��G�j	�]v<�����¾�h��k�C����-��Iq���	���q�@�	��B֣QV�������`�a�X��/) r��>5��m���h&�J$5s�>e�)��,�񒣓Yn��TI�bԉ�wW}�qm��P�"�2�Գ:�Q���c�F����߄㿌��R��/��Tq�W�]�|ջolSN��!I�<s�d����U���"�@A�'���!�S��Rur0o�{� IS뜾QW�c/Mő�Ցf�V���ڕ<���f6���g�\7-	����}$o���{���v��5[���/�ҏ������Ik�G��H����.�q����ڍk*�mRA2�tY��l��g8�Fr���p��z]�.B%|��iW�*QN�?@��;����c�'���HO�5^�� yT����[� G�a@���짓us���(��\k�6��;|ʢ)�
M"�e�(��U�v��*V7���X��0Ҟ��d,�ϡ�
,d2�b�gt@���3��U���Y�}�<�z��NT��H,����u:u��v����	`Щ��T��k��Ww���h�!B^"h��}���qa�i�\�g��2�V� H9S�X�����*�Η�����
l1�.�t=	RS�RY��	&�8�5���;�	�����Zg(�B��;�����rM%��m�9�ĳXMʋ�g|w��n���/%�̦�ʪ�Tc&����"��`d q��G��$�f	J��ۀt#2&��1z&<�f�Zh	���|Y���.���=L�s����0D�K�}߹/,"zp��G�3�Y����6z����,.���x�퀮sG&���$�ۈ���4�u��cc��*|��eg�;�(�I��J�e��5�wf�"�;vK�5�����)�Z\�g���q��^�K���ݏ����E6.�K������}�붉,�eYi�_A�d+���Ȼ�e���C��rȏ���� �֠Ԝ-y^����"��I�%���E�
1��!�s�q��n��1;�Ґ�yV�r"v�jvƷD�	M;���!E��D���d�2ç]B�HJ�( ��;"+��v��0k�����.�G�A��m(PbEI��z�)�������Ɏ�A�8P�9��%޸��3%���ȣ
{G������aUվ���8���b����^Wɹ C�}����z��;b�4�$Hܸ1b��/�XHS�M\2j5�d2$�׵�pb�f�bC���4�� &��ѓ_�,z�>|t�w���`A^�
�
Չ�ż��P�mo� f��iĳqU��q�XGX��\�/}J���:K�p.a�r*�{y��':�s7S�T�o��l< i��_�U�Ci���n26�X �j�F\�=��J�/��|]�����S�|��h��e`���� �.�b"��%������1�m5=�O9�^�S�cY��bY��*��v�p_����f*۳(#�?�L�ۤ����@�(Nw)r�#�	�~['�灒�J��Z��3$�N�kN��S� �/$AL�:��=�d��hӑ�,�0�n �{�L�Ԓ�\WV^�Fc@-�
�̗*��%�%˫�ɼ�q�S"�ĺx&~̽
Jy����I��G`��m��%���9%>=J2�TG$�����ECч�h�R�p.�^f�~�Jː�JB����?vy|�E��F)�!�����x�˃�E���-Ͽ�k;�5O踘�hwڏ�>������	��+[n��L����<C6�)к,#�[p���S�(s*��1��e���\�i��#!��,L&2�q�	�O%�4�
{e����ͼ�?���y�J5��x���#���9��|@Ze��]T�~M7٫@0������p��Z ?���+uv	\�E
k���,T�Es���c\].����P�;�4��0�D�~0%(�������I�4���6&�?��d���d��+۸��A��m��o�F�O�HYd�1��b��n#.��[�A���9^�
�`k��5}2"W�����[%k�^:况���W����}�sz���c>��Y�ȓ�>Y�&j Q�����C��_ ~�♋��p�����.�.3��8��<;��5΋F�m?����<���Nz��I���cY�&S�=�Q�����=��j���DG��7�K�41�vj�p"�I��^(��N�f���"A�(�֦�p�P��c\����td����Z���I"α0sQz���Q���H���;
C��p>�w�+�3z����p�_��{��W���`�#�td=�#j��^{h�'&�~h��i��y}��U��������A�I�R��~���ܒ$+İu�˳$�	d�+����}����/�r��Б� �P��@������}��{+���	���G̟�S�C��l�����
ַ��þյ�U�J�R�cz�p���rrܐ[�'��p�~�m5^^nun�Rd�͔-���R'h�����>��%�`����m��!���9��JOHAZ	J�ϟXђ���x�[��G�	�6�����*)�DH�(���>�Q1��Z�]a�����v��T����ԉF�"X�C���lq�@�(����:�̺�榱�2�㺡_r�5���k"�088������2p�M��t>�B>�ս�f�/�%�= �q�]�it���D�|a)z�xt���2Ɛ�9I<X��&:�����!0^��EE@� l�,���Ǡٰ��[I�z��q֤���i���6�0�F���&�=u�!�@B}�*Hb��tF!�1m�	�3�
kUҖ��A(|�L�cp���L�_��R��QfT�%�NJ#�n�"��:
*���r�
�2u̕?jϜ��MW$�u}A�G�l���ﻝ/�����b���G�laa9�I/�H��W4�V(����%�����B�����2�D[�%�b��%;�PO��%��JS�@y���>?��=�g�Bg���fo/��Sj�����kp�Ҏ@0*���!�����������{rT�E������?�M�\�B�L�곳�aj.c�1/^����
��b�p��"]ԵjH �s�Dx��	u8��"�;Y%$v�����8����QM�T]�
���ҭ�����d_�/6�U������ ������C�%h�)�TEwxs���Τ��;�R�A�B����d�!SP��\�����k�.t� _�A�p�e�f�,i��4r2�zOX���h�mw)��(�rr���<~��d�߆���7q���m��oo��-
��.U�?&��.�z�]�$�>�2�(�~����'�W�B������=�1��.G����SЌ����7�A��:KA��XF�����E���n�@�|�c��y�ɬ�PQ���|҄�1YX�jX/�:�r!�l��} �p�h/�|��a!� �FT�^�<Ư�^I�fn�<�W2��%Ηmsxf�##�q�ǕܒK�&�'΁fȠ�.���D�p�L�4l�n#���z�D��O㑿*�<�S�唓�x�p�,؏
���SLw9�#+���b���[�6�J�*�=����q�^�)�RI�Gh�?�{�D��_�F q��)��h���\f2�E�$�K���.�ߊ���}%��m�E��%N��}�Nֶ#������u@�G����ek�c������A���k�(���|	��p��Aœ�č��	����U9^���!��*�ku�8i���Cw^HZ�Ї���g_�a���Uha*�"������"�c;�Yي;}�e`:]{n�;��\:�:)-ЮWU���M<���xN���mo���5g�0���*_����A�1%���ǉT��e�,yS<���개�������K���!)nk�P��ނ�E�F���,���t`��v
٭�S���鸤�/���rƓS}X���+0��#����5����oJ�W�`�T���˵�(ܗ�zZ��!?�(�<R@�q�� ��� ��!Li��� \�I.�4�-��f�h�]W 99척-��e�g:�c	����`A�Y��qzb�2e̹�|�C(~��+61�f&(��t�|,;~IBQ�{ٷ����늄���/���b�`���O8Roפ݄�]y�m\�Y=W�cʑ- ��W�o�A�7��䛒	����Sw#y�2�;�������n �G�T�.�����y�$x;�u�@�2�fZM�~�D���2<<�;��b�F�U��=�@�W|��Χ�8;����'N�����v��v�:6薨,�9:@@4�n^X�ڠ2y(!(�t�m����V�D`���#l�_�'��$�����̗n͔*E��������&�s�)G�/���^w�Uac!(�tN��o���e��&U'������Cw'pB=[1��pӧ��?��$�.5�e�}��['�H��ɪ��°�5�Q��{5SJ����g���њ�[W��=�ٔ��N�	�ʒqh���d�\6�+�6��M�m!�/pɗ8�i�+ݍ�'wv�Lj��"6i���n�X�j����nQ9�K��uH[:�sb�V�`vm�kkl�X�^�>Ca4o]��>��ȸ��J{����:cp-�)�9�M�=Oi&5 ���l�M��a��X����>�"{(��� �[+J&�r�J$[���6P)������@Ҭ�/�Sr.��rQ� ,tu�^�$�-� >)��bU���<�Z3(���2G�0�^7�&�������r^�U�!j�ϕ�1���о�8*�7�L%�x�
��t������vS+U6���봨vU�?���.��'}8߂Akع3�t��J��b�	)H�P������
5�4���:�%乫�->�<u�g?�Y��)����u��]�H�lk�Ay�{������7�Z��0Ţ&9�
���y��	V�� Aa,��	DU-�/�r�I�ª%b]E�b��Vd����f9\7�Ȏf=����V�0"d�0���L�X\-��t�P2���q��,tm���3�e ��R����_�JU��*�������Nxjv�T��g�'6S�8���#`[@�[�(�К�vY���[��|�"��v��T��B]c�2[|[�Qoنz�U_#'�P�U���/S6��V
�Z�`���`f��O��Ӈ�:���r����0}�JTz����T�4 @�����4�Ŀ��ڣ�k[�s\�e�S� �m�K^�ͨ��s���:���JR(_�X�SN|�,O
�*PĔ�4�I���p's1zҋ�)ʌ��4��DG�	��fD��E��~ܧdÒ���g��{&���s�	���� �UuB���y������V5ˎ��j�#��JV���.û����:�z�
D>�ocЬ�5�+�0DR?nr*, �j�������\p݈*VEHP�g�.��<d�0�
@����+���T>��=��P��7z��X�2+)�"c�1$��uk�h^�I|E!�ir�a�&�$!�i�w�s~Ӹ�r�������V#:�	�|�-��n��G�[{�� ��[9�������P@�kנ�z�T"�)P���^Z?�\H>]�țYl�I[��Jl8�R��fk��"�W")i��U�����1a�	��}b,�>��ˎ�q8{Ä����)0+Ti#i�=Bp��g�p�N[4��>z<K�m�i������k[�DR��u�>�D��t�{��8�!xsa�Z,V�Sq6Z���yL�s�Jڈ��)s��R9-ɝ��������_^��8Ћ竾V�\�i̵xx��n�0�pE�3�ݥ���}ѹLN�g#[`7������8cML+���e�GI}0P���v��{��w/��ݕ^�2�������gj+,ŨK&�/���P�J����c�#�����
��'T�}�8tN���>��i�-��®�]J��m 3�P�V$�r�"ؗ'���C��Y�����C�(�de5�V�և�7�1�8�B�THX�p��J�nݢ���R,#�uDq��Bh���AL�}S�rS�폊1��ס���ݾ�z˭�+����z����~�hK����}��)ڠ�V���%5;�>��!L�U�$[)�?� Ei��?�Fkm�/E<����^��;R�;� kKU
.�Kg��R��'�7�(�D�V���=K8�.��E&�\�
A�-��A�ʊ�&���i�}��uR�#��U� 0.���lp��Ŏ�#�{�L��Z*.�ct�b�����c����T�ժ�{%�z?�c�XH�۠���\��E�ជ���
Ug��'�R�U�>!b����:����l{f��Đ�l��|��j��Gb�h-�W�N�p?;n1o�\��h�M=�5@x;���$���a@��߈j��jo���R��)�i���!CN˶!�2W�5�t�~Ѯ��z�V*��U������v�u��t_4*8u�d��,�D����{�){�=�	,W���ʮ�c��=�iS��ݙ�̥>p]4VڈzT��Bw����ŷ��́w��i�[�v��d��^��碁��X(a1G�/�	M�iԁ��[�e��v^�:>7b[��Z0N3S"���5���BR2�f�*��Dd���7�^;�t9R_	��vaz\Po�)�ݐ��k2_�
�3��*�L��؊:g��{]��@Yä�5ȵŋ�;��`VlH`t��.�$�BY�};��q��g��U���"3� ̌ͧ�^��
2|~G��M�н�[��������ި�I<饬�ei~��ip5�1:��B��}�Z�c �g4<��Π'Ux�� 6�S<t�t�
�B��7�+�F�%l{Y?f��Dq�S�������l��Ay�ۤ|�.���C�����&���u�r@�x�;���M��e.������Rʰh­��4�H³��8�T	�� ���(Jp0��(���;�c�r�PKS1(��{���`�@D�*���}Wh���ު���({B�o$	��O24�b(���P:o�$Q��
��F
a�T�Cڐ�s�ޛܕ ӫ�<3�;���p��\�4�LRɬ�2��3a��Eݪ�ϒwwAHkؤ���q�I��b�c%�(�bg���Z�ےS�\�#B�)=%F*:�	�Rq����N>�)��ս��6�-V�2����o�5�QLn��V�Ң�o�\R���h+c�7�K1Yz������#�3�a�5������I7��۩l��v�Hd�r�o��8���UM�{��̃ ���os��ੑ6��<nd�"�����w�[=#�}�_�e&�aG!Pg�[�s ��X#J=�p��"(�e3� �m.T��Y<�����,���[�tK��$�T7��[Ś�ynCB�z�ge��s������'���w�J�A[߷d^V,�ϯl9Y��`9���v���8m��6X-��e�3R�<�<�U��B����q����l�J�_����VC��~>�|0�mq
�b�k�ɒ��f4�	�T�犯�VU���w������p |�?j�߼]>b�v�g⢟�������sC�@�8��}��W/����D�b����眮��%��H�jc�5QV#`����9�*��u���s㜅{t� �\��pi�~}Ǜ���Jb/W�~�a�)�l��5��n���i�κL�d5kU}8��Xۘ	���bͅ�_�Ws|ND���8��r2T�궳!��!2@�6��u��wU���i�c2�e��[��K�x"`D�t�n���,�q%�[�/B�&nS�lW�ź��e!dgv�R���s3O6
)�->�)�?�ۡ�}���M����`X�M?~T0xO.��F�o���Wc��!���4���gQ3
D�<s�j���i�X˃ �Q�"?�gQ�
�D͵���8�%e�A7�{Hx��у��.7�{8�3�ՠ<Xj�?���`�D�
K
,�!]A����\ϕ�\^ �z͑3�^�����7�j��Sݬ������t�	�;�����:�����������J�iZ�_xI�����
�z��H��XIf
�ʙ;�"�S��.ǖ��i�^zSٽ�C�}�*"�zu 'v��EVK����b��2`|�����Mp "��Q`��xl� #�xww����'�L�e�@/L�%"��>�a�ǜ�w{�k�3�I�dlX���~C�$U��sV��Iܢ���+�'Bg��h+�G���R	jD���.���7�3eci�p���������l����s�hmc�ҿ��4��=E����#"�������,L	��@�DP��݃S,����B^ؗ`4ȶ�nS)��2z@��M���_�eI�l�H�����ɞ䛄��k����\������X�3&���%,���1�c�}��3�~�w�5��U�a���p��ʍR�З$�� ��v�π�F��`����,�Ń ��8���c�4RWbsvh��	��̻����B�KH�p�&��i�}G}��<��J�0M�㫔ÌwyLW���$`֔A�����E8�X ��$��H	rR_�i���V��:��ȳ������/���9�C[�My�a�{�QZ
*�lʊ�yО�0[�n@�-�:R�h��Xz�I(�"�RNǣ*ꖰ�F��|���L�n3�T�|��m�4�P}��e��8���oY�(*K�M��f�UiSq�1WR���H�?�I�k[<��t&�_�}�jݡA�=OmmŐBw!M��^��Dv��N4e/�<U�q54un��r(���?x���x��F�ɓ,��i�)�J�h��\&D�ծ�B�L�=��̗��n�Dÿ�;�$�c/��s�)RO�3�w�"%�=�r8�bT\�v�-Q_Ba.3y����|aHb�iA�bʠ+���o�ٰs��]� �rρ��Ϭ�O|qɲt�:��V�H��D�[��T��z��\����lȏ�4�X���M���f�*��-	�`�3[�w������*�6B�&�:Mꁋ�J�k���Շ�t��y�&;(����.}1�!���k"w=K �l���Z'���Gj �(�x2/u�6���-�[>�ޢi�Ȋ L�� ԹK�2�S��`י�oM���3�ao����U��ׁ�rp���zpZp�!��q�[�U��.�m^�$��v`H93V��X�$�(�tN؁�V�������������da�h�w�Ob��Cw{	����#��4�����3�jf��'��t`ج�g���P6��!�=ɬ<��l��9ʉ����(g}�i��:"�����ђ/�q��^uus�Q�L�J�u�cg�#�����7�;�إMfh-�*@K�^j��:�"�.n���oUw���4x�?�D�H���nOH����f`/�\K�:ksXkxV
����Va+CY�CO���;sg������2(kʕmYlY�o4ː)!8���$��sK��ꌕ�>��������_�������Z�re����%Dћ��Z	�r�#W֓~��g�5��D2"�]"Z����n�sb9AQ���\e(������OK�(`w��8�Le^�{'wO7�u.q����4��Q���VkUܨ�l�G����&��R���	�$)([�$]�����4YG��k��i�#'UԆ!���0��OO�=>q�:=]��<�b����r3wVe�f�j�?l�'|g�`9�e����+��.����vE!F�;o۰��Df�p�&iA��&��jV���=��P>��
��bE4$���*�S�����\,�|b��aGS j��8�֋[�8<�¼:��.�2���dD����k�L�ܤ-���;�R�a9~�{;���0�H�?d:�,�ض����6��[;�F��X��D�^��I%��⢕��a���N�2�x�-�#\ 3ѫ���K��Q	v�&�L��jӱ�ɏ�>�1�@�iиsh�M}x��X���g���K��fd��Q.��dþ�E5��7��@��^NZ�X�:W
��/r�35�����X>1����	^a��!��@L���5�i���is:��u���ՙ�����3�qR����wJP*�n�N1be�#����8�lg�0�G�dw�R@^� ZQtQʺ��a��]$C)���`�¹Y�ǐ!7�tv�"˙�?&)���n�kX�,Z��T���b�K�{���%K�S���.t��8D(%�u��v`[�zl!a�`\�Ȏ�ɮ��A��I[�b��>(6�-b�єx%���y�uu��)S���� `[G<���J�@��zr��h?�Vċ{D��sj�*�����|rytq���	?��*�i�y��}��pMpAr1�P����U����E�\�߾��PP5�M@z�ԅ�g�pG�G>󀜀 a;���E��+I𶊟ʹh�Q��~@��ō���f䮋/���E8<i�.�6�/)�x�G�C� P�u5��wN��[�lN�{o�4��F�/�4F;�T�I9������xM����|���[�`ITD��y�Il`��"�x�u��IBɿ2�w��H=�nv��:��5�  ���s�Z:���#Iw9���>�n��+�8�s����m ��:�L8_�)<e�VX�f��Z4�<5��K�>�.��� t���祁[K�~Ld�:����jcaQO�[���`k�~��A��`�\ӉhF$���%�q��M��u�9��J����<Q�j5�qJ��`�I1�S�&�	j�F�+~��6t����-ӯ�O~9 ��{��{��h�H���͝u����Bb�Ǩ ��VIe��^��G�%����U=�DE��yN��"��
t��Jm��c�ٿ3�N�˓=�t�$!�E��D��^����s�nQ>������H{�u�$���X���X1{fa!����:nd�%QU(gk�H�����3e��K���X�E�c�
��d�w鞭n�(����ŵ~l;LPr��������/L�ȗ����?O�p�>m;��T5��jEt�X��5�-�:G�m��Y*�)�[I�%K~��6�#�aO)d��r��R����9�pk�>U��y�&��BZr8MbO�ȸ�w�=���T�;���>�ڷ���(ݶz\��4�p�8��ҹ�G_O|�o	3;��Ǜ�����0��gM���S�4O��|��^_"~S+��*��Y�R}�ɾ�p�T���2��02X���Yr:T�%���E���E�� ��ֹg[��M��/�V"����٘e�w,u���]ᆂr�'��G<�g$%����cK��N��v��Y�+�9hYmк�d��\�&��%�\��Wt�T�!�\)�=B�B�l�5��=�5%%���?4�L3��P9Ԋ�YRS�a����������to1�P�8c�Qzd���cF�x�÷��0O���L�vJ�o���"�?���NVQ�חb%jw�}F������$#^iG��`v��Z҇+�s%����E�&@�F�F���8��-�$O�o=]դ{�2i0�b�<�AҰr\���{�8"<Kh��+u*�%zeY�amP��K�b4� h\�I	�p[X�23�ee_tܩ-�]$$�q�Xn`wz��zO��ܦ^aR�3�=洯��*c�UR�d����bk�%�-��%����Ч�7l��O~��}�J7
%�~k������9�<NGj��
���mWp��O�;5|��:��Y��H��N�r}c��Z�C#A#��5OF��yv����h����S�|��C3�/Q���+�7�D�>�"���cU�:�6H�d:�i�k=T� U�aݕb{��,�Ó�F�e��)�V��$����7)�h{��F�e����Oؕs����`ey2?��p����#��ۛ�&Ĥ�T��e�{���){�e"�}��:p!�)�=������ݙ�@@���j ş�f��H�zz}�h�J�	�ħ߳���+���.���lW���4ץi`6h �W.t�K�Pk#@�<�����&�9sI˦]�D��A��2�w��>���L��M�+������;ڙ�T�&"�g?��G����b��B5L��j������]ܜ(��͵[��wbo� �|s5�Afψ�tU��]� �L
KK�]�pnFBZ+ܯ�����!d<=����j�=���Ty����:x�]���h���n�T�Lt�0	����(#P���@�C8��+���za�MIW<�U��[t��PJ�p����E4�lsj�'�skTy[}+���W�[�~$7�KT���b��M��d����e��&ԃr�XX���lrŗq.e���I8 ���[Z� ��}�5��ߛ<�I�O�ЊZG�T:�_��Z�[0?����E�Y�8�w��� ���������2����D�.��C{�~��9�5y�pX��.O�PM�1���D��1SCN���z�vK�-L�04��?j�Nwn��\�g]^����qH#et�+��	J�6Vt����������O$�1�Q0���qg2��S85�X�כ:�X�Z׌+MC��#��ㄏ9r}��X����c[ʋ���6O��S�X�I��6�	�K&�/+7�~5gĒv5y���,�t����S,�V%׹`��'7�q���6Et���{W��(�%V���Ņ�ѭߣ���E���?�Vk�y=u�ĝzR`m�~ŀ����h�W��Ϻ]��|15��A��1����I7��6�n� D�EV�btns.��P���C��+���y;��~��y��*`ѧ4��9��|����d��vr�r�Z�ò7HZN!���(]���g�6���z��'� �r��!�޿ ��muגu;�����'9��d�:����@��36�������̙T�u�zuQ.��1}�G���0	{�n�T�}������M5n��8��ɏ���$ �"��j�Ԗl�*˫�+ �ǷX�Dy��d�b~�蓰m4�sb:��]��-0����{.�N�6E������v��H�M��\��s�����E�@������h�)�?o�ȱ���;�g���|��i�����Q�w�f�|�Q�~�=�R���j�r�H��c��{���3��b��,�/���s���5��f�Y�& ҆�垔
���6��D���g�Z����b��䠎7h
�g?zl�h���ype���F�؀2�{��?^~`��'��+�֭��y���C���6��J�_Z�ָ�j�7�Uilm����ј��F����6�y�K�o��~�e�X�f�y�����~��`�Y�j/_���ͣ:-JB��%풐�%3a��c�T^�S�y���xR~T�|�j��yu�����)�Cᒹ&������%����q ѵ��c��t��	��̍���ߢ����"XH�p[���&ғ�J���%�n��ՙ:L��kU� ���_����	ܢ#�>A�����O,���U��6\_���@E�dkw�(�$�����	�D7�)94>ç�#O���;u��Q��;����mٻW��/�p2��,ݗ�ͧ߯d�� ��ma ��^eiO<�<>8H�,�тJH]jG藡Vf+(
�:��&<�o%��3�����6����	�[�j�F+D¯��H��ԌS����CM��+����B�m�2�	�Z=�w��������)����h]l��B>��j(�q���NR����]_��'Z��ۙ��7$gk�~LLoNbS�6�i0�6<	9��`�̌��N��W�a0�Q*���M��L�}�R�6��r$�J���^fyL{22>6�7��dGb�/7!�n��'�U���0���B R�ݟ��<gd��%S���;V�H8�ρl'&�{zf��8�F�_]�*�MC�@��	Ţ\a�!7��G�jcg���3�@�!Y��\�r/D�Oӎ����xEĄ�(mJF���HLn�I��I+D�.o(yn���J/`o����~��h��v����=N=B;��͐9�ua�ٱ�{���"�����6i�c��}�i(F��I�e�l�+ˮ�pm�4=h+�-{uR��G|�̗etaUm�g�/���VqA)��I�\X���5�B�0	QR��Em�؉E�K%���m���<S���^�s0kV�Z��ח+y��lE')�zG��z��Q���`�s�`HHq�S�� }�f�R>]G��ע*�M�+Fd"�J	;}^�Up��"v�&�W�%���;!u�͛�F���T�ܗM�:Ha�R�5у�R��'�6��!�H�H1��@0��oT��\R����(ŵ�:xc�5bS��&/�(����m�e˒�+F�%����t�ajw���쾹q�'�{!n�術��TM�]C!�t�Χ�vҮk�~�~��K�*��Q;L��y��.v�h�Q��Wys�5[OKȏn��j�'9(�]I9�L�m:�r"Y%�$���i�xD"u?R�!��Oͼ]�Ұ?�x�Vx<�):�D��M/�n�|."���T-���;	$g��4���oՉ$/b4���-�eX�S�-�۾����/W��iP�gX���6/cd磿�A�,Ѻyܲ�u��9+D�sܳ��E�D�䀯2&˷��
��.MKO���g�M��#���RZ:���S�d��p�q��Y�7��Jd�w���f�X�2����Z�W�\��yt�[uu�~��vڷ�@���#=G�8���q{�o�j��4ަ���m�Nn�7����,���:_�3�'�9�?ͼ<�N�p�F���=N��7~�|���-3
�c�~��K��������?Ķ�"�J_��0�	Ik�.�W�C�ӭg⠔Ӳ�g#4��4uR �K�8]Y�aS&Q�K����(�y���p'[�?�F!����Ȋ�Eٽ-NY�M'z�����C�/��X�s `+���P%���*�Q�[�Im�jZ�g��^��r�݁8/V,2���u�֭\�v��V^�����n��