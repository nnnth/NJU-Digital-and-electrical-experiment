��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o`���d��]�v�1d	���u�C�[?�ϗ 3��kNm��5�/,��JH�Rw��$e NMF�K��w�h�0H�ai����I��@	Kx�"�l)s�ŉkKz׷�
��[c��������l��u�_��Ss��"�7�����K�Y��F��-Wi�ؚ`4���P�P����ԻW�2�V�gO�z�*qn3��|ע�Z�e�g�������!��4ωG�7{},T�J���5��Ƒ�~���80�F�sH���U+i����:U��7X�R�lR�O�T�p��d�v�������@�y���>r���N�U��h�N�e&ٚ�j�����e����-y�{{���m|^��}N)���-�u	��F�_Nu��F��ʊ���Ns>z��=��)m�"v���a�@ZP�I��UP:r��i�_+�L���z:�.��rx��\��*�c���!5�{s�_8���{~,TL 3��Y
$���w��������1c���E�GF\q�,7������2�Б�Ø����9Y��+-EL�����徯賛��5�s-_@��J*F�QZa���Iٯ5�g��-+ŧ�p��@�R��G���!�#Ƥ9�����Ц>:aC�3�mj��������O�z3����u�R�;tl���/���\d�e���%F^�̿���l������$*�E����T��̻T�<4L�Uȁ(k�gW�<{pU�����sZ����2F�.@RX�+��۱�($�kO4r[�4���.�2���Ɔ�8���ɳS��QRwA1ˈ�G!�N+ȱ�u�f:t�k��E��V bԻ�>��~�]�>�ٹ�&��¯aX$��q4��\2�����ӓC_]��Tk�-w�m���t�e[a�N����.���"�� \���	� �������F߁�M�)�������2��J�~qԨ���}��������d?�u�k1<�{	#-U�t疅�{�Ԍ��w_X0p.Su���@���m������=O�t��9A|�\���vC�1<�$�?:�����y�����.�#����Q�9ڥ:�@�G�,�?ΕэN�P�<���<�V&v��;C'I��bߕ�8���d����HZ�]��:i#d��>�l8���%����^(��j���ūp)�����r��ܷ��q�(���: ez�ޝ���?X�̬M� �~I.|^�ؐ�L��]ew�P��T��i��P�N��vv�u�ӿ�����mN�$N8���a^���S^���%M�S06��!���&����$-.�Ht�ߩ����<��@��Fӯb����;����c�|_��`02�y8'�䀫�F�!'W��o��o�1{+���1��I���@���mW�ٺl�:��h��씔�v�=(V�@A�I��K��{�;H��!%4`����d�]i���U&�)o�P��5��hW�,=*fgjP���O���0
��Nɤj�jI5���/'��)m��z?Ýδ�R`��ַ�jr��	 `�����n��:����1�zX����e���d��.�lT�����8!� \+�h6���S�"��z�>D����ǽw���al��&�c�$ù��V<jA��ژ��8o�D�k�+����5����kӅ:�$�A���Ew7FG	� �Ӆ�P����]>�N50O�P�F�~�?��"�_��:�6�f�7��o7º9gk����1���;z#*�+5o�Qsp��U�d�A)�}�-�5�82_5��q2E��έ�h]#�:9k�|H��w��2�t�b�aV��zʍ��[�V�bA��5�4�޼�� ��[�\����i�6��V���Fӌ�Oy"�����]�Æ��4���� Yg�B	5S��`�%���@�>L�d���d
���� �Q*~�h�4+�$v̀DI�M�h��؋��v���5�9�m�y��W��ϧ�����N���M�����'���4e��\���qGA���,��X�y�,G���9K0
{ߍ��
"Ly��3��^�� <��f�IZ�E=f�=\V���Ms�dx�X�k{�2��!�H(}H���ЁA��쵓b����T4��KT�3������Iu�F�Y��E�9߳_cp�W��g���.1+4)��]Ż3�i0�sł��+hx�dn��f�0�F�yw1U�?1�d�1 �Jl1E�j$���?���˚BC��G�]56j��=�ၣ��)�\�ۭ���:f)��7kP���<��-�*״����@E����.�D�bN����ׇ�r�3���n�8�ewS�Y'�B��~~����$z)�/�,!���͞>�`��`��Z�d���מ�|�M^�3^�r����Zi�e(��%�v�*j��|�[�gg�%p�ɀ��:�C/0��]�"Eb�ͱ�b��\�'LW�v�"��ת�f���T�H���j��lE���v��;%_R	\�v������^>�g^�l�ܵ�=z�ǝl_߅a��0ǘrKBO$���Jiy@���1[�߄j�ws�yf�A�*���IBjq�D4�)x���9�kȼDDF����Z���"A���U��-����[1(�l�d���I�=���w5%9��
n�w1 �J�t�B�*R�� ��$[�v�豕�U�I��+�L�G�C���q��?ڃJ;��=Xt`B&�j�p�:[aT������5o��E?�߲�V�uK�^2A�Nx.�z)�Z�%`q�k�8VH;t��^x�y�w���Z�o�7���X{�:��Y�i�q9�U#I:u����\!��'�;� �k@��� u+:�xi�:S9�;Ҽ��7�<����4����R���Z/#���%[R}c�G�Y�L���u*�(��<8~'�� �}���w�g)���H�=־{s^DK&|��b �ʝ��^w�3W�팃-=����"��P��L�O(�擕�R�#5��P%�/�7Y�� �JM.�x�Oߞ���-�Ԧ���QX��7�`*���	Z0��������4��V�\h�QG�.�݄[/��6ED��%�����������} �$��X��R�C�ra��������ȳ �0�����Ù%��Le�I�@�r_u��t��]�n*���8�4o'%��I���P'�<*�F���M�>8�M��(}z,{y̪���w)���<����Y�KI��Z opp0���j�a2�x�E#�'@:�?�^�q��Tʉ&��t��x���5"���eP$��z�'y��հÎ~�mB��Q�h�s�&^2�����������J��#t.+��<�BT �:�ԍUBG��Y��cvwPOS�H��Ki��M�T<����X�e��<�q��]ߒ��S}�����pR�R������G�`�Y떬)E�e�84.��uxZ���ڪ��X[)���>�E��A���ؤ������\��"bCq��������T ca��@�2셲CE�}��"�x���HPj/B�DdG��+�/������|� 0W|t3�����6�Ju����z�:�$�0V�%��"�zv�$��ԅ�|�zdg���%a�s��(�ohj�Y�gX���%�Ѹ�3[�M-�a��r� WI;��y����9���;V=�=]z��7��k�6�q�4&X�m�:MT#b=��Sd܆�&�!`�w�/�B�W`2�_���[�ŜlF�m�qS)GZ��a	H��7��+�Z�ۨ=�YAs��CL)W>|Sl��s���Y[�,)dJH��q��bz�iTE��P�C����J�s���~�ᢏ��c��H�aF�ob}��v�
�g�V���Vh: ��*�N�	6��8��p����T�/����B�a.��-����M���#mG�`�"���޲m���g���{ޮ�݀p�%AIR9%����#�)�w�#0��E]��'�M�֨���Z��1P�%�xg��TH�:��ă���k�J; ��L�e���0�5�B ����B芕
�A�f��8����<��n���d�<�uw0�C��n�/���.������x˖������
C�T�[y��K.�>L=K���J�C���f&w��n�oe�oؽ��Nuu^��p/7c��,Q��v�k������;��<>�y�'¼�X'��8�%�pu�oT�G`�N���WD�Ҥ��X�e[���oUO�׈f]�y�������M�G��m�Ms�,��-�ۚÇ;y�;��*��z��vKH�0��<�.n&�����:��-5!�7-;#��@���kD�)����I�g�����0g����p������WʔA;4/��< �����Ħ�<��CnrkB?c�����p�ǃ�5O��)���O5�4�0�b�:�����ȁ����D��~����g�や�*��
E�^�u�fa\�e�y�r\J*��]|�� �l��Hd�GP�r�x9r:>A%Ӟ�Mӳ��\*L��I%��Yȋs��y��`��z�]�\�?����ϛ-���4M`N������T@����׭��n<>"F`�n�23?�)�@�:u��]U�N~�k$�=ܹe����e����	}���6�
��yw�TQ�	Y2�<���F�jפ5�˔;@���#_��.��L�;!
XU	F�\���φ��J��P������@*L�h/g;j��؄n6*��x�w�������XhP�;(HC	?��<1C��+��?�\�
M�~���GK�y� �4l6D��%�^�D�暬*�T�G)�vr�>2��Yc���"f�~h�C�m�������15�-!8�����MA���A4��/�Va=����%i�d�d%&̊��_�d[�c79F.�ek���&Ή��z#"t,!��:�zoF��/ϩ��'�����$��䘀#:Ȋ�9&���$Ax��l����`�8�fL�uΛ��Θ�1��i���áS�n���I����O�t��]zz�2�eN \3H�6ɀt��m28��f��j�{o���2��a����A�,=2wv����B(�D�BV4&��Z��*�$ʖ��yj�.����<�\�O%��b/QF/Ûʂ4_1L����&b&�t�73?�/��ଟ��`���J0���k�!��7�DtO9��|	�R�#�҄;���4���@N%�-���"��T1\IuO���vA]pHՉ�4a8b�� xSq��b����ht�����v���[�G5�hC�q27S���2���G*�%go4� �����CM ��D�x,\�:��'�V���]�CٴN-
�B!�k&<�_q�u�����ݧz�v�����nᾒ���wW�n�b��C�-DE�%:��`Ѫ��>��J��g�OVǃs����39�f^�q�E�5��V]2���n�>&+zm`��ȟ�{|H��`�[�����8hM¡V����J��>�ÒȨ�Of��������B���	��(_KL3�����Ǫ�!�}槳T
.�- r��U��G�Qr�G������Yī���X菼K'H�ӷ���#�x�w���V7����q�/��\m�Z��U�޴)�Z��C1A8n� �:�U�4�[�)+F=�È��[���rq�*�:��D%�@��5�a��/��,u�u���OP���5�@�uy�d��'u�"��Z3�g�̻�EhFX
�5t���J޼^�|ɱ;�qTv3�Ʈ{U���|[��\��ε�Jfܛ��4Cr�_P��?ꚻ�A���^ݥ���bPz����E�C�Ge~*"���6�nb���O�D��l�&���M��t-�z*�J�0;b�@Q˄�^��aS@��(8T~H&���{M���)I=�<��zw^$k�G�Y᧌�Ȏ��A���\�;"`
*�8r�*k�c@ϙ�٨�Lr��� 9������n�X>O1w��i@��� 4�9G�@:��11c�5Oϻj���0�8X�8	�젝jٷ^��E��+�x�{L�F����rK�S�u%��X�v>n��D�	#l�J�[�"��
�R�%��J�J�q����e��YF�"5J���U����U����
����8H�F�֖5O��aQ��n���E#Y�3�F�E׻�>�������{B�Bb�i�3GI>�����}H��";~֛��V����+I- k��Z)��WC���V��V���B��"}{��j���86�~���QeO�+l0t�Y�$]I�2��/����{���W�br������ �N�&�Z���j�є�䟆$$p�]�`n΅��=@�W#���n�;Ӵ���w�IFQ��P��P8��]9��c�Ѩծů��I��t(��b�������I�3�ݳ�"P�&I��^W~4����5�:�Rlk�U�< c��ǹ�o;�#�����730�m�3O� _��ۢ�x�d�W�,�Ro'i��U;�h���c�O{�R3���ᣔ���CX��D͉P����Xlry�A7����	���d즚�Bxآ��݋� �b]]�b�� ����+���и�߬�kZs1|r�X��"J���������%1�F�Zc�����A��v��p�WE���[ 4�V��#w����xƭcS�ggpMκ95x��fܨ:��,����SO`�{��[��)�o��h%j����ሖb*f�3������F4�R�+�Q^�{�xW�5�*H�k��w)T����r.�Ѐ���{[����&P�=��~�:.�����嬭��N9v������<᳾QI*�o�ܟ9��%���%U�ax:���N�W�x���gS�F���0i��F�Go��t�# G��k��̬���6x������?M)d�x��,�o,�5k0����ݺ��nZ�f*}�O�L!����K[HYV�c����,ʹ")�Ze۽�?��66K~�%W��(+�Ƀ�	�����R��6̂���ZU[�po�R���R���Ȕ���Т��#���36RF�����#��@�Ͱ���M	7=��5���x�#q<��V�U����`��zsl�n��)��zw��p��͓��`�Y�M��![����7rʷ(�N\aWl̥X'�x�?:p*U~�@e�4�ʒ�cw�q}�Q+� d(-�5����_����]L?�|����"�����SĮ�$�2��C�XM��]�G��/�s��2`���b	Lb�-bI����"<���n�n�`��9f�qǕ�	Gq(�]\[A������9���>�xD'��'o '��5�(�bCv�}���q��y1�Sgb�b�O���NP�����فM!���4��'|GA,(t�1�B朥���X<���TԭvY6�b?����ݐ�O�;�Ҿ2�;�UC�=/���ϑ�!^�K�8�%'��k��!�B@j�޹o�����u]/V���OWV[���:���2���sxv��t��R=RZlj�X�Bn���e���ۅ�ӡB9��gj �Gx�g�N�nxZW씧l���h'�p2���M�{��{Nн3aC����*ƶ��<���Q���+�E)l�d;~-0_b�d�;2j&Ǹ�rȰP�-~�� ��
 <םn���j*������T��_S2	{z�)!+̉�i[WQ��5p`������&�1�+�
׋��B	�,���.G5�j^�u�6G�J��⋪��i1�n�Y�4���5����3R�b����u�`$��~ ;)J�W<�礼庾��h��6F�X�IV�"�H�~�,q�5��l�������.������<@�Y-����R|{"?en��:��T��I;	$hb\}����R�n�\��Lϻ��r�i��'��7�R�`�P����Ԑ���
?S��4�ju|H���x����{Y��rU����ę�ߚ�����g���i�R��_�M휘�X�/M���ρ� ���+G*����C�힆h)��:�5��q֛���%�CE�� ¬�y���AV���3�sݲ�eQ;���r �y�љ��V����q���{�1�7���q<2��z�Fz�$�(y���<q�.�}'�����i���8F�3�S���.�׆|e��A��&mD��݃�$���RӋ�m�t�o�W�fў��|�A"̻M�e�/��h����y}��#<��8H�?{��_8�YP/�O^�!n��yZ�ՠI����m%-7A�C}j�,�Eu�4��e�p�_[�ז�����#'c�[�D#��	H痝}�X t���<��ukT9{��Q����.і��Q�������)ʩ!fT��m�Y>�2��ϡ�[�*���7��H�`l���9䫏����6u� �Tf_W�#�Kl�5��(VW� ��z�J:_��)z8�;۟ຬA�dt���J�����)��):4H�I'�:�[Q���tƃm�VY�7vW��}�Ǡu�N�eR�e��䂰�xTc�8��6�|c[��{}Q�*>ɉgʻ.��y�cG����gMq��9>�ـ�^��9�h�}Hn� mX�;^��_�k�JJ�>��� n�0�J�bK)^!�f�	(��ܝ���i�`���B�N�I�59-�xPF���n+�y4���7ɂ8����D�3y�ʰ��5��w>k>Q�IC{U�G��H�t�0�����u}!V�@�,�Q�Se�"u��V�������KfK����[�q`=h�6iß�Ʉ6}�4�{�0i�Y��m��tA��A�H��6��:��E"S��|M*�J �����E9*� �C��nbb���g���'׎\��B��t4���@$�0�g�Ø$^r�,��1�|��%�f�{k���l�.��"%��˥Wl�,���.<)c��]����_��2�ic"���6�.2�.:�z�{x�.Wy�Q�ˌ��;��&�[h���`_��C�^�2�0�&'�<%���D��q�o��VT�H�[�}D�y��	Z4�Ӽ"�쉑��xD��WQ�U'ɡ�k���cؕJ�@�R�F�S�:Ҋ��W3�Z��@�5��8.��ab�e~�OǂQ@]��#�L��
 ��z�]c.�j'�
�T�	\ͷ�J���:��w��qLa5-n|f��nx�M��נ�����|*�T�(z~��ϛ�>��h���q�?�\l��N"���B���ߤi�PU�k&��?6��Ҏ�\�%s�9��-"ߞ����K�
x�Qkr���b���*cyK#׽<]\�u�)$���,k����`�Y�g����,���ـ�˃�{OL� W�O��nn��|P�0ԛ���v���ި������[������^@����A�;!	�� n�a#1J�c�їS�@������aeYLY�vEB$*�"�,�������k��9�C`޵}!�~��)^8UM6^�k��|����El��&J&ʽ{J�����Ҹ�n-}�-|2K���2A���q����Nz01˛�����jMw��pǋ��n��Ja��G]+�>w5U�4������\^��YeZ����%��t@+>^���'��g]&�S�mJ/�!T4~E�׃K�Z��Jr���&8PVb��&��JD�^���`�=��a}O�ܠgo��˱-�5�<܀�6> a�bx�|��A\p:�<�7XH�d�)�
-�"q��:�I�1,�J�&x�?�C\98~���{��o���(G��W���Z�Hj*��V�"�h�Hv��H���rL�'`UwΏ��J|���h"���@*f�����ؠ��" �DUJ`��I[Fe,��}���ƚ~:P؄�~�q�6~������d����+"����]"��'\Ԙ�
k�\)�S�ܙ;Гk	t�z'J�{j��f��JA�� I�8do�Α��8��=�+0SiY�=��K��=mB�\��?I�O���߃){^8�)���������I=�ѭ��}f�W��}e�R��P��ؚ{�	�ֻu�UU󌳆3��`�<�d�\��n���6��
Q�_���>ٙM���Mc����6�&��ς�fz�n��GF[�t#k�]�����
���H#�L�'I�*I+�`���?P;$>�ڌ(Y�vH;�w���N ͥ��%�gW ��i�/}���u8\$����c���^f�ȏ/>;&�?�J����<x�_��q4æq�؊&j�3,�_��,���*�3��EIE��8n������ܫ�,l�'1��I�D���z���wçܰZӘ�+	��z�Wi���|����8
A	��ի��@�x� a���鉼~��=h@�x�vee�v�<��P�����?M�{4��;r'��g=k4b�41���P^��~.?nB��98ʡ�p��YN���c^7�̬
4�%o�c}�!ZN�3`�Dȹ,Q��C�6]N�b��H�@�BU�����������Û�<�Qu��{YI�1��t:��EE�}HzO���A5<'�����a���x16�]���-����D�SWxҶO��ϵ��#�D���>��.�ʠR�O4�K��Y�̟|kNH��FE���Fm����G��䞛0(��E���U��9D����TJ#'��w�Q,��2�0J�mlW���nӔ~��IN�a�����O�M�zL�AO$\�v�s*�De0�H�Q̬3��8(�&H�shjj��k���`S��8p��>�������RǸ���I�B|�L�P�:ފ���z�-�v�܏���d��r8�<�"�ą����r!$N�����%S�@W~٦���|���؍n�ߘ�*�!�opB�S݋��w�uK'�{�5��j�����L���a3�G�E]��20�dC1�K��D
���b��$�95�:`��%����<ɂr{X���qP��e�/u�wd���kE�4��}QX|��w@�S.���l�U�r�����UxzZ~