��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t�W��M=��!�T ��V���o��Tz�Ӫ��ݲ>4@C�@k��Hs+���k��=s����$�SN�,�0�<s1}����K(I�0I���3%��`� �5Ai�յ0�:,_�E�`K�U�R���7kI�d�)��(��][�S�����ЅjT�x���Q�#ԙ(9��%�!��
�q�%}}��yT���l�<��D��U���p~�
�1
�4���o�|bNӄ�X3��f4�
��4t���Q��\[�_d�	I�7��v���_�¿�L*Xi�-���	b�b�)��6r����l�X�V��}�UcCb���ۺ8���S���/)8

'��	Z����ԷԬ9�ʽO��P�kN�e�v�S�1ߢ��o��eH���f.�.��'h�,x�ןg�ې*���@ړ�5�[{��7o}�'�H��I�uZ!q�Ԯ��v�I�
	����Z�C��a��6^��pz���V���H)�$�E>a?2��ƫĽͭ�վ�8�M* ��S�3����z�N��K����'��W�����v24e�rrÄ���тT!Pw�ӎ]���bi/�4v�;n�psX�a���]���L����SK� Q��̜�ش�$d�����b�NG~8ڔ�4B<�x���J���@��9�*��`�v��n�m�1P���Mڤ{�v��b�O�F~�sX�G �>>�W�yɺwt�g���������H�$�{����a���B*qN�10l�烝��w�}��;�f�)�߿s��]�0َo�g��8�N�L��`6iyk��p(a�i���
,��z��F_U�^@����N8�T޽}+��+v\\m��D�ݞN���!EE��F���,g>����.�do^!���å�c7�V ��O3�2j��W��o�V�U.��I�'����M�4"������]��2f�]xsO*���FDDn��VP�(�(�)�M�a��>+�Z?ӣz<Ӑ�9�=��pרI����o^	�a4$���iѧU�6���/Rwh)c���<5��ޑ��?�{�'G�)����Ȕ�E���<�ױ�jF��� �Yg��C���݌)��g4���x?�P؉W=��p3���
�@�SU���ٷO�����z׫��Vɮ�U��礥.��Q��V�a��ˆ���c҉��P�
�5HHj��������l,��!/#@K{,�\��bZ]<���$G���w9���)K��$��w*�,������>��EQ�����Gv����K
����;}���>k��9j����#�|y��$a���-�``.��mc�.c�Vp��xUg0kM��t�+f��?B�r^�8�
$v���0��뽕��J���S֤E�����r���M����a�\QFFz�þc�:�j0I\�� ��붙��Z�9Y��DK�����U����qer����#,Ej@�������;��z\�N��#�w�_wJ�?.zm5B��9���&{�rsO���Z��'����s�b1P'>��|�a�\r|�qƪw\�{����^�#	x�u>�w��ּԗ�:�6�������Fj	����,L͇D!���� n�[N���OĐ�Y^y�U%"W�!j.SP�*�7xTM����$�v����W�b �������k�����D*|�>��XI�F��,�C��+|G���˳g� [A?�џ������ �$�H=?�������H
٢�`	�A�m�=H[�CO�I^�Ł��D�u^���sy6�l����`��, ��-䢃m�T*��_�%��\�(���@F8��F �9B��?�)���M�{��wDhQ?���*GW�]
���p��A����}2��_�bݐ"�(�����E�)(8բ��Ť[{�7L˗�X��zM�����1T%@��d�� �|L�'�MN��4R㧳����2��~�d*�ANL�����ʔ���ۺw����?�ăҲ�w����5�cs��Y�o�������:$Q�È+�� hof=咲D!��S���I��9�F͏T�R�!G����&r�TX�l��T���Y��*r�)��d��^)�
v�~��bN8,�����<e)�=��5z��alS�ҙdQ�g�8��>�(�݇m�qA��g2�lc4}`9PUr�'������%��;%/A��Z� U�?�!��\q@�4�d�`W�{ַ�5=�r2+f����[W�E�� ш�U���ۥ�_j�"\F\H�KLMN٦ lؘڡ�̾�	ZG��zR�w��1����:M��cWP��m�	�I<	Z���*����u�WZE{�]\��(��EcSs��Y0�Y�
�"�%g�w���	��b�Ց:�G��3��g}ǌ\���u:	��W4'Nͥ�Dv�y�OH47����׉������{����|�-�V���"��ǂҭ�}]��B>��0Q��q��3� Q�U'�]O����k���*@��^?fJ��O
�1���J��]�Ϧ�����{{޳[��]���? q���Q��(���T��a�Cq}�-�i-p"�$���Vn��8�f^f�u���޷ͣ<\��clT��h�՝���P~���V�%>Xg�!d����Y��o�nv��S\�e	!��~_2����{n�Jy��`��"m5���z����!��U�R^�`�� u`��t�2�/V^�f��,k�����R�|w2���� =�,�ǇǋCێn�2kC�����vR�Y���t�X���>��Ix7����?��-��x��;"���/��6,w�%tw��h��m�Ֆ��5�)�u���;��×k���Q��3���U��B�f����$/V�Я�)+�J+F��&��:�DY@T@�\�3q�:{Ny�����9{0Nv�oD�{wk2�H���x�~���e}���˒�ʝ6�r� ��,��aƷ�Hs�M�NP���"�C�m�y,�s����cw�a�c���\;�c��(�XڳKË�B0�;ov�ـ����sH-�k3[jb�ID����A[�2��=]B�t�ߴk�ٮ]�� �|���'r�˫�=�YQ��h��d�9
q+�b�����^'�%��7���(/}�	V谸��	p�-)�Zg�#�5�t�Ǘ}��i�������[AC���-l�L��h�Ue\N#;.%��"34��U���-ַT�D%G��O��L;	�]�,G@�}�P��e0�Z��6l���	]"��������
���ɪ;��Oa;r��ܵ�5�F�\mT._���Ye���{�jGM�e~��a�8-����[-�$OE�������=С��k%��2�@E�W��I��-HBWUzH�|a�~�:5%��㏎w�8>-�qS��0�C9FP\���;�>�
����q����m����k�$¹�y�+9�������"ԟ䚑fk�d鮥��X�@�B[�X�~?��>�R�%����H��U��1�\���r�	��	��䕱�!D�P>�~[3w5���WPT�-V{�-#�̪�)�����H��9
i�R~�ߦ�P�E$o�[��ڱD�'[��Qxc�d�*+բӥ
�A)b(�E7P����?�n=^8(lBZ5()��:C��QJh�oe�
���d���0m�&10�ke*$��"Xb���}���>�FL�@f#T��Z���Gv5�a��˥���$"E>2V�<�(0
���ߍ�3���g{��"��b�a����қ'%m��fzBz�k몃��m)&�>�\�6>�$헡�Z���h�^���gN	�d�N)��r��|�A��<~;�y��W��������Xcn��0m��;Zz�C�m;��s���C����J�7=��%��A>}���J���'��0�6+�������~��)9).���*"|W�?ઙ\���\=ݻZ�xz���g:UdƳD�Db�D����P�{���ȞJ[� g�~�i!����T�����a��="թ����>2�&��/�{�y�6��U{3�|�3	���m5�c��%��7�������F�d;B�\��U�$}lq��jl�Vr9����L8�ޗop�_k���Q�|W�J���q��C��o�N�L���M��҃>�څ��V�V�F��f��HNaF�Kkn��X���&�)���\d�	�z��auL~��<yk�;�)�%�H�)0��Ѳ6uKA�������7��w�4#�Ӵ|�V���
��&���lՄ��Bʏ�|�yN��W�˭`�V1��TX�>��� �9Ӥ��B	L䝐���޶�3U7����0i@F4&N�Ҏ��[�EroM��$�6��ȅ;��ʺh����0n�w��(oz���(I��`2�1ÕTv
j=b�)��pݢ��(6s����⼴�-�J�5�	�B��N�EdZ ���ǚ|<�dK�9O��M��Ɗ���n��"���2��  ڑ����0Y&��-ܽ��!&��o�V�Fh~Q�LJ'��ht�����{�	��7`B�у_���¡֛y�ۿ�AC�L#L3[������n=�S� ]��C����k/%K_����0�!Q�U �@-3�H�>���e�^��*U�R^�\��IO*�
4�Y6P����9��"�{0�M�i�O�+3�7�K��R�Mu:Wx�ٳ���I��M��Ϻ�4
������s��<qԤ��PsSx\��Y����ִL)�\� y�;�bϾ	B��ʱ�1�1�K|��Y��z�Y{���G�x��,p%�t������Yܫ<~�=Y�)��j|8����086m���v�H{Κ|M�a;,��͌�qMJ&��-"�%�P1��{�,�����/�i�8˧��\�$��F����тG�x^Ej�j7S��RcI����T-�$�5�1-����p��Џ8����7��5���	2�'�}�ؓ���6
�Jr�O��9��\�ܰC:�@j��}�� ��m��c�+�%�
��b����~}����^.�c_�K�}�`�XO�%�I"&1kmԳ���~���s|~3�_�xdi�?i A����gtR��9
88���~Z>)#Dî���m�JCӋ.����,o~�,�Oڋ�%J�U�_�!�ڳ��X��-�x�?-��%�270��OK]�oO�g.�WS;�M��G΄7�P�e�t��]�i�%����X����{��l��A����U��h��1�'�|f��"|g^M�����C??��tr3q�R��ֵ{��~>���%ǲ=�qI�ڬ��I�����=D�pNb(�� b'��c�eM��qׁ+�m��ܼB�N�o�;�n.�ʶQ#ʜ�m�$��D�QR��UW�J�[��8��@fR;Ų(��~�+z�92�^�k�w��Z���#����R��A=⓷���)����8�'	F�_!iǫnf|k����%V>�z�$���\��R)U�a��K��N�+xٛn��!�������Z+�;��s������
׿�N�V�84B���eo����~�I�u>�L��5�>Zt�g$<â���'�hAd���1'���!qj$�f�k���m�p���|������SM�lH(��>>�S��0ͻךhm�������aB��k6+��+X�2�lNO���1�b5����m����/�9_؈����6Q���ǚ=|1UˡN�'�C��ڬ�V#%�� �$����W��h��=Qp�IG�c��ξ`� �LJB�WAX���)����)s�>�����|Vg��A�K����Ϋ?��+��W��9�����0��NS�T�gl��[|���=L0ZR@�Y � %&��ф^���n�Tr��7�%�7u�����zՍ����9Í�s�)!���N,���� ���FvP[�T�/�`n�������l�\l��5��OA�1O��65����D�_�O��ߝ����HR�m)4�*#m�g�Y�Z. �NrX̪5{��'���qw�qEu�^.Ы������c�껿-X��� *g�q.�X��ܘqZ6A���_�	��L�����K�Ul���gk�B�:wJ2�䟨Қv�	�r���9��Fl�_�֘`*�&ά�r�T���d�8!#h�+C	a��`��2�q�;G��ɥ�E��e$��Cr�@%%~�L�7'.BYW��i�X��l�f�5�I-`��*�(}�Ĕ�a��a�ށP�`���g����i��ۙ(�"�ϵh)������'OmE��KB]2a�����mu�̌^�<��`M�J�sS�(b��@�3 �kZ��%�w�-�q�9ݽ����D!B�}���H��jϣ���Om�y.�T�.>�G#�=�ԅ�����
M/�p�QB2߈���]��_�T� Bb�9�v��p��py[<V�!?���?��6����r���"�r��sI�1�Z?�&��i�fh6�N��������}�$/�k��IuL����ۡ�K���G$!gh��^��O����C�vD{��PROÛ��oq�lw��y;��16�Ү.�78��z�)gOa[ΰ�{�*V�^�I�A��<���y��{O�N[�;�s�ɝv��*%�~����-V�����W_Wt�ʼѯz���1��{+`�ݫ/���7�4egp<R���<5�8'�3-���r&*IͫJ������E�!�
z����#��R$ b@~�٪�L����e��Ë�w�E$�X� /�¬�;�/��'�Z]<h�42��P]��ۦj��� pF&�q�:e6��B���ɿ���,bx뵠����D��lh��´�l� �`�@����U��i�����j:s.�{�q�+� �Z��uɉ���2cK�1�U���{ד���}4�$��L��0��G��q'Y^6��,#�Y
X��T<g�^?LVx=�D}*+ȋ�(���3;1n<�q���J����S�FuL�V��8*�8C��HYCR�L�d�f� $:�~�s;a���\qc�F��У�ܲ>a��-0q=�^
�Y0�����M�o��>�������o���6@��\�!y#{��r�"�f��}2�h��g���SߌFi�i�z�m��A�`S�����3��hX����Lz��(����5�,����&�5=��8�0�'��4�Ҳ��K���S'G.C�b�z�:�E=�{TEC	��%�������<�Aߴ��9��x�Fq����}TQ\
���-[�c`���̝O�W,4´�� nẹ>�%��cr���l~��.2���3G�
@'�إ��6�$�.݋⟥�
0�5Yx#�s����_n\��z&���F.�~H�a�U5��=���sJ�\�b�r �m���C��*H3֬kk9l���۟� ��lSn����n}�`Z]�R���vD�D2��{΂�R�GPx��]c�\&�x8�M��zJ�����" 
!Pu�S�|S����˕	�'��6�|bNg"	]�{B�'A�2U�Û�e���LxE���T0o������"��n �hp��%�(�y����3E�0r0��-����ŠӞ0wP�Å����/�3�W�i	��j�a4�k'�/Ѕ@!?���}��������f��bi棢���Ѧ|a�	G�6�4}�?�������f~��r�2�����#O	��w���ԴC�W�x���V/����7u���#�~1�#EHX0f����m�+��������d���Ȩ� �J6PG��*�M'z��E� �>MB����hh���=�����_��^YWX����L�����tqƹD6����|1��+p�:s�K��������t5�����K���w���|� ��-�`J��'%1fM�I	XF��`��5@��X	�+��6z������_i�����\P�_N�ig�ΥH4��0�<��S�p�t�)�X�Q�����/��Ի" "���	B?goiή�"������*�9��zƤ�2/)
�<0c��m��<ĉ�opK��f�e]�<M' ӄ=O�:���R%���܇��K|D�mM�Sf�b9ƀ� �g4���c-}�
4?Y�����RA;����7�̗�̘�ZB��T��WݒgwPnd0������:���z�ҪVI���4!F�RS
3���Z��pt��n>9�5�J�g$�-����X������`���e��z�!�Ū���,�9��m]��$���;��������;��P{����}�%������M�]�|�5���O�����&4���v��@	��4H:�܀� *)�~+M�M)`~2��g9Ψ�p=�P6�9-�riQ{}%\dH�DP�Ar�4���XGѹ�*�JH��"���$""��0�fK�@՜5sғP�]���Xu��R�c2�b!^��r�T���q*�B�4�VS/tÎa?����T��xgʰ,���¶
��k�u��>�X������_Nd|\`]Y���!R�z2>մN�sb��ʇ�v���N�m��2��.7����i��bp*�Ĝ*�c(j=��KW�%zgA���Q*X�i�e4#�z�lrk�v/�.*�ds���j��w�y3*>
�\���˺`�zT��"ݬ���3��B˚gTq��Ԓ�:�6�=�p ����c\�!�p�4����H��v|f�5g0X�:l��!V�"�=��$/;"�������|�"~��uI=&�~��k�X!�p�N�k�+�	,a'ҡ4��y�`�Yy#%��+���=(&�6r�6gK�~lU��F�vR��v<q����o]i'|~:6�7�����g#�!��)C�Af7�kK5$��NE�<֚d0%_�{ؔ�[�
��h�Α��ኆH��,��-��������	R'����w��t��9-���8���<�M3�y�VڙW�m��U��~A�x�%-�E�W����-,!�� ���P��v;�Qo�fu<jר~�շ
�a���uR�����R*��VVl/,h��`=Fm���j�$�i��$�C8r�q���VsQU]X�P��a�A� ���p�kf���j��'Ɇ��*ci���b���t>��粜&w��������S �S�Ľ���ݩ��f>��j/��FY!�$`�]O7<�~5�{�YS�0�p൴���P̧��:l�F��R�;4q26Dz�=�\�l������3 �{���#�p}�1��4������EOJ�By�\�F��risz�����O��n!\E���Z�$!��2�P�҃bG�I��_�q%��Xo}_�Q5��gI�m5 ��~���4��%�-�����o������Y3�ݰ�j��Rj�v�C	�H�I���R����p!t��{T8�f\0I��e"
2�Ejh[�`F�:�����-���qO���MR��>�A�,1�Yײ j������	A�6��~M�
�V6S�a�4�Ч8�8�=@�s�}��ŭ�&��`<YG��4u4��D�S��`�-����w�� i!�_"a��6�(tש�J�����O~�n���u�e�L©�
,7�G����>tf�ɲ\m�s�sژ�x�8Y![*����â���#�
����^�gO8p�S��gzԴ������V�S�q�*�j��iFa�\�@M��O�0�k)=� ����Ю��R���(����gfT�� ��A�t�ǹt.���'�Z[�9��>U���g�a�ƵjsZ DD�����-jI�`��.S�ҫD��T}���Z���C0Kݞ۱BD��NV���iϽ��5�7�+
b��g�%�I�~m:WN5�js:�˥)-��ia��Q̭b�@���4k��h��2�r�\�Q�e��HJ��鉱�TjA<'P�7I�Q_�p�D��u��c��������8',�A��<}�	��ǣ�%�_��@��=���FͿp-4��ʔ�Q����d�L!o���L��)��vcJy��g�bS�L��Ƅ�;v�D3��[~"�\p�M��2O�xP�v�����Z� ��)��H�rns�ӻ��姘�	&㦈���r����k���e��~+� �g� �D�{!�����"�'��	�4FN8���P��̣��	��5�y��v�,�����Tq?�g:Vd�m����@љ�1�A6�l���$��5�lOvvJ��aCE*c�a4�@�j���f�p�>�R�c�a�{-�a�OA]9N�AU�T�i�'k�I�ut*i���A6q;�&I�P��5��(ȁ�8�%�{Z��<��q��l/��o��� ��������+K-4d��j%����":C�[�Q�s��W�@D`���,�麈�i�.L�|/Q'���j��%��� �D�[�����W̧qI_S>��W���fjr�	��ΜJcH����$y�`]<�<yƴ�|�D��K� �zqa=�h���&�U7�j����Bs�fU�zP ���c����3��l�K]�71������{|�a�����r[ w6[��
���1&���rb�\M�&��=C�pJ�od��ު�X&�����d�Hl�$��H�k�����B��jY�/��E�Mӕ�����g��s_� ?g �%Ncڶd�a� 9ǡ=�f��2��9c��|z��o�2!M/-&=ַ�3�9�$n̀x�e�$2�����9" 	�Ja���ǌ��y��DJ KL�ԞJ!X�'�<������d���v�)ڱ{'�tg�.=����[������q��⽮rl������9ciS��o��2��B{����&���� ^k#Ϊ��'=v�A9�5�[I�������Ǜ�Gv