��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]���:����~׳�jB%�Q�*�U�&y�z{`@�t�#�r������(��G��?2�F@l!�j���Sx��a-k���]4&�B��C��T�3H)*��E�%�J�
CC���r�DB�e`���?)[��
b��傈��� �+C4k�+0W{���1$w�P��i���o���y������;�u��;l��pvqՠ���j�LL�(â��e�?0��#jW�3i�U��<~g�o�K���4H����s.�Q��Y��#8"4U��O.���#�&���P�'0wb�3�)Wa»%V=?oհ�z'�&��.Bw�]ܠ�"�.�����< _���ن�l�y����i�8�lP�� ��B��H�3���a7����-�3�#��)sP�ny\3!���ˎf��M�����8���-y����U��U������7�1��עG�{�;��{<kT��՟疦�D8\�+I�~W{ ���P�XXd������"�����&�۴�'ϳs��'�$�0���e*�U��ŸT�Z�G>���NS-ս��0���N�QIam]ck���	���r�G1t�.��}cZ�b̀@��B"���ʠ[��A��d�JGuP� 8��_T/lh�kw�I錀�P1E�4(!{6�cR }�=5ʷ��󜊶�ZL��=}�5����T�M/��,A�B��J���*w��7��I<" ez1}�V.�I`�-�~ό���oS�<#%k�̑B�$Ѿ���O5_�.e,�Kz�Z@��D�����=&jF��#\K�����#��7��G�0T�(;eq��:-u�ۀS��R$�q�'(]LWU�Zq��].�WBc׿7�tf���亣+�3vg2�3)|a�{�����=�/t�UP�[V�-Zj�����bco�AM�	B����!,iN����;�-~,�1��d�c��l)�#:���Y�rF`�yD���eZ]%v���� �[�1�Z�KkB�F�G���e�6	J�3�lt�f������u7>�x�.m �le�)��fu���%���M::�X�N���ִ����$�9�7���d���.�.�L��&s鮏(�%=�Ϻ�L�٣�"�p�}9c���������ȡ��OC��Z��r&����=5K�0�q4ۆJ�g��+3\l� 9� T�R(�����/;��-�B�G[�{�SdD �d%�c�R/X�UX
�y�&��XGYn��j0����l�^$x��&�	n0By�JFXq\H�E��EB��9�K&F�b�М�A�^�/����@'�[6�2��{k'v��!p��K/m�n���z�!	F�K�b��sQZy:+ƧqXZ%]Jo'ar%��J�d��T��1��}ˍI-�H"�/�S|�Oؽ!��� ����u�k&��q���z'�v����EBgA���m�bJlE�]�Gs��&F+�ftS���M�oC�EбwE�3\t����f&XL[dL��_�Q���Ia��,j^?�G��VHݦpKž�	��^�nd\<�-o#�zwؗ6"�<j��}q���r���������.��Vv�z3�W�`U��b	����O�7�F�_��v��\057�A���H�R��5�Z������ľ�>���?�-{$~�5a��;FV���Yq���ݎ
����6�l��=|�u�n���8�e���r��,�!m,��=?�k�~�MLS���.Ѽ������.F{��򜹄�(2���є2�s��-�X��t�>u�~��� ��ҙl@�3	t��_��B�A;pr�u	�}�4!s���~{ִCn�����ա��M��#7�T���~P�q��l�������tb>'��[hf�|��\)�M��qq��V��dWDd[�Ih�X��sW �me��'p!�`�gY�Et���>S7�	v�#�\[�{����(�ǟН縲tݚ� Q�;c���}�ڸףlw����0��Q>�H��i�JX|�v^Cd�K�2X�s�y�-�\Βhb���ܓ�|�7�e�MX��|��8O� ��j�/�<b8�,V�՞a�c�g�7�\Ť<���H�����	������ݱ�7�n:�^�����~�y^�NL>��'1.�JP:%�3�G��[�P0r(�,��f�\<־��`�
�&���gQ�-�T>��6��Gs�����% I��/ŧ���R1��@ �
����(���R��*���6qe�=m�B�b�QUm��rtB�N)� 6�=T�G�ǎ���"�<� ���r�4�����gR�-��,Y��z�F��t��Ah�A�fo[�g㑆�&�P�D-�a8C�ex��B���
����6:���Te�x(��v�f�m����Q:}�+\\A�(QwKTW��$���$*P ��T���s�D���f�B 5؊fo������oaԠ�g�-B���C�N$Ȣr�"o�58I5��Z��=�aR�!�U���%�#�ѢC�6 ���k{�^����rř�?���얘{5�!"#H����?��QR[��d��Lq�\"��W�KGf.�D�_D�+_t��l4g�X%0C�޽:�V̍��|r30��=
k�Wt�$��P�'�v��Jo�����IK'K2��k �%:��V���jb����%|��hFo�h�1JW��k�+��ޤ���\zq5�E�G>/��Ab�����[C�,����e���-���GQ�S����ig����F�";ٯù ���o��,^�=�D�,Su��,_7������h"
�~�ob�t|3�[�'ǖ�S���Z�2�|���74G���P�S9?Q+�5}:�hn������\�=v�*Z�#��Ԣ)�{nP���j��y���W��|?2�h{o��e�0����9�LF�c�	7p\�4K�KB�7�9*���7n,ю�a24Fcòl�%�咟Mz��4��[�$B�9��sH��wyⵈT#<_+?�*&[�f܇(j��L��m����(�o�K�j>=ܔ������5��PZ��7�� ?Sx/K�$��"�6Ҡ^��{ �=��I#�3%��G:��_ʅi5�{'�kC➚.��F�x�Y�p�%�Gd�4-K����+�Ʌm
Az-����[ ��'�K��9�^��z���zo`ϕ�Q�O�����0OL��J��w��(���UE��P"*HHm�JwR?Ȅ���Eo_�s��2�V�@��4��)Xv�?��U�]��T!l�6"x#̟Z5���|��8�����g���	�BC��5�ZǓa�����o+B!�B2ˇ���V�#�d�ґ,-,L����R����y=�#9+ڧ����������ڎ�*	ȑ���HP����M��]2�6���4q?Ohފ�^�ф��
9O��hJ#�($t5�_�?��Ʌ�S?6�ֿO��p{7�2�4)���=W�)���޽��PǤ:w�$��[�^�)��T��	��DS�qq�q�����j[w��̠9$0av�g�:��e��z��H'�4��np	U��)IB���'�PÖ���;��X����������a��u��5�Z��;������w��=�h"������ڿcڠՐs��%{޼��Y�\aa� �:�2d$ե�?$��^sL�}����m�-kr2�(�2�2��k�Vf�ʴ�|��]^�r���2l�"v!�ni��cہs���,1�� V�!EA��G�����q�BG���J�6�'�K1�7]��FG,cH��wd!� ���tء��@  �KS�^�>P�+e�š�V-K�jyd��^�B&@A���!ҭ�T*#(�@��I�C��|���$pٲ�u����c7����'���f�뮴 w��w�=�Y���r��!PC���[�yآ2�����]���f���\�5@�݌�{5�Vw�\��E]P�<� �i�\�W� !5�H�|C�c^H�㺊ec�a��*r��. Y��P���Gr��8�Ja>��}��e �G�5�K&8sX�e΁��KL�I��߫��XӖ�������r��@�^ª4��%�������,���Ǐ�w��٥#�f H�P9]�����Z�i����x'��9BY��p%op��~1��MhLI���ByS�/~��w[�੔{S��U�<�8t�ݩq��ql0$
��0$��@kͰ�[�}���m�K�+�;%♧Ч7[�(�̈^ʌi<ְV|���p=3�Z�������ަE�lv�[���\Qw����bgC!#rWz�ءG�F����d�J�<�/r���2T��t 	���ڑ|NIRjS��S�����s�Ȱ�L��N� �*n'��I���� N+�{�ށv�W`��H?���=)�Dl._�9�!�ޅ�MI��`��y����O!7ܞ��%M����C]񧒏�]�Zץ�"|�@�.Hf�!�K[q.�!Q0#,�O�Q��7g�v1~M�rG�|�!�}3��]�uh;V.g��%�|�� �{/w����Ò��<{�%;����.2�����g�;�Ry�4��3X~-����P�@�R{}�XC�si�8B_$!���d�o��P�~ߎ�+q�ы07%I���K�
��Ϧ� >t��V� y�*6Ŋ�0:^-TmH N֜e�W�1�c}�,��\=3��y����!��{�
bs\z>`�4]�AL���1�bu�i��fj�P?��6�ֵ��;]tL!�t��i��t�8 kW46�Xm�l�n�*@Tp)��̕Tu�u9X����b�>J�k���g3���'֙���AJ��.L��xtc<̮մS�L��f`��j6}q�� �i���F�Z&/4�̋����KD֍�-�Ŗ*&A��X�GD(����G նSʿè����ġ|$���8���d��(���a8az�0�z:��dX'� 
��I���P��I�Ig~�ݏ �f���?2�Lk��6�A����1Zj�u�:�L�� ��H��y3�&#���������ӗ���ŗ��n�X^�������l�PV@B�zS�MNG��\�-�O6����������yo��������6�����[3t"
o������;�I�vĲ�4(��a�[����U����:1���8I]�tS3���1uƁ��ˬK��^�X,��|��IND(�>[&;���ۧ��TaةL��ŵjK跩�`�!M�Å�Kīa6DkgO�u����9'�����V��&C�gP_�GU��T��J�����[�.H���n��)�-�����D7�9�2�ʰ�wU5sr�S��4�=�+�ۓ���Ԧ�k�#���c�7�D��G73�l/c�b�)��I^	�kha-כ�a� ��!�$Iѯ��47�{��[��[�qD�]ho��*ne�qp��݈)��i�@�G܋K�K���g
5�"yW��<���dc0C:��c}HEF�1̨�	c�	�Q/�"��v������Y�Vy4j�J��^�d���3�"��od  ���2d�	y�#��m��d�5�p�������-�ƃ!�~���Bc�N�E�xo��p3S�şJ��c�V��]�N�%�"��]�[!��Y.B�)ɫ#k��ڔ#���p��3@� �`F���L�����I�cdt�&邴�@&*r��W�G��ꩉ֪a�����LE���;��6;�ݏ
�Bi���W�`�0�ru,0T���=��"��Q�X�am�k�֧:��ߥ0� y.��nLu=o_�r7Y��@&ٵ>�̣U�$4��jŘ�nMY�We�9��!N��o�������J��8���[�Y�P�izS�E�R���L��dGT�-�>,¾5�W5{�T����q8$8���a ߅.8�K렪�SNx��lx��H��K\rJ?��f��C�`v�
m�'���1a������뱈:�m�[JE�N��e<~��ɻ��!L�ãr���Es߈I�BX��M���� �ȇ���l���0�)o�@Hhm*���
�2<�����Hx��Ȥ�l����=NTGU�;{D�=�?�}��ܔ���р���F1<�4[�ղ(b�+L�?�I���ո//�����<~\����{B�BƘ���O�:�>g��о9=c{{f��N��������[a��Qˉ�>�k��S����s���0ņ�`�����XT�Rt%�.�gu�7��z��tQ�1)Q�BC���-��x��J)ɘte,���E���"��1��2O�t�l��!�S
/!�._��iJ)���,
���+Y�D�Ug��%ˡ����s�)�L�C:��-�c�oS>yLd��-;�_fB:B�������v���.�f�`��7�c�%P"�{n�Н��n����F`TM�D�mR�/�&�H�O��9(�����sᅃoa���į�s
�mZW��������r���pr)�K����F����ܘ{o����`���3 ̺�K�!�gͩ���X]o�䖪��8U)S���C��S4�Ed�7%�k� �	7�j;��(�DR�R��$zA�]�i�UJ��s�n 2�g~j�����)^�G�N�\{�������R\0<�4r=�b�PD*�>{Oy�-�};��q��Tk�3V�m�;6�r	{����{�,�(�L�A�jH��޾ڵ;k�Z��� {��|k	5�,��!k�5��o�5�X2����ޓ_Ls2������2i�(��}��tLԝ��@Mf+���L�T/���*�Q`{�F��4�Zq.��v�'���[����\���گj-��]!��$���b�R��p����ܲ>�iM���Lgz��S��J�`z��%����z\�H��:�N��I�>[�Uw�(��׈�
��UqG����E�)�S^yJ*�E9�9�@�� �#�K�n�?�g.�L�S@�\�l Z�k����P�Ƃ�x۬S����[f��H��4Op���&=�O�t������,�nP���������q��s�MHt/,A��'�iB�	�h���Gw�־��G+� ��;�������K��E��3�d4ӠF��&JK�jx�N96d�&;�z��7|��sJ�9dX�D3�q̍��@���/6d���2��Z�X�]��k�t�=�M��BF�?L��ɢ�Mv]t���f��#d�&��؅�r��iP;�#�nP����ka�R��s��I�A���7(�l+?߫g>(�ZJo�մYf���M�U��P'�1F��`X|��*�9�͚�$�r}6j��s�j +�$`�:/^W7:����)V��&3�]�H�$�WT�T�}��FΆ����y��������1Ɩ
~>�Y{!��LI������B�$�R�jj�6\D�"��8���S	�p���{U�=�ʯ"����2���(����dGL%� e�'HL31�����#�G^9��[��z�����P|���f�8�Ch�+��t�@0��*����<��]-�X� _�C�k���C50zǕ���S= H_��ya����-U�AY�g�*��qU��䨹��G�>��ẏʱ��:�sz�2U����w����0+��_�~�Vy�B���}s���H�g�l�Oۦ�#F٬W�Y�hïG,�!����j!�t�����ᓔ`)�{�*j�r� �����{ǐ��]I.���Wv�K|Ͳu��!�;�  ?j�5���x��0�MQ���L[Q�����3'1���v��[����dȭ8�R�9'��[�X��c �uUz��v��v�й��P�I?��3���@{R�=��1c���n�"ь�ݐ�ٍ���l�����#��]��h��Ψ�':��������&i��	�m��Є@��f�#���OU�a�i��1~
��Ay�y�f#��%�/����A��s���/<1�2���Qa0�?6���\d�>։�4�+R�gi�\E�Iu�+��p%��y��>���22�=:<���ck�I��ڕ�<y�z�W���_a�u?���j�8=tV��_��^ݿ�w� ����Y��� �K���|�Q�I��\!ek�T��ԩC�%湵�JF����q}|�!bf�m䳕��~���k��9q�S�ɭݹ��>X�0���~t�C�rνĴ7*˲T�[%��&D������f�سs����{�g�P�n&;������Ϭ�|����˻�	�q# 5�<e�^��̮��b�Ǳ֯#�����NgR�
���(�a�:�_�����fXQ��g ͚�J��B�߅U��Y

W'dov\��N(�&�W��o��V (����f�#��=�'|��<ɋ�F��wٝ�j�"�I=W�ذ�(|�Y�I_�?@[I����y��C����l/]`���OWBђ�ޙ^��2�a�l4�&G�z�)��FH����I�xc'��s�xL1@�ش�O ��Ҡ�1���R1��	 %,�o�LeמB( ��{f�ɭ[���������3AɵZKD�"�Z�3�#V^�B�*�~�q�4ɶ�[�Z:Ǭ|E��]V�ɥ�ڢo±��/�H����f�#W1���	|�)x�UPU��q^q֤�K��Z�|��Pj�>�~C
JzIQ Ns���D��jٵ�>s:_�<�
:+�	��Jy7zc{O�S5v�K�������B���ww��>;��kG^�c��هti�m2s�x�C+'d�r��H�2�|�w���%�V�E��h{������qC�v_��k�!�x�����A��z9��F�7��Z��nH�bvS��r$^����ފV(?eEV��j�F婦=��!.�h��"Z��-dG�>���CN�L� *o/�*S����	k_�|;��l�1�~E�{������˚:=�]<潞
�Qf��X���RZ�z�~��r�8�=�["��>���n-����U&��Y��WxQ%LSz��+F�2pÀPS(n u/�E�]F3����l+�-8���J��Y�����xG_�&;��P�a�>�Ы���14�poM��yl~9h����
llֺ�2�?���!qr���D����D�[�-�@�8�+R��3�x�{n�|��*�(%��
���v��pm(p`��L/��jgx����xxq(`��t�8��,��Ad���u��ZL��A�/���)@�d��p��3ӧi߂Z]>�H�E��� u�%s��E�X쓦�&i�������P�Vg�k��hx��J]�)r���jt7~�%2�ab��C��Hj�I�x�N�W��j�Ͱ�l��wPⱣ;V�n'|G�S_:�nZ�a�8��-�D�����է��a��ź7���N�z�Y!���o���rz����Yg�*�җ��Q�0�����R�����.�����\Gy-����D�2�J����X?Cn���~�$o�M?���UOS@�Tʡ��%I�LfM
4�ʛb��!�Q�B�>�m��nמ�!Ꮅ�P7�ʨ:��9G��eX�]6Zd�7�[.��D�v���>ig���ů����13	捝���^c�u{�"��`���ǰ�>�0� ��ؾ�6ܘ��&v#���=�H(7n0+l����>L74����JR��d�-��R���cH\Z�곲�K�Ɉ�y�j8�&���9�IR��M��CX�0x��`.:�b�7�*��E�������Q*�ՙ���[�Lh�x}�����S��V ��4z�K�����9�O1���[Z��ui�T��+"m%c#ZfW�:k��	d�^V����t!E�"5ŋk=ߠ#!�WrIK����O����(�-Y�
H����e��z!oG�P��{v�� �ƛ�zg�"���^�#$-ؗ�9���V��[��Y݆���A���.
��M�޹߄UE��������9am��
�cإ�����2�(���00JUWFR+04�I5PI�)j���$�'ib���"���q���z5�T\;�eo�����1��B�.[�w0�C����D��f��d����Q+n�3���ZHI��sv�A	���Z�5�vGV{�	+����X�Y��6]�F�-�[�f��*��ҡ��Y1֞�.W���[�So4O��ற���`J.�
I)I��o�,[��Y�<�^p��t���Z�g�.��}:�h�!T�H�b/��@c��1G�������X�ۡ�n,2�c_�i(�=/lpr�nf[�p��I��W���c"��X8n"��쏷vH�B����bכ�D�!m� �Sl;�]l;�){��.�E94nѳ/���$�Ii�����8(sX�f��*Ϙ��x	�J=�:�z�g
f��� 5�����b��}ߋ�bį6rG5�:�c6�b��B;�B�.K���uQ��#d�K^�����nW3��^��1J,��Z^���Yb�=ml˸�2�+CGm�8K�'9~�?���ݵ�Q���'�'�y�!�|N�;�0� �C�������i	�^y���M�T��?���ux�e�
������_���Nndx.��1���P�[肍z:&�����>d��t�w�T�*=mmOT��`5��z.���u�9欮ޫ��FQ����V> ]�kI��}_��}��w��������o��3ȑ��W��iM�? C]��}�����̞�>(ʪ�m�]=�FnrA�)	�g��w������P�0�@�X�@L�`�cvX�M��Z�]�gT��SD�oղi��t�
�_��:�^��^��`�ׂBc�s�-�޾���齭B�4���^:��s��{11s���Ľ���^p��V�i��kЬ �f9f�gg
:S9�ҩ�fo����qb?W*�o���7J���i�'�<�ӯM���%Ds�)OI��"]�_]@�dٹ��H7I�<������5.Oգm�O�'�_��7���=�Q�X< 8�C�wB���}Ld���G_�T�4g���5����kF^���T��zF��L��N��;f��)��C�3Nr{k��4��)/t��m����p�3w?T6 �g�Tn��߫Z�	)
�@yQ�� �H�#�e"u�뎰��������V�O!�!,/@p#z8����S�JV6@_$��G��5U��0���82�,2����1��a��OƳh"�W��ڛ�]�<�<���}V-9�BA+�:u>\�
���<M����y�nF�T�7	ʕ�n	��15��{����	�#Ouy�F���.�A-�:�K��)���OL����n������/�_'���e��^��n��3�4DT��0NL0�/���9]�_���k��r�*���u�{]s@�n.���s��h1��/�P
q"vV|*��)��EM��-�W?��t�=d�\��"�r^S�9u�(AE�|c)4:3^�.z���c�4�c�7�0���z�Up뛝[�0ڈ�&[u�T�_��sc�1��'h�-	��6����Hn5K�M�����*�$zM0j�ѽ�\| �~c��j��M�xH�������nʄEtj{W,��&��۾XI[M=�'����3��i�,� �]�^��,��8Uȡ"q��g���6�D�����I� T�Ʈp͎*Q���
�T��"�d��q������ �t�k�Ud����3�R��AtF�׼��©��|%�3n(����
KscNx�Cw�'[xe��b��P�/��!1)j�L�) �	�m�%u8|CN��6׶dBvǋ^%bf�H�!��l��c��'d�,e�S�9>��7��o� �h#7�CIL�������ĆW��m�
ȐA������T�#��ǝ�wb�X����Ǽb �Ju3�R��sXc#3����lP}���6i�y���-�݊�ߍ>
_�RH�o��9��:�$J\w� �fE�HĭK2���L+h�;8HrD�+{&x��;:<ɶY�쁑u=a�.��;��^{]�����,��<���:	�(Yx�⥻=1pN��%����C���{=l���粮	��6�Q�>�7X����3l��ޏ��6�����.4�Gw2]��f�(�]�x�f��a�]qa����#	p�c��@��!;x%5���)@6I��l�Qm)T��}�>�BN�VKꩯ�ױF��j�b�Q�j�����;�`6_L�5��Y�Ѱ�d�]�mx���.1A�|���^S�]vp�"�g29[Jl<,��iC��2��t%G2W$v0�]x�Z�����-=_��߬�<��$yf�'<�A,�!d)2��k�Z1�w��A-V���ۻI_M��m���7f-p�u����|���1�:l��S�)�?:�z�p)��th��v�P����W<D���6Xu�o=)�|��ƴ�_�h� y"!!+�� �@$��3�@Y��?�g��Q���:���ʎA#�dD:OK?/��*=��Uo�w�,3R.y]�E�J"*�cyt[��
�Q�^�;Z�M�jE�0�'���oTm��ރ�s��G�������_�۷�����̽+�+^����Hq8GT2�dŐ(?t��9F�=8��8R��ߩ�����W�_�`���	�gx�}]�e�Ο�O��}���i#c�h��h+��+������t)�J&��ӳ%��~�\���C��HWg��q>��=�������w�8���Z��M��B�� ����WS��5.�/˟�~��(�L���ef�Rs����E���?oz\���Ub.)�O�G����� h'|��$m֖q ��(�����܅G�G_��*n���:�����&���J<0u�L�1�X���K(�~a~���H������nB%MZh»m�ͱ�.��˜ �%��Y�"�fY�d��۹vA�[�]7X���a<���>ܓϾ��̤�;������hC�O*�:����m4Ry(g(�ʎ^P���6�g� �[�R��XFk�X�ȥ���Oh 6{�S5�K�pp�ѯ�=aɇ�SC;�h�H���_�jw
6QH�t*�4%�!�&tPq?`/�^��lPk*��ԇ��ޑ`�F��U��Lk#�J@ ?9���I͋+^l ���Tw"_�
����<=h��G���jĝeǺO�rh��Xc=�(;ʫ
�F���g�k�4��V�Z���[Ts�rEB��c
��@J<��� ����$��c(����/����B���k�����7�7�3�r��T��+:�R��6;�/L�A��*�(y�P���%h�T�7;_F���@>Y�]������s �K�L���4�"�Z�_�.�r�����h��"�N�����;��M?�]�
���(���'�� @��K |-����۾���P�r��1��?_�� �M�z/"d\���-���uÅ����	�i�6��'C���c`�7�Wk��xe�V%J��C(�Ֆ��0u�gv�&������@��9��%�Я
�:J� LB`����ǵ���Ut��Ŋ�^�k�� �,!BM�����A�;�T�R���Q���{X@� }��$|��v+җ���rZ�����Y�&����+j�F�?��!����6�YmuT�pT�!ډ.#��W�Y�E�`�&!���K��ksP������ز�쭴y}�p|Qe�k[�a�Y�4�	|DX�4�`�7DM��($JΘ�#O�8��o��0K�ekh���`-`q���uS�-=P������f�H�H�� i��n���ː�f���9`�#�T�0��O�oA���*���V2�]K�.���b���1UZ	�s0��ꇍ3�'�Z��&G�{����߾A�X-=\c�c�>Bɾ��~�����wI��ȯt>Y�U��L�k>l�n���x�ѩ�h8A�ё�^��3w)�Y�a��l�ۖ4��z��.��h͌���
z8�� jY*��5�	�Z����:���C��"�r~��k	�s�/���b�'V:&ٞ�w�kw���SEH�3�Udp9����G�����=�Y��c`M5�σ��P�
m��+�*F���E�SkEY��w-�3L	�����k�cq}�qp'B??J޹��Q��sd'�]��Q�&����<��9��香�ꅶ�:�C��mSn��W�{����~���c ~���t�؞��B��zޯ�_��c����4D�D�]P쀡��_�"��f
'��mHI1&�]��9_+N�(��U��5��ax���,�e�Bϸ^�*=Q�E��5���d��f@AvN�>`e�ɒ��bL��bő�� ��˰S�vؒ�������.�-D}h�"&�N��6}�@��^��0 D��q霞�D!�}�8_��B鴛PR�|�q��a�,9xf��z�K'h)�7�|�-�s	��=�Y�m���%0t
�Z8���xk�6���B�)������y�|��x̢�]� MS�������	����1S�Ru_�T�ê��;�i�YX��`�2`*�8�e5�E���k9ӻ(��nd�)(n|�A�%w�A ��S��Ѥ�M\	�iv��!�K-��xIw�/$�P������8$5ߴ�.I{Ô[ɉ�1�z��ߚ��uk�|�P��u[��b��r��S�?���ԏ��=������_�la��?�C����ւ��fzk��yA��tGt�!��ܵ,�؉�h_�R:��3���Bc�>�����@"�ڿ�CQU{���s�W�K�F���;� ��е&�D�O��-�8��/��� �e�	dO��>��Jy?j�]�a��ż���?��w�@X��q&�6Y!��x��I7���uX��g�x|��E�r�V���`��G�
M7+z½0�C�x��z(��������U���	��f�)�\�:�EO�y��$�t��7��2�o�%�U�sd�{�	��ojh���-x�V4�J>�j�F�dT��.7��Mn<���<�$��W$a*�uD}�<�I�������1�͟ �į�YP�������'���#
nР�!h�g�0���;�,LC��I���8��	8�$�ᶌ��2�>��PC������7�:q��-zRҟ%�퍝@J$#�q��qʗX��7��4Tz6bƤASh�08�tH�+�K��H����'�fc�t,z��	l�Ɉ��l�Bu��H�]ecf�J��:�a;;qʾ7��ŵ�^1_�TnC�
��f^g���ǅ� �9q�v^(�Z� :������|�w�w�Δ#0��4�X�h��V�uN1�����E��#ş=7�R/]�0g�MD+݌	��$�J����a:�лSK*�Y+	G�h��u�U9�}�q���?/��&�̥r�����$OJLi�ؓCK��5�m�3EKR�_���JaS�H�r�V�sM�I�=�_�ԹT�÷fΊ���!���&/8��B���ϳ��XhL��A&y��5�����0/���!�}�K���,�.� O\��Q�E�΂g��:X��GC�J>��,��9?#zZ���bI��<�e�:3�9�z�c�,k�LH�c_���Q����n%d;Dq�d�bBWK�W��F�ÈQ���qgپ�{�����N.Ն���=�J�Ku��]��+{�Ե�3s=�ި����A�ΠR��#3!G{B٭�rC��(�vЁ��f:.�Z=>��WL���-�WD�a���Gyu9�o��6j86\�`J\$ULCG��;����7�vw��6�����md��-�S��>�c_#JvE�X�n ̖u��>�(h�Jf�9 �����v���U�����`�{��c�4G�a�}��������pRƔm;|`��@4�^��|��`r���\�
[#O��wI��1���?�[&y��-co�1] �3�g�a���o�)`h.*�w��J�CH|����� 9�:���m�<�	�ɡA`���Mw/��<�L�i��&���1�{�s8��J��~UgK8��j!�~��mVp�_�uF7�?��bf6��|_߹��b�q ^�r� �T�)ۑ|�C���L�7�gB��c�J*�;�v܃����I$EF	^����Lod���6�G�O9��_v2+����)�?2{.��}�����3�C��Ǫ����o�:�j�Iǂ�Iu�2hG�T���O�wB��]ߎ�zK��&�Jx���Kj��B2������ʹ]�:�'I��9��۶�/
&��S�=2B����D��pp2Bи<�dv]y�-�V�pOQR	[����-a��u
��*�˰3Q�yjW��b�>x�/sԫ�e����s%��:�Av�R��+�5����K�>�t��������o!����_O1(�P�'��3Ҭ2�n��0K�)JhYR|��F�-PpxS��"Vǥ���2Y�nrn�L{5w�닔p�'�b�I�)���`��2.�3�����9&T�dk���A&�%�l��x�R�D�Η����4��4V���=�����FXb��V�<\���s��F@�y��v���B�Ȁ�D��?�$� ŗB}�����H=^ k*����0��x�Ǩ.u�,Kg�@v���p�W��߰<��%��������"xH��'|p���	N��N�����^���ۥ�0{�n	�\��֮'w�EXy3RIϒ�&�\lΏ�v�=ܜ�k��4暎Q+���3x�L�Z�@%��^�[� �<� G�a)�f��?=�ѓ������1ĝ�{��tf�0��u�lI\麃	   �,g�+�&4񏧯v+=���ܨe�MT9t#T�Ԍ�A�5��d~L�G�+})���2�%xYMT*/(�:�������J�:��f[~b�{�����m�}�w�3�\کH�[���rm+4갭��!��1�� �p7v4�<����8ʩ����de���fY�Z!8��3ם�qv�o;�Iy�o�f��h��r1�'V��+#8�gæ��t�0Y��_>�8�'ǃ�f%�1���.^�4�w�F� F<�=��=D�j��i#z���(�j������"˰!ˆ�:X�o��V����:��NH�8L;Wy��>�k��-iw͢?���8p���u�9��W-����a��bfٛk0'��"��5T���q͠Ѩi�pڴ�keJ'�y����%���{�֛���ok�%iR��,
�.a�T9���1�L��2���@j�_��&;��7�r
a��\�%f��e���B�2öWj<A�p;�����XE�.K+J9:�T�e���'�� 2�Vmey����_MH>z���i���R+�?r��� l����G�p��'����i�|���:e�SN׶h[�mxJ��D�����C��
��脦t�-�`���8�ٶK�c��55��iT�{�ӵ���C��ܸ9I_}�26[�^�{Z����p��-oڕ�v�G҄0��l�̇X]a��}Ѹ��7leZ� ��-Tox._��u�eWMI��Vc���k�\%FG�Jx8�Z��<K���ɂ=m,)��[`&>7��Б�P�I�ݾO��ݓ��YhI���2W��ň�B$�ߤ@m3�������o��	��	R�\W�0~p^��#�]�F"���b��'y,�u#Qz�f0�&���F�� K�sMJ�`��"�+���d'��/<8U��l�Q	�lH0��c
]�-U+��}��ԋ0�Zv���iF5��)k���2�;8�*�ކ$~��3����p:1��0\�@���SPۭr ������N��gi��8p>���짦!IY�&�� vnl����=zfĪ6�I�0���;�%�7�-_�O�'�*M���S�Hd�:%�����>�TN�uy��صRI�B�im@��qa�+1�ץ�WD�j��KR�2��dѧ;O~"	Gono�ʡ�� L1���=B">���G�;<ɴk5p�M� ��䔵jRZ6+;�	�R�i�t�\Ս�����h��N֍����/��}FGc���1Z���	�q�ˠ���D%&�ܓ`�8��=50��|��7��,&Dq�A<��)ܛ�nVA�V~�6�'�[�U�͇�\(��m��-⬽��NJ��S��G��g|f��H1�A+mP|P;����]��o"�o�Y�q:�%����W��H|[���F[px5w�Y���nʷ�wF�#+�(������4�-��ӄYp^���kK��N��JZT��3#�f�B��Y�4b]�$��﹎��uߺ��M˨�%��"��<\�`.�`� ���jz�z�*aؑs-���R�j�aukor0CŦ�2�V������������0����Qp��8�B��P��rW�n�;���;�4 �7��$(����Qf��� �>.��a�p���j���2"F+��� PO	ʰ��'%"E��j�����*�ބ��:`H�&��O�p�BrGl��Y4��'�D��i(����Oi�p��_|������3����k��ZC�(�ܺ�;<r՘N���_��1�̡_�fZt��u�	%pP������u-�5�
����>n�r;N��\yY�+�2A{ygA�-(	��B�d� ��E���g3�W�o�(#�\�i�/�:���.�T	V��ߴ���C�?�|F���ֆ��8�@���f���a�3=���	oX���L�5Vy���á��w*���9�op��/>z*��y�f�Z��!rԅ�L�E4�Ɏ���).�)r2�O����D�8��0��O��]�����h��0h�a�6�ʤ����g�F�r�w�^9qS�2��IU'1<{�-�M��G=�Ec���,Z��>�.����1���>̓ʫ�ZjOI��-˕*4l�<�Dc<2ơL�Q4"�tէ���0�3$�[4�K��-��,~�+��դ-Cf�[��3���Q�fe�٘$b�,�L;%;��ވ��f�l0|(t���+��h�G耯�+a��b�vߧ2��s..�_B���s#0�%t��� �r����e~+[Rs \?"\����L�A�P�$���1�rK�*rhM�($�ބޚ��s�hN❵9����=C���Zs2�j^G��$�4�.	]7cp}4[�wHqnYx+9a�3��Z�L�(mJO��R��V�f��$���5j������N]�	��ϵ�o���vB�Q<NJUAKIOk�稔�7m�%Y��1�#i�'��!b�J�yo�L��JO����E�x��׻�����s��r��p��Q�qbNJ ����&a�R�F�3�L���d�#��h�Y���C7�]�aX��}�8v	~�#�['�!���5����υ�|Zn����<�E䎣-�ф�@�;k���0PxaN��/z q^+��JA��r��i�n��y a�9)xx(c�9,2��L(Ƣ�uq�Q�3�a�٦�fX>Y�*ju�*��a��'֔�Bo�J\�����4��AG�L�(y;S��5W	{�/�d��eں9Z(���f@� ��s���3,'~�O`K��+��%4���������9a��csz�X�,�ֈUg_FT���.�>b^�(��o�����g���0T*�;D5!C���"��p�oԟ�!���X*�Q��F�)xP����u7���/������8����e�^G�u�!/1����T�)�55�x?j����6í	{
�\��qw��-�� c��11�B5�Ll�&	oC�]4D��0��2rGb̓��e��2��29�%C�+�V�o����~���ƒ�����:�3�ҬW]�f����E�\[��U�:z`��L`�5���F��I�����,�4Q_�Y'��Ǭ�U�P-��+��c�H�c�|�tz�.��ⵝ��x#�c
^?->ٻ`S����Z@D�h�޳��Q�T=��E��r���Y�r��.����rF�'��*yʥH1v��T�x�����/9��ƣ#u�?Z��
����I7���[��ro��v��R����S�Ϯ,�%��R�V�&H<Pr3�b��]�9�U�j�z����Er%��$x{��	��S��M5�^��S4�t�x����n�H����k���	���9�|�ŏ��P�B���<ZI�,+`�M}�yם��1T-�'yK	)�`��5��Ls�%�?}��R %<p$x�<��h=��U6n����.�Fj�"g���`2m]��x��v�C�)�_pT��z����\�@�����|<h9�l}��,��I��V���"t����7��^@Q-��,f���G&��G�����n��n�by�]���Hz�W���p�y�8����}L	��/&�u�t��N��S��3S�������-7뜘��� ��$�j�°-���v7�'Y��l�u-߰�(u����������u���\�'Z�IJ����D7�zkun��_!{�00+?fmtEv@n��(<�W(�N$�ڟ�����6c	l���Leߐ?��f�*Ͼg{k	�#��Mb��g�~#m��=��+V���`�\a�8� Ym�
9�E�<N��A����9�o��&�'�����Z�~y��d���Z7������a���˰a��(�#+
a;L�4N�$�ğ���*�c�)
BD[�ݨ�LCdq���!��%N,��;�f���F6��O!l;�ӶA1�5C�_�ϖ�����D��\�c��k)̯�rr�Z��c�#��蒯��mn�����k���'\���Ms��餐J�f�	�7	�u��`SH�*h�ᮃ}�s1W������=L�����G(&Z�&��m7�����`�N��MID���|�o�#>�Z
�MZ�ߓ���Q�]�7#0f�a����9�2pԶB����7lI\�0�E˙��F��>�44�^Q�=�W��\�=�\|���4�O ^�ދ0,�X����'g���36Sۃz����ު)o��##��X�"��q�P0��e�k�g+i�;H\+�A�G�)\����� ���x���;��WPz���.��\��8���B]__ ��H�p��@ O�\,�%���wC`�u�+���t����H���I-c�ū3���6z��k�oV��*��b��M�Ǚ�۪���+u�����͝��;G��_4/�����X�df�w*$KȨ��f-<�q���'dRܽ=�L�K�£��pS��@�٩!�	Ȗ<ۡ�J��<BT"6Tث��D<@U�Hg��p��9��SEv������ѹ�Z��%�b�j��\�����1_�rF�	���lXaC�5�)ͻ�+�y\��V�4x"�;3�"�����}��q�{��/Y��K��~=�i~A�@ѳK�o��?G���un��z�������J��7�tI�|�/�x=s��%�w���������C���~�i##����,��@�j�����;���Fu>�����5u����$�����$tu��uH�&���}㍖L����ΡU���
�Oٱ��*����+�Gӌp� ��A64����.��U賫��/���K;���x�6�q���p��?v���,�F>T<�x��]'�	Jհ�
�h��@�1�K0:�E�?��dR^�6����F7B�����X��\��'��#�5���GI�`s�^S���ʑì��gc���v�ڥ�T�L'dڴ�jqn�-����/o*�!L�69&b��AN�#�A�fӌ%������#�B�l���U'M�ژzYi�8��]Jcq#��J�^��z�e6߂4�}V�����V��/��l��_�&��Bk?���M�f����
_�_Jf`eB��xE6?C���~F*o(6$�~t�ʐ� @�R�k�.����K�/B��*=�	��?��nzC�4PםA�.?���~C�i���94�3y�m�*��Q� �BL�W��\N"�Q1�0�S-*}O��ƭ�R<��d���L�]ԇ� �fy�}�M���Z;Zҭ�٥]x��BJ�4��g~����N�0���篙#i�o�>�Y��4�B�U�g�s��9�6K��#�����s5��/��8���'��>��
|�8J�O���tR�A��cg�zʔ��5׃��%x���-+i�=r��ٌ���b��N�΃����R<�@&K�C'�]�n{	��4��@�KPr{���������"��6��j?~�9���D^�r;�l���MW������oe��A�S��0<�7�#�k�4��1�5�����&�V����2�qz�Vb<��?�������/V]���M�e�%"�!��UB ��IԃȱF�<��_^N��?��|-�cbK�����HF{���)ZQ��֭P��a<�e�r��x7Q�g��*��M���ΎH�w�)1vGs��W�8O�Qsbc�g�HR�hrW�rM��C(gk =���V�ғ�K���Qa_��Ƕ���P��n�IH9#�|���~Sݮ\jw���Y'H���$���� �a������|G�.ǲ�Vq�)�*#B�.�/3/)^ͽ�z7)Q`�!�,�(O
�ǙB���j�^�W�tQ��Zlj6�ٰ�t�9t6Q��)P���E'6���r�^G�Î#��o��x�{��ؕ8̡Yo�K-Su�]d�	`�C��"c�o�)	��=��������f���	��sB��ږ�������Z�6U_9�0 ��^X����!�p����66�W�e׵r��!�&������|��o��J�)Ͳ������:���n���(�SUHH�c/�TL7�uOS`����&�(���.���x���}�5���~�K��a�L�������آŀvձ����@'+��wǹ�䦜M�j�N��ˠ֮e�/r3X����ڹ<��Q�XG�0e��ڧ)e���糼-G"�*�>f=�w�i��i�C��UD�^�ehj��HN��\@�O�E�6�~�? �Y~�<�^���9��[V����j�	v�%YI�*�$��ӆ�f�M?x� �����4��5�6M�#�홟|�ge:���;9@궽�c�5�g���t�"�r���}�;ODp#7�����z6xF���l���b�@�[Mp�8;c��[����g��_�7x������U�/L�U���D9���Ǯ�YWl���Lp��׼P�H�MW?5����_�,��v���P<�j�i��U����gm�~�pf�;��]����E��*쉦�D!~A�i��LlI�->d@\�R��ё*��F�b'gܞ�P�-���WKa��<�&���,������SNa~��H��Ҍ� �f��rHs��NYxg{�Ɩ�PiA\����.�,FO;�/��pvt�	m��˟��ǔq�E@o��j����&ϱ��/��^�*�-Y4'��پ���i�<U�$�>	�����r�o�����mVa���'�z�������H8(��ukݖ䱠�g8�\-���:���)TO���7T�6��k���(�����x�>ǲ�4�����4+e$�3"�������t��`�HF���_�XvM�*׶tU��f$F������Xl��c�1�)�hSi�+#�]��!����Yy��t'�)��]����9�i�́݉��0�5���_,e55�oR��1�f��13��G�p�=�Ѷ�z�w�������0Q͊�����s�(��M�\gN�˭s�j�3���d�V�gW-r����EE�rg�DW�P<�����ĝ�6x좏Q˾���IA܌��<n�B���ux�=����A��ޙ(��zx��7P�� ���x�
�pav�+��
�Khx+a:��cy���aT�:ǜj� :[VXo�xPZ��_@�V�����3%��_���~�El�|�=�V�~���8�V���{����m�z����u9��*��	m����OhX"�X��Q��z�7����QIܪ���;"�q�#���q<d���,�*�@~njzљ��C��c���6�P)q��(5
#�-ʾ���ź�z�>�:x�=�0�?u&��w������.AB���͛�w��%�N~x�߲_m��VB�xS�}~��AT��9Y�j���<{�0`c� ���D���[ŕ���b���oR��@D8�{b�,�L]�!���$ODMAyr��Q_�gJT��8\u*�<ɵ��8���9A�`��L��(a*m��r~T�j;�9�� p��>l�b�Mއi�̦��fO4�dt*����r���o���u/������wmk$j���]I�	ݧ��$r�t�0��.���A�T��r�~���Dɷ�pj9QomM�����3�.�O�:.�%%A��_�b��.��M<fl����2�{���+��~M�03�K�n��N�8���Yx�bU��g�Y�|�<��yt89��V׈\O=iɪZ�	�`f��Q���;�6���BǛF��8��r�V���ے~39��5��p�,d@��o��jL�r9��^�Ҁ��g�g'O�����{��G�����B�-Q�2��Uԗ3J��m��b�ċ���\T�誅Y"�%L�U\Q��b9UM��2���T(=�S�i{-��bE���΁��@��8l2�~�7��'�Y"�e��my �������'���A��ɱ�pX�k�w��30�b��V���]��7�!���ܪ�xVΟG}}��7~ĦdJ���b�	$U�Y҆&B^�m6��E����aߵ&�P*$�E[�T��pڸ*q\��ud���HY2�P2�3%ye�۵�c5�_�P���_u�L�s�Gi�J���ZP.,�� kn^�C!��'wŚq���(c��<�{YV]Rv�Q=�o@��6���nք������l��d�X�9�g)��J]�����+���F�&�E֭h+�ǂӕaOE=��L�}6�g�"ȷ�8\/M�r\i�w�Α�nv=�&v�]����p��M�B��J־�Z�;���z�sq�ۧw��R/�)	C�~.�:�%*�·v/��p�Z����&��<!o�É�l{uj�5z�����(�9s��i0Q�{�0=�N̟�-*D����D:&����0���,��c�g�[>{y"��_"Ƒ�g5�Y��Ԍ��W�15XP��=N����k�B�)���-L���Bۢo�?f��zs���ܣ='�����Ld��_�+S=���¸E㟰?�E*�V��o�1n8U;S>��D"/.,cC8�8�Ҵ���w�B��)Ȑ`���@I\�����ݸ�9 ����I��B8oH?H0�'� BZn���>�2c���ʋ�T���"�f����՞^��T�ٿe{�7��v���+���i�\��:�������E��DAKG��O���A/�8'�c�`=H�E�`�d�μMu�=����(���"�K$s�!\*����Y�ɤ��3@V#� &�]"!If7�L�m}]!V9�h��c:-S����"G�Tꀇ�Ϗ�oc;�4o�T�Y���	i���0a3���(�u���_�I'��ߢt�"�:f�58�:�
���i|������_�?r�K��a?0�0>�,��š�s��O�nEv�45J
��"������{j���U��e��ſy�=��>����f�fu�����A���Đ���._�mc=I(�ż�2)����l���M^M9� K�,� x����m�<��zV��!W����^2�o�9[����>-�B7&Ȗ.��ʖ|��;� �M�OJ=
�Z�6]����8���:27s�D,ʄ��!5�ʫ�D�#H'a:B��^I~sOs�f(Q�`����fǭ���p��n�xl��p_j��쉵{�b���es�"P��:�������ܯ�u��h�_"�o��6�x�c��� '*�>�'MPN�bZ�>��]��/q�$3�O#�@�ڱ��Dql�ڿ�ЄÖE�,����Ί�k�"���[�`�u��4]�9�FbC��/@���W�$G�v&������>}E�R�4E�;�����{o�J�o�1�ąg�tn�1zF�B�4��0lɾ)(f�ӯ��j}���GM
�B�����HW�k���>�9k�$��_�m�tt��W`��v�˧4P��J�� L������E#@/��(��_$��(��з�G�Q�{t�$��	/�Y�vC���Q��fi�aAŽ�*:1����7�W�����r��߱�$���X����.<�� �̻��gbI�A;�1,�ĮIC�13�_a�EK�?�|������3�v���i��+3�f�UJ5ձ���oƧ�z�;�AtKPѵ«��?;�a҈0Ͼ��@@�-�L�g�K,
e�b�YPpgBE������ޤ&�f���\�*��s�f����WpVN�4�Y ������g~�`����"�E�������wG�R@$S��g���w�L����:�h��|�GB����O�V~�h-,�g��I�~��L���|*xZ9���^`�:��� �!WH:˻f���%�1��+]c�
f��>C%#*�򔰾c�5߂���&�#�Ɖ>j>$��pUq�LicI8%3?��.(J����Y���U����k����߂}�n�#�@�a��z�����aP�0OXᅲ������i M�ڝ�̜h���#�wLЙ̕��l���41�ަ?�ғRA�˨0�qQ�n���0c��ӟ����!z�Jh}d��`�,u�aC� ��Hr�W3/� Y2E��������?�۠��x1�D�$bS�V5F�j����v��U
R+��~�?|u*�7Y��=8T���b���{z7�n�����	���Vsc�)V��ײY߫�q
K���볉�}<&�mS�"~���f&�m)�g����&�G�*���O�������b���Zs��#l q�G�]8��J�\Go���-� �"�wq��
\�{�.ʫ�Ө�ъn���N#�ps�ڊАH��v}_*:q�<�Z,o��1sY;?ʭW��i��n�������킩Ya	��܊�� M���/��^Qt���RopM�kA9͝=
�3��
PB��A�+;��ʃ}�_V$���@��^ais��R_v��ҰC]6��
�Gq-�&G~
�KTWō�V�6��IO��h��
�xRv;i�>)���k�Փ�O�]a����t\]<���,�����-1��=l@��y�Mq����ä����|��C��H����9�
c�Mr�e�`lɠ��Iv���а�r>k��W�I"Ȋw2r��9y,���!1Q=-%�(�?/i�B�RY��FgQI�}�N�\����:0�IM�g������]�p�~�Xy�Ȣ<p4�'�1��s��S��:�rG���G������K���gV#C�N�z�p#�֧}�őʮ2G��ͭ�^�1+�2�D��g�X�y�)����6��a��De͡�#B��\;e���`�v\cN��Q�&��."l���Lt�'D|n����ߏ����T�:*���p�H���.�NI�JQS�꺕�Ke8N���ǅ�,V�x�8!�0�De�MB�;��`K��z�O0�n���JI��c�m8�p��6�N���1?�QGF���aΤ��O�y���z�6��x�/&��(�5B���t7��^�E�R�B]�����*�Fwn�إ�,;���}? cޥޠ���?"K��^ܡ��|���j�%��l�6쿒Ֆ ���fϜ�0�c'��U�`����q����I.�0�u�<�C G����5�u�I5��t(C���\G��#�=v�r�|X(�!\��(�u���/G�ˊ`�p��)IDy���?=O5��?�WAx~[�R�WNR�&%~�˟K�tO��WH�N�&���nh�#��lub����#g-��
Q��V�1���Ȩ9�ْ�\Uֹ��_�d�] ��e}f����Pnn�9�㐠�p��1]*I�&.�O�e��}E�Z�9��3�I��j��iv�Z�H�(�8B�d�E)�&/, d�Ŷ;�*�O�=wv�z�������O!�M���s�"Gݨ���i1/x�� ��C����d��"���%S+}8��d-ɷΏ��I�7����T-�7�/,�!��
0�ga����玥���$�0�S'ƥ�*gN�-��Q�j��*���ukf�U ��FwR�͕lF5c��VN���9Ў"�+K ���B�}]�����c�T�F�oCr�w��F՛�����'Z�B��u���=A���U8�N����:R[���@�4�Ym^Nv�����'�������oA�P�i����/����U�m�?�h`�~�Tj�H�%���������elLl5Y��Qh� ��=h�������K���n��BJA�m���9� �Jt;���'{����~��A��Oo����5�
�kG��u������9��_c�6\���th5$��d�m���Bx�����^�;Skq�h��Ё9+��kyކa���6���� �?��Rz�SF���P���J��tR�y6z?���1���ZJ �D��!�u����A��H���^��_��b*̂e���I�)#�h((��쪘�<����x�/�:�"Q;�N�Է߲<o�H��B%��?����룒�Eg՚\H���,�r˛��gf'�ʨ$[���/]LC�G����#@G����Wr{ 5�����q�����Q�O�I�A��8;G�x���,�(Ӝn#�$x��X;Q�y)���W>�R2�}.����S�G�m@����X�_(�����}N�L��_ �̌�٤w�x�{8�)q<���������s+���O�V83J���O.1����&l���X�%��0=����[�*��O�
�2����;�,ޑ/������v��n�B���h�"��(O��2� ¡B�{,9�B ��␹�^O<ۨ�&[	�FZ<I^��v��(�΁U�`7+(&P/��Y�8(I��&gg+y)w��J���(���ޱ$3��	�K�J>��ݑ*w�Q��u��aqM[�2(�Nu	����C}7����f��h�RA��$2WE�Z�>a�Z�5��"	����u�N3�l�k}g_�uT���¼������nEٹ����a;tþۓ犟r&\���gc��]���x�Ri�|i��։o�z��|��!�l�k���Su�^EX��9^B����6�I���#���9ڲ�'�cpr��(���*R!���C7��T�^������8W�~����(���>�eJ����!�As�çeˉ�p/M����J���k�h��f�1P�����X��K��Dx�����#I)ڽ�l&j��[����c A|L��������6f�v���Ҳ����V�z /������/Lr|w�)����^��LkX�Ő�2��Y�3�����oBV Hc�_�M��7b8a;�:!(Ї���ߢ�N7pg� 髷�j�&`���҆���EU�!W@e§d�f,؅_[���;�y�@�$9��Ȏc�|�8RS���N�kar�񱽙Y��� ԜK�
gu�\����e~�x O�9u�R�7h���q
.��-ͳ0W�i���8�����p[K'��G�fG�����Y1>p���M/Z Y�%�7yN9�N�Z�8r*��J�+�ȅ\���%2�����c����X�C�[m=������hɅ�P��׉��G�RA�͟t�� �e�y:G�2..��v�kdY���4���� QbT��o1���*��TSnC5��`&$E }gX9���9ǷGǟG�tlh��c���>)�|������ ��&�<���v�����Ǐ��|إ*�a%`kH�)�1j��� FtJ&xu}$C�1M�%�]	c��~0I'���Qj�����+�D��k�9:�ߕe����*��T���|-��|�J���x�F�wb7�JQTUt�"?�ZT�[vJ�L�KP
��J�U����B�pu9�L���m�w�:ƥ�U	M�즩�+�T�ֹ�����]���:�s������54&T&Lvý�4K6zNeYf�SC���柣���g�aq�8,>{�frZ��W:H�n�3�-�&������oُr���TPNec����/��U���`�P}�� G�����鉐�d����M#(�S����MΨE������}
V�\���̝���'�Y	1����6m�Ա{�(.=VA"�)�٣�yG
�ڧ�-�7p���A�������+T�*!�ȧ�P֝O�Eү��IH���B�v��jT�`}�Zj� [���a=�!,��VS.�c%���ƀpz󒊥抜�"�Vr�U>���\�Բ,+O��v�>d\�s8���2�)��l��sbݦ�!��h���{]B1L����b�?�G&)�*f�x��2)t07�'č��ىQ.,/u�N�z����+��� v,!B�md��:1�pF���.D%��	6��p�$��h\�P����9v���)n9mG��y�D��zK�	7x\֤�GotvܤXx> ^��r��ޔ����C�H�O(:K��)D]:F`��5IN*b[��/+'"Qx�)߂�A�e,�|;o3��{�M�<Q0�t�Ke@�!i�l$Z7��M�e��ߺcb��L������V+��M��F�9\4Ըe��8"}��-�^J�g��A�7�s�j^pFi���y�%/>c0�W��]�ޟ�0v*�֦�~l�|���n��_CBS��k0m�&��D�kQkۗ��O&�����Q�I|o�9��a
��*��ߘ��n�
�bfb��/��6bM�Ç�f xp1�.~���4T�ϲ3xjXS��l?��Y��I�m\�|��҇V������ѷ�.��J��I��4�nY��On�-�n�^���.s5��0
����(�\=�~�j�/A�')����5}�"�q� ,S��^��n��K&�`Iy��O��]n�k�/A������*�]�2�ht�����er��t�J�S#��n�\�:�y���������jC�LF1q	�G��	,.E�6.y�Iև×b�N�jaB�d
n�m�2-�j�[������i.�R/�>#[��xVBC��UR"�M8��'�W-��
�Ղ��4b�+'��$AS�l�
�m&��s�{��Tx�9`�H�����9���ȭT6w(q���SRQًw����&ᯖ�+����y���,k�����M#)�cu+bɍ�4����,�E"������	�������h��=D�0��C���Y:�ұs2��� �b:���ťD"n�S"�Y<�a3d�:�<��d;�K%z*q\�-�Ͳ�=�6:��Y���0�#��h(�1�x�z�HD���X�	�k���������탃˸�|�Db~#Y�:7ᙲa�1`VC����&Y�8�M��э���_�e�߅��R����!d�L�µ�.0�Vgg�l�6�p�	��ݞ:��G����º]	��J�U|PH���G�B�MR뭚�5���	�)�(�!����A�=U�-z�������M��&�?LX��Mk� ��F05w�zTW
~' (O�?=V�C��3��x�7���(���γ�`���Yj��R�6���uu�<����`Zv6�vT%ٲ���h���m�\�9̝95���Z3�mU0z�3ug�@��@H-��ޡ����W�r�3C�x��%�x��\^S�h�+��{�-���k2���F�q���jp � ��?��;Ą�]��rb�Y�4ۦf)�s��(�>
�D{��_#V@֟����pk�H�����Xy16����EGD�h�Ş�U��a��#N�-��;!�������ˬ�³��BKU��#ۻ���:2��p=�Žmm�Z�g�	��"�S�+�Ms�5}�.���Cĩ{�rW�����)�U�Ӯ������X�	�2yMa�w�(��P�bR*L��D�fd���]�U9���RfYd���8qh*�_|l�z��%j��B������n���	�)Ǻ�)9,p�Oi ����dh�c	c�a�)��fs��^��r�%�Ք<�>�m�^-JjT@�bVË9H޹B�t���G,�s��tzC"�$p_��W�F��*	TT}���oG!,_�HJ���O{w�]��]hA9[��J��8�7<�������t3f/���\�oo�)�s��o��;���nr,j[Xwx�!߀W� q6�:.�zs�_V�[������� -j��V�@��z�E�i��cf>Q�)�賱��VrM��ߋh>���u��^��J�gN��G�z����}�j�EE�@�%9����H����a5`����r��� ��Μ?V��)Ӳ��]�Za�^>>���<��8��.��8��g�{_��/�V��:��6ˋ��LtG^����6�Ј�tM�ed���h�������}��1����<�V
�����}��-�g���ߔ"^K�_�ӭ�KD�hM����/�(�_NB=�X���@�{��Pk���A�eHn�k�^�E�x�p�5d2�{z��h������G���`�T�z_H!TR�?�nz�،y�j�%���B�R�����T���grGA�[6�������Cے�+Ɲ���g�pa�,���R��9�DUR�U^s���d�y[��٢N�?�&~�jy�aaB���۵:z��E���u��z�+��	�\�τ~� �I{_2E*�i˃#�=�s��0��i+R�|Kd��<I��1�Ύ�7R`F� '"���3�_cm����I~���֥ ��"�E�
��=�����f#���{E�����~�0��o��*k3'z@#�$��p⽘k��W���`��3qJ��.f�n?�7_��H��`I�奭���JŒ�
�eǅ���W�>���:'�yD��V�5g
��w��`ٴ�2��6*)wǵ��1��dT��E3F�����@�Fa�*��W����m/�)�q� ��
��<�K���$9�[������	o
F"�r���q�t�Y���>��Y����e؊
��KIտ=�a��gĸ�%�F��q�;����ʴ,C�[u��
<��4e5�ȡwA���d�l]�
��Ŋ�!�?Uu'�����e�.[`���pۉ��g�=��҉����&�3�� @����!A�-�ES%)�Z��[��B�]�}uh��$����h-׉���ﭛ]�
[�~{ga6w�0�	`�mҪ@)���y�b[�g^?�����������y�T1��L��O��	�uO�{}�G	�R_9`E��hE��p�iH�Ա)��Ig/��b��3�(��Ď�_/�>��Y.�1$�dI��X��e���%�3��BǞTV��<��g;ᴀ�
{4�c� �ʐ@b��Xg�y��7kL��ˇuDE�u]���Hv����2��W�\j#=�zslԠy���WX��\�&RҤ�*��~2�W'r��9�ʳ��M	�mi�=MkjB��=�Jp*=>t@SY�%l��{�Ӵ8�	sօ%
O*&����4 �~�{���wO$�k��!l������~� e4I��1&X��u'��Ճ�1��rEe���t�̏�<��^�~�x����Ո\O4��'B���[w�捼م^�`(��;��+Q�@����H���_��_������y{4�_gw_�c�A<�r�⎮*�������e����AQ��Q|��q�Q'�?��^-����p�7o���i��wI��<�����	O��zp�0�uC�)Q���g6�2O�B����k	,������/�%�I�g�t�3M�@�S̤�Pn��M��2�ŋDx�#�-�T����<�M�,�C~�[;h�XD�_WF����-��\T3FZ�!��VBՋ��΂�h�d�ؤ���a"5�RgI�N��ܿ��E�	�J��Q��2�Kf1�e�ş!͒/l0nm�9�ߋA�@f�z�f҈�ZE�x��b�ܠ����4٣�.�/p�F+�j�2;۽���CA�jK�H�忾��Ŀ}��L�S�b���r�|��Y Y��(����xy��d|��B������b���R:�#$���y^����c��g�r���Ԁpe>�l�r�4tw�|M`5��N�o��I�w^��G�$�f��A' ������a�Xv_$v5g���9��;����짒N�ke�YS�'늠:ڪ1H��{ý"&��2��4��E���I��齶�uG,��`�}�t{R���;a�ъH���OwʕQ
�l��F�{���6�3�z&S>XD�{5h-��*ܫA΂wLU�Mʸ�V��C�A�+*��l���Wo�Z��އq�������G5�ۡ�v���$0i'��}��(��3�D�;i�O��+�h�A�дn�B��p(vte�}�z+GN�ރ\u�`M~G}��3�'���} I�H}j�M�}3��q �������4׮�e44���� �}����n�٥S�D2.9b�0Bф�1�2L>�xHZ��Xk��̙�oc����S�k�.�ֵ����n�q
��{�k���D#�7$؎�1�}�rD7Evz=� tQ�v�a����<���80�_�<�8�>*�p�D&��cO���;�Q!���N2θ��壇ϝڮ�|����w��m�PO]:�X�@��C��᭜��~Z�]�����(R@��q�,�<6K�E�o��E�ђ��7���Z��T$U�a�FcG\s��j�J%qw�˨�������[Կ�}����	C�Ĉ)���EE%�6ET$S��mx����05ĩ~��� ⑬���]�Z+ �߈�}@��������$�){�L�Z��&;�wڟ� %���8K�`����ف�g�Ҁ�ȩ��-ь*���O"
��.�̴o���M�4�)c���_�J����«f+�Fm��]mq�[p�?�]W��,R_��T���K����1n����9�� Q�u��G�R$g�G�g)��q]�7޽I�� z��BV�'n!�f`��;�eMQ��8)�$�"��6=%�:�(��]���MA;#��{|��VO$K@��v{[M|����6?;�gp'�4 �7&��P���r�+�s�A � U ��У�X�.z7��@���Ю!��������%��<�sv/��ȁ�o��1<�ӂ_���_K��N#`�
Z�$⽵���O5pt�1"i4p����~����k��%/ �J��'�����������vp�aOz��Wd�3͏���c,������h|nޓL���~�\�x�Ŕl�v-���B���hoA�fd��B�#��n��^�\}y�=!��.����a<ޠ}��?r�W��*QgRz�<x+:��Xv��W�������(�7�H�z���s�lTT�J�ܰp��LL��S·��`�aL�����lr�i��@�r�aа���2yW�=꾌��n_��-���(�؟q[ю������]3���o�(�8�����W���`)�Bl�y~������p���22H|�$��EŠq�fXL�}�քf9UZ�#F?ݯVK6"���ࠧ���t�b�{�>T��W$��R��.�ᬀ%A��j��~��_m���z�[���P��X��Z�����8���<�[�Fx*M��%�#�^�Diݖ����^��ۋA�<,�Ǯ���*����)�J�.jf��\�����^`�v3,����o��?	K\��4s��ҎD���5Yq�!o�?�@8ⱷ�5���H�����*�o/�����zD��� �#�  ��C�N�6�yQ�_�%|����S���S����M��iX��o���o���R��� i��2��4�+t��(ω�u�|����^fT��|���nfTy�S=߷��cM�d�̈gv����bU:v�,(��|�r�K��\.8�sx����l�������M�t���������\�Fڟ�S�"�M���[d�z�)5CxW����Z�1!�i���L[Ŗ���T^�uq�P��
���j��Y�_�w�^O@��k��;�[���D��S�Yd�'����᝹{x���_���a*ۋ��`�Zڪ�a��Sb�>,[�*߸�P!����d�<����lBa��Cqgp6��I�1���k-	@cD�>h-���@6�#�u^��� �'�?ǐ֚.��li�{A�V�:�Q�tЁ�vXt�@�Ҙ����*��p���Q��o˽:e��mB�y=�^k��
����$�diX��rq#�����U�C ɛ�ߗ@����|� z��Al��N0��?���px�g�G����Ewg�s�l@c_w��خ�I⻕a��BܽC�0wХj��s&3�Dl�q��������/�g�s�C�����]�9_�^R�UB��@� ��r�p��Y����a�#�H�g�L^3�MU�u+���\Y���¡�y�]u��	~��vŰ	zՄ{�B��!Z�c� i��E���3�lVl�`e�����O���TSo>���)N��͂S�����=/�
kզ��\�n'����d$�%f����W��Ep�B�+�3�Y-����dt��d]{7�������cEY8Uވ�Rڛ��LI��/_�3��"ou��C�@�:-�DB�HX�����l�s7՝��l����B���������h��ܖ��"I�G�-M\��d��V\��8��l����>����>9������vjYؙu�;F��y��=cj(�	qߺ�kj��.�y�9,Ĕc����zb�g���rl��x%
*�FjnC��%��	%�쩀�)�K��"�;l���H&w��fM�?���Q��@���51���l<�*zVB��-q�\����vJ��6�)������ӯg�f�d��4�/
Q5�y��y���A��2>��Wq�(�	P��QL�cx�V��\y|�ѓ�`�Ңв�F��@���"��q0���H����j�Z��aW}C��x��ŀ>~��r}��B���	�˚���E'���T�=��(����e3���Y�з�D��e���L,��_���B(�}_?��M�s"t���]EM�b<�7&��%�_h�ڋ�2mc�	%5���k�{A��c��3.��Ƥ�ZyI��2Hk���_�{(��G�=�~Q� �O�c����# ?�c,:/��TS�2#ڴ�](�L�
4�6����, �?'�@q���,=��o���K|�mֻA9a�L��_Ԧ�< �4|`<Θ���[�lVю�Ԣ�4�0.�%�MdĶ&�Oo�_w��*�i�{����p*f~��%3����ʘ)I2E��m'�k(
��u�S��a!��J8uJ�*U=��Vw�v�-�nkA�����g.�W�M���J�i����2�c.���怖^��Y�����}X%Q6>��U%?����toD!��J��pR:�+m�C-:x���6c�U�pzR���mm$�+`䦅�&�G����7躈��X�V��� �Q<#X{����{ލЧ((E��.J�������}���ۘ��Q�EZ,�-�>��|2R}U��X����Sp����32 
���H��B��%��}ﳊt1Me��ǝ���LG�yHX}v�i&��z��Vn�b5M�>8��� ��GB�w,ݍz 7�ϔ��0"���XR^M��S�����qՔiai"�X�s`ֲꀨ��w��U��Ѳ�l(����JB ij7t���Q�0�u6���F(?yh�⨘B��U]���G��fg!��e\�E�<��[�۸]������,��*��H��3*����2i�Z[& c��S���U>�:r`�A��p�$�$A�&L����U�HG�8A�u��[&֥L&��#{զ��n����"!�{?�R0�4�;�^4gh��' ��cվ���y�XZ�
��BLk��U���]�R�Fy���ʴ���_oj[뚸&&R�1�iU��sJ̄�k��M� ��ke#�����|��"�vh�j��v)�=�\C���P'%�G�2F��ه��p5.g{��~��;�L���-�0�Zu�N�k+�Q��i���KS�O���~OQ���b?�O���1B#m� ��*W��S�?p+O��W��"�;?8�
V��&`��j᳒��&�8m�U���ɭ��j�O�9Qx�z�˜�d�eDw���5��rl��#��XÀ�yw�A��pu1�}�=�L���=dk_�e:�ފ���*~�M'D���X Թq�"�A5��)�?�S�V�Ōh�v�vs��Y�Ɛ�yn}�Ȍ"�4�!�l�5d
��1x�lU�MBO��n�%J�൧��tȤ���e)�+GA��@+@�n�cН���.��d��D��k@$�����JX9i�	��Ep�I�sَB�TKd_��I�s䁸8��L#�x�o�'�vĤ;��Etz���<�|�?l�g'���S�����9a����P)�E̋7����0�A,m|Gn$4忀�q��	;�x��`�ԧ�ql<�����ii�ˎ�+���	�I����7$N�U��]~`��c6��5i�DD~ۀ�
�d$��(�9�9K&b}K�/X[~:7G��X�9Yx�M}ܺt��'��{<v��x\^_�