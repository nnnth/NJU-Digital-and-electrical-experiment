��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��h�S�L#��4)��L�6��b�
�U-Go0 �
�A@B�_���av������U���"��-Qéj(a����p��3���T�l�Sত��RHx[	|��r>_�7h-��h���0��CɠXz������l�;460Uаh`��o��h�R$�`�)}��_j��ԡ#E��c�a��@�u	Q��lO��ĭ>��X�J�)
�D$\�m!w{�����1ͮ�֌�4�Il�õ𾵁䭶�vӪ�^$&ʠ���x���{۳˻���	>�?ü��f�85;��R�K��6i)h�+u��s�B��ɉlo92M�P�Z�tU�ұ�5�R�g�?j*θ���S�OL����*O��`�6ȁ��J���}zo��*k���j^� �"\J<�Mُ��09�=�t/�»dq���f�l�P��FI��r�!n��3ߝ|�=�L�f�Vn3!U���� �9|J��h��dپ���A�#r*���+Ep7�i�}�c��F������1еN#�6�&^�(�O3�o~�oZj�a�{t����W�I���3G�,4�ڐI[�jx�0Mf�0�)c�ܺ�Ф��w�a)M�|�tn{[
��#v�$�vH#�v���B/ɲ��][��$��[tfS_�^���&p��u'���}��].ߠ����˺��\d.����dT��[^o��9u�qt>J]x�F�F�Y:zʤ�g���< �
���#�n/��P�FC���
�C/g�5�,���.��N��D`�۝���:yԇ�kƹ��s�?h�\���u@Y��x�]�T=!bCe��:��
�5m�\���<�<��@э�1J��>|s@�[l�[�?���㘂�+���R�>R�L��,�=7)�{�M9�����3�kUW���e���S|]a�R,��o��#���{8�(����E ,O>��р'#�n�=uo����s���Nu�(���_C�)*�}�3�C�'˘۫�K��|c�*EH��ǲj������`7뀓��pI=���G�V�û�-��UT�$��������6A
��w���NB��ԪL���t!jL�M�R��M���b��v,�yNp$Qڼ��I��G����e�ͯ�/Ӄ�l~Su�]w�R���Z�����o5�Z��[�-POٗ��,V�[���:�Bc�X��ŶH
!����M�p2F�-˷x%�7=�����s��Zf��	8l��H5�n��P:��#P.u��@��ϓ����	�����黥�������`	lnG��Rɼ�ׁ2)#C��-^�c	�9[r 1+��,� �s�	��fž�<ƒ���s<�Q*�,�2�}�3&�t�	��6t-�(Q���ԃ��+8�o]���c����$r<���W�L�(!�'8�e+\����<tbbO���=uz���*��}}�D1������ב��%�������/_�\>�'}�%t,C�ߞ78��9!�k+��ϑ�j2��)q��ټ�$Aˬ�)9����3�2�m%��F!���?}�6r���l�>�1�tF}�iC�M�+T�l��T�h�����HO�y�	\W=g�n��!�����j�4\�����0aU��E(��8f�	c��6�u���Jصm���OzR,�J�3���٬���⽶�5f��ھC=��`���Uu������G첏ƥ�|��e������5��C�8yO�Ұ�q�Y�F�����UDxf�E㠩��⌊��̍���wPpI�o�����z6[�u��d�C�%La���������F�:eƚ���<ڧTS�"�[�N-'0�ծr;�7c$�ׁ�˓�b]'�B�])�#�{x$D@l��d~{[�~�����*L���u�S_��,,��~�iQ>�����L?�{
�Z�A$�Qn+n`X���G5g��udJ�����}oTQo{E�(�o����*����eL�w!������$pCp���{��KnP�I�y,��2��z�p��OCZc�~���c�^1���4���~N�} $���y��Y�_ ,��.����������;8�=��)l�T�=J��A���,�_ B$d<��eF�
�(cn�u�ث�|�H��^�u�������{�U�C��ne�X�8�?.x�&+���1����ئf�W_,�G��C�	 s�\U#�����Z�hN`
��?,o�>e_;9�Nq�S�� 4�q�N�(PWO���x��>�*������@z��L�G1a�93�f�hhC|�GΙ��Wf�];���L-�<����E~��p�'�f�7�����bU�3�=R�v����LIu�ȗ5��c'`��n}ݲi�|d/�r�~���/,6G�M:���Z�nJa�x~���e6�K�9��W�Ÿ 6��'�N`�
Xz���5�OŜś��ap� v������^����^\�V�2ZmZ:vK�^w�s�o`AFfz�<�o>��P�%�[����eP����4ө%[�ΉS%�L}91Ar�H}Џ���]�~K@S�N@R�7�̍�����=�5A^ф��;ʴW�&���`�g����a��\��Fk|�R7����Y��M�	���:nx��ێ�2�6_ۛ����~#Nր��8�Nh�0HZ�qT"��ɽ��u���;����[R�J��!�5'��>a��������/�D�j�jM�>���,+�b¼<Zz���aن��c�S��yx�7%RFE�mï���.޲H ͵�-��������c=$@ V�T�R�a:��|�9p�D׊�F+�zIX�!��6V|�H3̩4���S��]�c�޹��~~�!���=|PF��\i��w���n�7�.��^י7�&�R���d������A������tp��_e�>���$�Vd/�{C��Hdn�m�5�z�j	�'�����-��	�+�֕�蟜��>��J0��m�(U���,�\a��� 8�룅�ج�(���Y��bc�U.��q�'�=�E]���̞>��p҂�ص��/�E=���~`��x���bUZoPD~�G�HWW@yh�� ����6�쭸�5&9��`\Q��3%��T�g��7ׂ�$���'H��J���0iM�Zp�g�����������[�2L�VHI���Є�)�F�7���[�.���ڵw��4\��'T9
N#׻�8�v0�GbaD0(�E�/QBz�t8�=~V��L�i�qբ+LN6�/��+��@��z�5�錎����l���;�ʟ�����T`�"����Ȧ5i5�s�/�$������UĪ�
i���K��:Ư�OT��+(�%{�!��U N�c��`s�ݛB�mRh?�R#�`#SN�nU����ݿ�����&S�.���#L� :����QtI�r�ޡ���	���-gM���4�9�6����h _> g��IM�9|F����1����S�O�i�I�����;��#�n�@��nl�p�D���7A�����$�m�E���'���@�_�ө�<M���=X�[�V1j��=]���Di쨄�x�+]n��>֔�������sY�w���h��k߸�	z�t���e5 �j\A!6���Z�5�/�#<EwL�5�d!-����wV]Q-?l�*��|#�Ir(kn�ږ��-N2u,����_O^Q\tGKm0��S/u�F�<+�ٙO�5@H��LC��qc7�6�i�LF�a'�XGk�m�!��1�0k�6~���U������兛E��hkT�s ������V�%��bʆ������)ţ�%�H�n�Iဃ�\R��X/3�hixP�ŽT����9�nW�1'?�CZ�r�H*{y?D��M|�W:	��+�+7���`6��Q��S ����:H���2�sU�7��9�l;���ud�:?&Vٻƃ��1��Pp����R�E�!<v�Zl��p�8d2�:Q�kM�]l��7�Lp�w�/<�EA��@�U.�)c׌P]�PlgM�x�N��7^��W]Ώ7jҲzM���:��C��B�cf�.���ą��Yʅ�1|�>�	�oj�n��Вw�.��Q;(��sd��p�*L�[��-�W�@c��2�@�sΡ5j��s� ѧ!W;�%ՍQ�����<�7LR���ZR��j��߂*K�X$UsC ��H�6v�A~̤�i�*l��������kjKE����:Ј���A :Mq˄o�\���C`���*��n#��٘;%P���v�g�ivS�ް���l(g��X<̙8��|M�HlGaf���iEw���XIeҍ���E��������s�A,8�}�� �}�[>��ѭ�2�ٛ�ȫ֡}f� ���T��I���!O�ؐ���>9Ø��n7 �-�b��\Y���f�Bc*;aR\���p"���4Ǭ)��V��kB�\4%�ե�/'��� iz� ��d9�:YGi	E�5L-n�h�̃4������c�V~�c�-�:&ԧ��š���|U�p��]�8:̶�򛗃�G�߱K$�|����m�B�����-�Hg?t�� ��6�nT�iv~i*���F�0(,�\�����_B�%}I_\2f6�!�2h�X�l���[BuO��F%�,���Jݨm���|v��V�����x���Z=�rrxl;��߷h��2}��4��$R��M����IBL�FE�2�:�?0���µ�*q�7��3���6 ��ر`EL�"��.��˧��7Z��Z�:�i*�c��B�+���_;��K�KV�>�G�"����,4=�S.�k�k_���4�b��fΰ-ZF�������NR|K�7���;C(����m���>B�B-�ZC��B>���lx�f�?R���#>���V��Ig���ߺ��]�/���%b��vNĝD�[9��(Bs�u4"�����Q�L%J���Q/l�>��v��7�9�,gSG����ݢW�$1�L�F�[��(w�W"�X���+xR�gX�����S NVaH9��kps�E�F�eı�^ �l=T&x�?v�1 PP� &�vg��:�����J�B_2jQ�[�G���������/Lq:����gs�k��	��tc���@���Rnkި�<L'j³� ���ߖ.e�ש��v���i��+L�}~S�c�o;��x����lSG:B�O�Ud5�zB_DQ<�u&��!��̫Ϧ�"Ry%����ɜ��:��]L�P��t{d������!)�$e��EL�E�E�����Oh�s�
���d�ٽ���M��6F	.�L���5���7n���2����}Di�u��GP��U�Y0#����H-j�=�Up���񄚱I�ta�#�>W�����y\#������t%-�q�ܑ�}X�obv�*|x�ͨ1<2���/�cN�l���3#V֗�:��-�Gz��3"P��������n�B9"��v	6IO�9J�#]ט+/�~K-�e�������đ�,��ʖD����ٷ,�T���f��s�����.��_�R!���qܚ(��^v� O.s��W�k� �'��H��B�D⎸#ݰ_�#��5p<�wп�km&`��KP���"�T�1�¬E��Oʶˠ�{nT�Z
�>� U�sI�������uK���2�0��a��u�v�[z�݆ӡ(�H��{3	��:G�ި���Tt�;P���O�:
M�^��������3M���u3��g����̾^;TԎ~͠턵�dl�<W=CR�M�U�q�>4cy�0�ڻ~��My(���~��\�Jl����0�2��?�<�mt(dd���J&,ް;z��U��_'���gM	�:���v2k�4���Jٴ�QDí_�_g&Α���:	7@7Y �F�p>�[C8���^��!n�΀?��'�Z:³�� �<ˬ��I� ZkLc+|i�(�݋)���d�#$�N�V�����C�YkFy���I���I�y+7��G=:�r-���J�ؽ|����]�L�LF�#�y��4�����4@Nj9��|;X��%�X��D��M��Y����a��j�|��Mw8Ic0G	�TR8f����C�'�}���ǟt:��+ö^����](��&"��28��G�ѷ`{���4�6������"U��׏�`���o����Z��)J�C���������xc�����8?;ڢ�~���.�:�M��K2�[���� ʙ��姥etF��\s5[ ���g��bl0��l�!H��T�ۙ+�'�*w[��	�����ӽǗ���N�mM�%�Έ��=��|�i8�3A)4ߌ�ey��W<T�&�X3U ��X|��ŵ�WH-��jL��U$�&M��)�|:�I���x����S��~ǜA�_D=/���S޺�)˿X�r��<�p��|�K���������̷�Jp;��-ԧƒù����ض�|]|l3>������ȇ�������Z7,��n��b󁬪T�@��	L-�K����3#��q�!��]�n�fW�5��Ѡ�55�Fd��A�W}�k�(�B��<5�`A�%0�C�-�3M&��`���J#�ݜ]�TY
�����d�� &|^Բ*<�ķ��#�h*3�M]����|����O��!��M�M#���IzF�J��S�!>����@�W��+r���$#:~�EDɵ�eQ>(���[߮�qS�> ��9G�I}ʍ��,d��S[Sq�j��?�1�*��G��z���R]����!6D��t������f�8 l<�ow1��_��G��+H6Ƽ�	�R���DOfQY�L��X�h󬁊>��4��/�`�β��1)���t��@i�)hG����ݣR4Sh	�T)b����1�waٿ�{j����Jh�l=-�VESz׮���>�6M�I�j"{��OX�� ,4��d��T���W��B�����i��Oy��M���d�H��6�Nt�I�Mbqs�n����L�U��y|^Zq_�>8�ﬃ홡 �aeؾ�|�o�'��İ�����i�b� ��	د�%�� ��K��-d��>v�v~�G;��bƴ��M�wP=1\�υc����[o�F�~z:Kݎ����V�����q��� 5u9y�g�MݭbWa0p�:r|/r����cK�轚Ap( ln���'� �K0��ݕ2N�E��ԯh��s���'#��Ɍ�l泃T^�c��X��T�����8�Kt���Օ�^w�A�#��e|�Rʒ��PT�y��ב�`N�'H�B�M�N	,&J�R���D��?�Q^ܕ%���[�v;r��I���c�q�mC ������5m�I,�S�>��ߗ�8�c'V��6�I�8�;��**�Q����`?�R�GÒ�'|�����A���s#��.}��������!���Ke"B��.q���Cٲ�7��Z�q,�]+�/O��2�GE�Kx��1W��hy�$�C�8a'�+r�
�׃H`�ᤞ-�����TF��F|2����TP��Z��t؜�P�����1Qn���?� &�6.&�XLLq�a���o8ƵAR#E]ӊK�gQW�\3I';�Z���@?�e�i�!2qj�0�]�#�t��$��i�C��oD��{�8�Y6�ҳ�~�=}tۖ�-�,��WQ�ju�ǟp�댗Q�-�K�rҮ���33iR�_�ґ��fC��ٲ^�{�F��M�9*�K��ť�HIψ(,Q_#�e�L[��%������ݵ�Z���剷���s��kx3:X5�L��ڈ�kӁ������,��}mT3Bu�����W�?�/ٺ����M�i��E���^��r��t���[��٘�>Y+-ò�\(��曩{�]G����ꎘ��~l����B��8���4�|����ȫ
���2�l	wsv<����iht��)a��km%ڼ�1��ѲK�k^�2��>����2j�u������7�L9�<���+Y�=���A�f�>9��	k?"�� �+iLW�Q<��#%�
��*D�F��8���`����O�#=36iP��A���pR�!��^�. ��Ĥ�J1�t�����n{�0����ٙ��S�u���#�EE�%β�Y'wX��BI�`V��x�)ǜ.q��˝���ҕ�����)ݫMw�R�tC�Iȵ3� ̹�p*�@�������K��ʬ#����t3Z:�u�4����X���DlQ1��yٮ��`�͠���@��8�7!�9D/���	������Q��xE�@uԊK��Huuw����^p@���{]�-۳��Uw�'~���.j����xև��������n�,�#[�zE9�'�}����kĽ�qYbS�9)s9�����ԫB��q#�.�!_�եp�Hka*�F�F����vA���%UT�wi��X�y��i)�m�����9)�[_�ʉ��):#��Z(_ނ���Pț���x�tVñ\*I�9WMqv���9������U����)mሞ�ӂ��4W��SPY�TM%���H�ڑ�*