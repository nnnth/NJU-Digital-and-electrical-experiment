��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{`,u@=.P�.L-|�̯�	�恫f/$�mv�Qf�~�{���,���[� �dwk}Cp�dp��Oz+��x�R�#O�W��	ӓR��SG������k)��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��\=@��쿿��6k?�u��O�B���gǏPt�4b�j�T���N)�J�����Fh[j^���"�!-;���3����⤝}S���ؼ�DG�U�V�&��V��~�=:Aa�}\���.�S�;�Ɛ��w��щ��:�c���K�]���{�J��݁~m�\��4�g�T9���KHi�Gv	�j�sK�����IYl�殬��:���!ȥ/!J!���wWr_R��"\��ү�{��9f��1�I�q��p�r�t)��b�Ep�2��h"J���qa_.���"����maM�>�h<�������J��Fߗ�vk�#J�W�"7W����j��@�i�͒��OO�mG�"���b�Av�vKx�T�.2�j��	��2f9DM��@h86)�Ǐ �ƖD�-�"3 �KO�� ���B&�q;�:��ŅF6Cn�wF �w]��,���$5���f�dI��^���8 "{t�shy����R�l6c����$4z����l%+�Pe-w�mj.�zX�DF�wڵ�K�:U8�"�}wNY�� ���,��rf��ؖ�3��(h����R�*�5��6��7Z��x��NȒ��&��4n^�o�~���(�P+�=>W��\���83����O8H���{|���K�Q�v�ޤHko�y:���v�>7����t9ï�����WB;��Z
�bs�b"�O��ڴҗ�x�'���Ε헃Wy���+�y�ȧ��1����	���04�M�A����>��3L)"=o}��[~$,li���*�UY����}-8�����\�xqI$���G,�4*G�ELb�\��,M�A���7����<h�3���C�h�d��J�]���"����l#�8��~v�+U��[��I2�En�<Һ�H����qj�� 9c�#�C��!<6ّh��o����i
	8w��Ӱ�5�dV�X���(�6f�WYb_��B�*�R����|�
hq�%,�A9P��^1y�LM(���+�Q���P�<�Bk�R�w�(A��%���5�e��u�D�p"2`�*�I�xfG�n�!AWP�u�vEa�+���:�֗�/n��ʴǬ>m[���K9���@z㼸[�?F 'e �T��J��BY`�c�<V뺰}},�ǌ<�N��G�%(j�i����ШqțsZe�_����y�C�H�C�u���l1ͱX�ͲxD�7
2��"�uTQ�ej�щ�z�S��}v�^v 	�� (I.�#T�+rg�S�����}���f���#�s@������)��{x�#Z�����C���Ԙ���S^y�ć�����)cϸP �CZ���z��L.*�Ҵ�@	#��"�$QKNmr�7ޕ�5qg_�SLIDU�L��lq3z��&,������l�gUj2�����D�o�D��
Anz,L�0x��^��
NG��̋D�/��S4��
X�I.�������ӈq(#n�|� '0��`pͯ�6�E��u�0K�O�)��ߒRhW�AT�B�e�aɬ�,���y�6P��ɕwt��CZ��ј�_,�w:�4T�=�b����@�xsr�g���d+����<['O"xt�%��: ��i�WԷ� �\�k1P�P'���0��!)I����%�I���t�3) }':�De�
�~�t�� 9�p}{_	�q<�D��+H7������p@cIe�d�Pm�ҁ)�y��I�0�{5),��9:;'��(�I)3���ƇP>rV��)�FF��&����ޛ4�pt��(	��dx�۬�� v�;�`eDC��K]_�v�,b���~&����_x̌���M<vڲ>�mϖ�� �?�} �3�ۥX5�,�k�R_H�<<Eǽ*�5���j3m�{4���p�S���KH�4���ͅin��|\�2'�8���qEp8/����QߝGuzV�yvX@Y��l���ۛ�ׂQwR2��}��P�xW�?�y^���m�"a$����[toYCN�m�����O��� ���v�z^ߙ;��zQ��G@|���ǠP��LI߮L���i��okw�zkyt����kt� ��7�/ȉ�cjl���;�O_�.�� ����iEq`B��
lAxmN�=��Ƃ�y���cS�<���t\&���d�V�S�t�:������Ѝՠ�wϔ>����A�m
����'�ׄ��B_z$[9��
6Z9�@�1�S�_��ii���>���hqg ��63A����[�����aB�`�@{���X#�L Z�a�w�:0-�rO�x��^1�:�4�.����hJ���Iu�V|�.�t5X�~�����8D��9��O��U�`�)`=�ܤ�4�5�`6P�{�������^T�m!�/�,�r�˄����6]�k���t�˽���]��(y���7����È��c�:fZHؘ|� 42�oN���r��,�M{�a8��@8q�,Ɗ7��o̱�8T�P�/Q�S	Z���e�_�~$�gEo��%F���R�Dp���%����Jx3����p�{���h�
�G�f�x,���|�vI鬣����le�n�LQ�b!n��� ��?rl@)XK�?��E���|����
�!,γP��1<�3�O�y��s���Z�+�!��[vFZu�)���S��zQ���b��P��J��N3˚�X9RQ�3հ�­�ċ3�ὔ~��5��Xa���f�y��:�p3c��W �d�i����MS-g�mP��8U�"A��̏���_��OkAd�c�����z�!=ǜ�%�	�@^o�jg4 �m-%�Y~5SG��1od{��_ �	��S.%�Z�kS�_x~�ݺ����"��Mbƍ��ʞ�#0��5������9#�(!GOP��qא���V���s?��h����2�_�]�eNo����ԬfL7b�(U��'"��w�ٷ"C�&+z���^?�%O����B�I�-�Uz��� _��@���=]ph8#�ً=�|c3��n擴߰m�� .7���hx���eC_���2n������jE3?-6�Y@lڻc}���O��r6"��~�]�tnӄH?>���4�4.Ў�<�hHd�q2��k��i]s����R2�pJR[��Qو�
��3��"L������6ߘ�h�ā�4�X,�^�n�&�8|���²v!� s���Z��;q(	eO��>,DU���ܡ!�bX�}Z�g��I1 �4�q�W�;�$%ԫ�P>��
w��f��O������!%Y� �ԻQ��=<�7-Q�c��~K��Z/ �����jt2s��߂���Q��&�=���6�t��f����K��DarsLgJ�V��#5�"K5�h�����T$rj	���W[]���s�]'*�;la���z�kJd���ḟH3�:sޏ���g�w�����'��m�/{�4N���\ǯ�Pv]9�I3j4E�@�#T!�0<�f��d~wl8	*��󖌱�"�h�9��
�Ȫ6c�?��a�@�M|��0�[��7M�a\��j\�q�0��M'�e\>��m�M�h��PD}����2e�w��%�v׏a)O����U_�?�WV����>��W���*�.C���\>�e ��)7��K2�:����_�=�C�LT2`� 6tÃ�����ͬ�w���.�j��#���a�x�����
�@@'�o`z���g�n�B�vE�g4Ϟ_^�����Fn7���ZD�b=�B_����x��9�l�4=���b��لgÁ�.h��e�H��ۯ�
a�/;�yvQ�,W����8�6��������:sG����3��Z~:c` ���������N�J�<��봓��v�05'��󽼞^j-�<����,=(	.ob���*\7gY���C��;e\2@��5�n�X.�}� 7(؛~z"��7!�����y�Y�߼���I�ɡWe���8���񯪷B�?�ixrFR�ų���>��ޗ#Z�\�(�: �E�����@V�~�L6V�1�8G�Nz��R�.�w�\"��.eg���;�:�@i�^�Vn�lނDS���⤌��Y_��2�w!�Z�)%)��~	�_�9�P�ք���-HV� q�֔�()��)^�Cs�.٤�}�����='�H$��,�se�D��Av�4ы�����cT��*|��{�+_���av
�w���~Ŝ��"�9HZ��Ri�Ena۬� ��ϓ��<pA�~��<���P�/A�۽��#�Ve3������yK������!f���´����]�+ߋ]|(DI%I=)��.�R�p����w>v�������B*��q_�OƮ1��v��a-湖��>�V�I��K�R�_қ�L�2��Y�~ݲ���Q˹��8;g6���-l����aFw�<�(�ێz���Z���ɯ
�=��L�$5��'��w��!���/��M�̾�<���o`�'"�+2Rf57H.��6O����i�����~aM����+1!�E�����Z����
`�����4���Q?����u?��W7P3�c����N�4U�)�/�kV5��§�v2��u�����?nT�?���+�j��/׽`^1��
[:q�#?�-��#������T$F��H,Qn��@��R��Ė�jb
���5u�$�S�M/�1jV([l�����i�ԧs��Զ�OǛ��Tѡc��W�.���o�v��ň��KO_WO��+O�@�yL�C��m���,j�DF��N��EI��J�G���>�(�_�c�����}�[�э�}[wb��A�d�Ŗ�"�(��;W��9��^A�d�Xt:�m���
L�Wq@ͩ��{�����u��(E���	��Ӈ��Gбa�h�JN�;p[b(�>�8��n3 �Pg��i����*ZR������B�s����tgIG]`4����p4=T�Y/�wm�]C�U
J���r�Q��4��LXz�3Z�8�S�Tz_ּ�c���/�^�[� ���9	��$q��I����C��i��H��G�6Q�a}FC�UÂZ���h���_�1&���y|gxG7^&p5���]'k�o�i̟' Rn��)S��C�a���,���7"Ǝn|n����&{*3}������C���U�	l�0����3��\6V�½�Z/<�>��$'��ɚ�s�.�֔�3m�xM�	j�$n���!`__9�#�'��D��+%�m�S%�9V���x<���u� �j�rk	AM��N�}�ˌk�u�d���}��8��x�2۱����.@�hS��I�Z��b(���;�5��0����1�O�������]���&�j�	xT����+[�<U�:U+Oa0F�XǛ�ȹ W5�M���8Q$������=��� P9��!�z;e��M��Ѱn��2nS�$�,?�S��B�iF��m��a�~�+V���y��r7��˔͆������,�N9�ũ�c!�l�**?��s�ҏ��4��y��Q4��������u��/�� ¢kj7̓uB�P���#�M?z���2=i���V�� K O�o�;��A��`��J���Z~�:7V����� ����T]�(��aHV��k��ɏfk>h������
͠�#�2���ev��� ��k���6�Z�KOzr�=���/��%p�-��,�:��R@T�H%�f����,��#Cd��v,	��.�4욧9I��#r.H�SKD�/��MEH�H�	�?�8���菑���±m��K�����.K]ΕN��:��1(����;EYRrb+�;�H�EJv]��\m�	�o|�}Z5Y�x����[Σ�Ʈ:���M$Se��	��P2a��������!�y��>��{��Z���s�t٤:!����[�H��L�l�m�Nu>R��dq�L�i��<,�6<��7�ŰE��l�Q�1]H�I���諮�VlW�I�kdY�A<�z��U���Zh�1G�L�%��D���m.;OX��Ҡ����/�tV�Ŕ�R\�/�=£.=�Y�N�����'��;�J�èU����/�u:l!��p�S�*��=y��P�ܾ��i�$X����C���[���~�-p1ùG�\2�L�pߐ����z�4���ǉ��ST4D̓F>%�ʗ��zt[Hn�7>A��k�N�^}?�#c>�Z���S���;}
��>�]�����s�� A�{'4�e���d��ՓR�����A�v���R�j��2b<�=i�&��Ǻ>�&e>����k��@/�E�b�����Z�/�[�_E%Z��TR�%E#Gb��c�P�+��i�H�+��Gz�K�J{��;@�&&����D��]�ߗ�H;
X�k[���rN���pjw"��A��p�>��P%���.����zb��a}�m]��}����������q�S��k�y�CgD�3L<V�]�Y��y*z��Õ�0��b�A��T�J%�ݝ����+�A�ؔ>\(�xZ����8�������lê^\T>�$�	lW��06����~Lr��m$�
�W~��0r�;��Uh�R^�4e>�"�d�=0���(#�d��z�~ٵ�r�x�A`��p���^E��H��qQ¥y5'��G�j���L0�O��^�9VcD����J�
_
���M%�q�����7�dUb�pȆ�s��ݏ��7	c�]F�����A�L�A��2�U6?h�}�:K��,�,�������!~���}2@{ U�bUW� #fo�t;+6PD�"G�W+�RH��")�Dt`~�k�}<O�|A����+]��tOG�`�q����`<k��v�2��1��Y�v�����ە�җqLCddo��I9������ޠl��TX��o�X�����ʻ��V��!	��%�4�f6�0�ۭJ	6���/ԲX�8�~�]����z���:��؎j#lݨ��+�e&�N��|���G^sz#IZ_�c׽?�]j�U�1���#��wh�
L�soų�=B܇W��.�m������\]�Pt��G�*���I0���g�R�B�U���n��~4v�V8��}~$l�E9B�m�ZwՔ�d��UuX�V�p��Wz3ms�	<��1�4��X*q�į�t*e��	�-�v�y����~׏�Hs�GY��2�<D��������x|�=I蠎9(�p�k��,?Q�=���	�9T�$�k��U	�bY���T�3!ͭ��~Xy�,�6�e�̾j�,a(�>C	�C�baI��S'�nD�I`pq�5�]��&�l����_�Q�,ş+`��l� y��s���f��+��V��A������z�����&�=����\�<s*�W7��W]6��z���#����aLYŚs�d}��b��Cmcs	z~�����{|���ꤪ�}�6�
{O}�Q�~���ۙ��ǂ@�L��0|�L��g6�x-�^D7�G���XB��<#(,��|��Hݦ�n��k^@��
v?gh��onQ����=�W��gz:r���a7#��8�����|*\�;(���O8m�>xţ�a\�B�]��\����r�$h:Kw��e��V{��FO uu�'��@�&�]�`Y�����0�;��.�ٹ�h����<����*>M���(�A�t���P��%��F��$Z��c� <�^ٽ)��v!�1����o�=�z#Gk��jrM�gr�tTAсbc�j#G$��� PPس3�:xmh;���3�&\R�2a�+�||�3����WEL��gΠ��X�L���U���%Uh=[��oZ$j��+щ��ڋi7�A��V�!�c���Xc��;�,ǲ�N��=0����
6��.(R���*E�`1�L���Hb�u����8�g�D���;��rh�a?�Z7N�6��\C�.&�P�7ҳMY�God��G����M�	$��5������ 3I�g����;��-R��-�ER\V�^�GLa�����K�����,c����J]�P�e�mp� �{)og%Iݽ�,�㾥CT*�������q** CąJ�+��N���oA���nI��`���*]/�<�QgW��ŧ������m�gU�濅���nost��J�G�Ex1��H�_���ηߣà��Q�&����YcS�I߈�ߣ���'?`��#Ki;�
 7_�:(x����^{D�op8(&��J9V�#����*��P�y��-�������B�3��x���&H�z^������塃;��l2��d&R��T��M��_c��U-����R������P��ZťAat�R�4�H�/�D�w"L�zb�&� aA�H��J*R0�~�ʘ|fI�}�^.��0��V��V����� ��Gw�t�R�=&�X$���\tnT�V�numl3�U�4]��pl\X2��XQ�\s��J'}0��;"\r�߇�Z�+�ۭ�fS��q�eF쒄�3���ouJD	֫�OA���rߚ����6��a�΍��w��(����j �O��ʿ�0uc�t@;%9�.����h���X�p��.1��)��xS$���	�R��U�9�����.}%)���|L4;fK͎�7���6��4����)�e������+�Ȏ7rw�
��_6k/�A�����2���"���C���^̥����TA.�ul30�@�K�n���`��?x����#����s�K����\%�a*�^dC>Ɂ�O��C5�Ę&�6��IS�?��i�4�Uۈ��cZ.%mP���N�t?o�3�#xI�d�fR���2w���+P��fl㲐�o��S�C�P.�g�CeH'��h��am	�L�U��V��n3�K�]����Ks&�d�0��8�s���<���]"�+{#�EX�@��@�����/ aXo�i��F�#u:��Jꉌ��̊��\ܻ��;�K��h�� ��)�r#� 0#R����)j����ʻ\�$���8	���X�#}�|�� L��~�: �0y?�ۢ�n�	F�N�Qd\O�����e��;��9�g���"/��O/�g��lqÕG5d���c>����B�mJ���[�˾,�-�>ei�Nw��8��M!k\O��۪�}�E�M5�+�(�3{��_��)<�+PZ���Ī���v���;���r�<���d�E�-��-MGp�
h�������.��B���K�E����/�ѥ�r��1���-& ��0(��US��C�<�ʛ��#o"����+���>X�;�xR���%O�6Q�+Ga�����<%�d�M��Ɋ�̎��*���H��W�M~ߙxƢ/�EdV��C<�ġE��`���+S<���}��~^�h*j�z��nW���P�.�q?�^hԺ���ۭ$�a�A�d*Ŷ��Jvqc^��o[x�A�eQd�l�`��v������C[��`��e��n�Z�i�5�1�N~\ߚ��ڵ��>�p��|ƃz�|�YP���0�p����e&�S+����I˹���.���)���p��f�4�&�$���ugL�RN��ⵌ�q�}S�vU���fa�}��Y
�x���L;�_�����a�LFJѲ��"KM��Ӡ�kzcJS��X��L��ϒ5�k���(�{�3U�u��7#R���/l��P���,�t��l�G	_� 1a�������P���ʛ�Y��qC�%�xc�#{�C�*v#
�ڨ�(���/KP�a� �ؑ<@���%e�pUd��Oę�?q��c]�Y�v\hj����U�J}:3]�_��X�ћ��ԽjQ�FNq�igv�eZ�Q�ӿ��4�k΍�.�����9�}B:��;�N�'�j0s;��kI)A=�<\����`Lk4������E�����|`�[p�Z&��7�i��۝;p�w����@r]��[˦�r�/n�<�D��uA(V���U���Z��N��P���៊ 8�k�����2Q���u)�9��c�/�(B��䁕�J6@f	r&2"^��8_�D��@����x�^-��T�`O���vQ<W͡r?����B�h2�
�U�����+zG��d�FF]?�S�z����q�4"T���c@�=Ʈfɨ!~x$�$��Ys�M(ܐv�����V�NBY�m,���|�m�Ϳ��L���k�?F�y�/{7�4�P�G���-�5���C�f�w�L�[��Z�`�j0G>�����TM�u��ޏ����B�~�|�/VP��h�s�&�^��R�"��di�QI(�M=Q�|�� $�+�7�Ol�v���B�~�SV,&�2��=S�Q��D.�貂�:�?�Wmw���=)�6�D����"I�j���T�J@���D
��2�Z�@/���D~����ڧJ�:�|;�B5��7(yZ��u'FI!��-�`���MZ��<��Y����ǩ�3�#)7/���kD;�]JCpO������ =Nr��a��@aUէZ���� E�_��E�]G!�/n�bJ!Y�E�<ν�b�ݪZ��	�_���r������tBj�����v�əM�;�;�1���*��L66����`�`];�'���	�����L̳�6��wܜ���t|���`%mX�8s�uJIoOW����etq�VAg=U7o�v��"�e�ٸe��`oft[��,�<Z�A���}9dĩ�Ζ|��PeLd4���f�w9;-���EӉ~�=MR��& 8�Mg``�g�_"�_��/�HeX��zV��^�?����{�9;�m�W^��W��F��ئ����)�G�����7��juz�XJ*�(J���������h���t�ST�Ⲫ�F�2/�������rRv���{:c6R{�v���f�B��N��c'���������H]Q��KU�	�0�>"n̐����	��Eb3��.th��D���6#�Z�m��w7	��,�٦>!L�}Q�N�/vN�6�EHdO ,�`�Nw���r~�F\�]�B������b@�H6ݮ�D��'//�R�m�����';G�1���{��W�"7S��_BU��<�<	4+r	Cn"�9��O�9߲eY3���K�م-�JZ���������jץ�����3�dI�Z�*t�T��ڨܲ3��6��@SV�_�O�Ug��N,�,�?�+���4�Ǜ/��zjn1��]Yᗮ�٤��NI�j)��	��߶��b�WƓ tɽ�k��7L�wu��:���x��q���IQ4�M��a$gg��yuR[Ո5�[7F�~|�/�p�bne��"~��\������9��k8`�f,c��}�2�M��w��/`J��!60W�ST�8�!��p*7�s�#���mJ�-^�N���{ĳ{/�;�6[�:�q�Fʹ�x�q�Z�<�<���{�[7i�2��ݳ:��0A�(�|=�",�Sz{D͙9IY��̔F�W���_�a�Ҩ�C��H�T���E�w���p�{�*Y����KcŋWA^����8��rj�N[��̀?*����)��r�}�T�9���k���d��U����T�9� 3|a��M�\���`�%�jd ��	6K�%������aφҝ۽�sg��5�Z���f��t�<��Ǒ�8M��d�u�1=^_V��\h��Iy�?����aG����@�#�~���u�Zm��mIv�n��y�w��t��1yī/P�^b��ܲ4Q[�������#��$����l� �0�m��4 �D@�ē�Q�1���Q[�����R8Mu�jSW+&}Lpn]��k�x���}橺u� �M��Ng|3hGP��Ҿ�֍g�1l��ޖ���69\Hd8@0Q��R����xrR����"f0�����	^� �v��`]5���<���9p���n�Wt�og�v����x�	U/33��}����#�@���0s�P*��H�}m���=Ke>�k�e��}qL3&����6�	&��$!Ȩ&&��E-о�D�H�'z&�\UMZ%1�Y����
Ie���.��Z|��z�w�!p���VjɌ{�)G�YG��\��x���:f���j��\�?�1�熃�����<ə?#ں��M�HrUZWҠ�$Y�.c��W�!+B�3�Dd���8�[�����
u�P�m2���6��
�"�+��ֵ�Ț�/E咐]n��T�e�'��9��-�+��s1��Bn[50_�ڰ9��b��BM&-
��큼���<Zy"�78���"fz��+��/�i�ږ��s�1�N���,U}�:V?��a#���70��ű��HB�x �Wޮۺ��ɉ�{���9CU;c/7�AP9��Zc�n/����R���1�`�`�Ǌ,gb�i�aH�i�x\V9�\Ua}��jl��������̲��C'��h	/
МT�u�������n'��[sA��ٓ]ʋ0Y���ҍ����
)��=y(jwEW�P�>�
���fd�D�N��',f'��;M����[�'��\��ж��36L���0�er�>#j��e!��/m�ᴰԓ>2�u}������?���v5i�,��lv;�{{�q�k0�=�3-�d�c����%�>}�:>����Ĵ���l����F�)��{<���Ļ�����&� 3���ܦ�$��*�IJ�=V��_�=Y�����6��h�,����
���SU5���| _XX�Q��e�><�y&?l�8?[�,��Cxv0M���q�Y�a>WE3�u�z�y��R����(	��(7��XS�4L ��`�e
U��z5�й���o"?,�3�0\�)��Ƣ�m�,
5��A�PXj}�}
-��
d쑑��~�]�uU��\"�I�J�WbR�S�.�e@7�����M��)[�e{`57����N\�"\B~�}��$�k�8�BK�������0��4T����{��٭�y����܆N}��ל�s��t����߱7�Z7��$J� "ϳD��j�8���K�k�����a?oƼⶋ�V�~��q��4���ګ�z�@��@�U)#�p)��{��/!��d���^��re>S�����Xj�@�b�Zb���sV`;u<�#I"˹A�ۆ�Z�NЊ�_�Hb��l"�4�&r>��)@x�$WB����u>��E��͠�:��w�תV��j�HG2�yӺÌr���,|�߮sI�6�`��W��==���ek���tj���[H\@F�cERm3�y	91gkE?���'��O =�=}�e	����s*Q���E�� �DF�2R�n�MG#&^1���E'k�m��f�[c�{��i$����VL�z�+C�wH��/�!�Q��Xʹ��0~P�� ����u���;$�}VDk��9}�U]��׊�>3�ɩ�պ
�|�r��}/���@$w����q�:�5�Լ�=�B�8��_[�q]����j�������2!��y"E�)���VG��w�j�����n��O�<��۰�,��U�喬�P�<��s��m��qlm~�����ؠ�O�wPAT�+���r�H�&N�`�r�:�h��N׷ٝyz�%�J�#���r�M��.�q���Z3�2�|�H�uI9�V�^���ַ��w�4܌�{0:v����X�;�&'q� �`i�"�	�m	�Z�XQ˴��������,4���QE�� ��7_����V�E1/�W���)���A=r����N��-`U�Sؐ���D}Љ�I��^ӣZ�sY��������tv�^+��� ;�w��5Ќ*7倪�|��nW���7�JHP�ka�c���}Γ�E�R��ؚ����Е,]fơ���HTW���
PU��O���:|?T�pJ�\��@��Z]pXi�oz���OC���
v17E?�J�O"rC������{£��ڂ�u�IP�w�*��%�mI]�R�����J\�q��#;p�]1@��LÔ�����8c� �C�p��	��V�6�V���a>���$Ɨ��q\1�cX\�Q8v/?���č�o�du���Đ�²녘���܌��n*A�b�
[KEf�>�WI��̒�[q�r׃�pFΉ�bq�g��]�1e]-3
J���:�ҭM}��W�.�Nr�1�{�XO�M$\>��t�r�:����ȞDN��*@���cJ��4���������b�i���/�7�t]�֮�a(�S��z�=U��}��.�n_hp��
)���/kKb�J1�[l!b%� yq�t�ti�2f?P�-v\H -���I�	����D���Z���[<�*r>~5ƤǠ�GUxmE&*�ۢ�e���C��Hww���eKN�c]#L@�&��;m�o&!����JN�T����E��;"4����i�]K7�0.�n�-<��\�q�4��M`�E���өhB������;HP�sU��P�?�}~*ч���o"�H�:e�e~��1��u�Ms[X89�h4�M>34�JM�~�P~	)��͌�6�R���D��h��뗆q�
Ow��̿=H;^/ �j����*��/�M��n�cb�Z b����>�����!�Uƕ�:��*c����s��x���C�]l�� cR&�;�NS�a:�iO�[7[X�Z�C�!�m_a��R��lOth�[�Ie���8��K-� �;��k�Z��� �@³OZ�l���I���[×N��[����g &�k4�Y��=��2rB�.xz^��{+�H���(z�T9�͆L����{��v��6��x�e��U���*�]k{���Lx�3�IEۓ�R��<�w��[��`Ֆ�/��`�|�v������j>f�}���Lo\�&BPA>�v� Lp>�_�C<_�j�˷%�	���yY]����_{"+�*ae�o�xX���Cm���e�ِ�Y��0��M��2ٿ��O����Ӯ���V�^�1�}���g�;ks���!,V?�F{���Ͽ�I��e��Q�'�J���e����!��+4�qQ򏀔x��o�Y�S	<�2K�c~~��aԁ +0Z��`��ͣEh��a�o�STG{a���{�!��y��C�������z��/$*�C~�<̉q�����4�j�֝H��F�Г�������F��5ͨ7|���%Zo���H�&��u��\e�m4L�]���(��$�N�e����8�����r�š��3��Mn^(� ���\��aw/$'��;J���&���4ކ*߯��@Z��vJTEz�͉<�<VA����	X���+.k㣲YK#:�UQ�ߊ�j�Y��g�v��H��c� �,�{�Z�!r��_VuX���6!�~J��5���v���(��Hv�&ֈ2�_s�-N��.e��k������/X�G�o���1�W��Tr��m���q;&�\�Q�Bu�*_:K�
S�؟�TD,�*(໻,��)գ����!|�&�vV�b�0�X��lϠ۬t���y,�TsVn\�ԃ�!���	HN�u
�З�W#�y�)[W�z�w����F=W���x7������y��<~����;�d,D����� � ؓS�3�|�t�ǿ�3��UlZ�H�q�hE��c���>:;���٭0np޽�̈!�ͅzcr��>pg�B֍A�p
�gn9 -m�u�cǳ�0�s6�u��42Q(�i�[ɽN��������.W�;�g�Y��r�B��2X��VC'���f�O���M��� ���������B|�'�d��yrF��(3�埗�C�)�xy^w��"��	���@��-��RьR �*#",�����ij�\许������M���9j۞����R�#�LbUVMk��B�ߜ��־�ۅ����`=��<)�4�IF�G�%�]�F��"�Q@x��t�`��kE��IXc#u&:�d�S�b�R���Vz���6��	����aV ʓ���G�;B'����J�ub�gK_W�����:�79R?��u��Z��~Z.P�z��Sцc=I��3��#�ȣ��@C���hЇ�?�}��>m�œ��lk�o���
������k�h�$c�>�?Xx#S(�2T:I���'����58ڣb�L\�Q",���&�ߣ[Ӗ�O��B>ة��u{�m�~x��v��ܔ�����%._\��G��_���׾�x�YL�vT��.���s��8[Bp�ZD�I<gdb�:e6�{���~�V�7���V1O�Ζ�b�T;5�u�*���Z��sU�s/��ɩdv{6�&�XQR�qD�U�^��v�]l����U+4L)ϳDw��Hz��s�b��;�+.O�=�2�:Q��	�C�yJ2��)��2 ���M��Պ�����B���{]FR�^�p�ʔ[ ��)MxP����Z�r������^n(�g�ޘ�oV9�bo�X����(�x�`%����RZ}ːF���(�/��N̘�:�KQ{e�{������:���Z�䯇��u�^e�?x�����6��њ�g��Pݤ�K���	�Je� �2� ������v�3�5�`�l�Ί�|4غ��:���8�u������$�1���6�3�����Ld�u��u��q����ϟ�,��8��CJF��3��kr�̋������FT7l���kiy��H>�`�i���O������j�g�_iZh{�$�������|�<��<�׃�'�+����H@}*{̣���������b3���2�&����0��?�����Ri�yТ5�B���9��?���D�o�i��yW�%�͍�	�G�e�\�8n'���J��k��Txy+=��Pt���NE`.\�K(lTj*�6�F���`a�a'�������2A����8�������S���ؼpsU�+=`W.�n���v�+��@&������Ω���`*HظBE��~da�97�ҁm[�ș��K�&ua�(A�14L�-��9��]}K�I�7��S�	���m7�&���6N7����@Y��:�D+�}w�*n��.2�Ky	��'�陀VR��5Z����0m�$�gED�E�Y���
��M�FvHoZ1a�*
��u�*���PVC/N=������2�͕���}w��嫻r�����¤�d������Q�/AniL}s��޸3�J"]Igf�'��j�΄p��33�:Y�p|v$T�[8�� ���I
j6�x^t?D�C{�e�"''��̛��=p2O/�o�~�Y�`��K����$66r���5'm�ƕ���ӡ��D@L�}�ILnu��18(v���ɖ�=20Hs��\�����#����4��4D�e3j�FW�~ŏ*f�hoܙeGG�P�ߑ=(���ʾ3�*"ϰ��h��*"�SH�A�[_A�@�2��^.%\�N�^[�"�9k¹�-�������h�m��6T�G�f�*y����E�g��������_�=&d8�)I`K��/ݴU{=n���/`@�ն�[!�� <>o	��h�_���#�3!첁X3��µ_�|,\i�X�ԇ�
����{Ja"���7�J��YӚ"1��ݓ�:���
f�0���T�f�ޘ����D�YVe+���Y�d�H Y;�f�h��Fa��LP���O�jn���h�gs,uXQ�4<V=���D{�d�w4i6C&�=u~gvr���UUMv��7lk[C�i��:2��.-��~\�<����h���M'�T��
�P�=v�T�<nBA��nd<_=-٪�=���7�Ih�W+�tw~�x��	�26����wT)o�a�E7ciD�.ֹ�ԗ�������|��I��'w\x�r15XY�n�[�'���몂)�Be�({h���{D:Cݘq���)�f?Lm.3��P�=�Z>��ֲ����5��]nTXEK�}!v�G
���l�8��a�����E1��B�g�����`��0�����p��+�-�������� ���`=]�̮h�_�����H���΀�ZF �Z�ɖt��ʅ��U~�;�VOj<j�A�#`pT)zр`I������D�n��O)Y6�༸^�C2\�eQ����-���}f2-^r";���� ���}���w}̧��0�qM��J!j͈W"/��9'�w���~o ygDȜT/�C-H��{q1���4G�	˶�`-��A&��_�l�&�^x:�`O@�6�??k[��-`M�\������4�>�[ 7��#J��8�{K�~�E�mkN�e{��з������{`�@�Zl>n�5������>�'�{9-a����ke�[ӁO����V��΀\Vv< �A�X�b�u�h�eDG����v���=�{��0�Ba%�fcNNjL�_��i�#��J:�$�ժGp��L@sD�`S�`Ec^թsK��v��B�"?YѦ2q-r�@,��3�C�����>��	��-�z'�@�p�ֈ�U9x����u<��B����%f|=�է%����V�]������l>����:��<��Bj��&{�+H.٧����I�7#0��.�Qՠ�q�W�]J���Wš����!qa�%����_Ȇ�.q�t������-i��+��F$��ٖ�mH�N��ꪛ!54Gн���+��7]��X��ȒC>w������d�\�pu�5[C=�&Q�O��ߔ�	�vj� ��v�5�;k���z�P�r����&�U��B��`�^���n�����7w#콇T���%�EA���Z���k$SA�x<���5L~s��*�=:�t��1���В�fBo4�O�9��f�����&��W���i���%���1�0-�����Yx�yդ2�w�w%!��v0�F[*f��Vf	B��a:�Ϛ��Uˍ�)�v=*몜���ᙬ�9Ĝ��~i�7n�	=�+R_�%[��3�k�2�(u&�V�r{%�\��ךl�ʗJĪԙ�O�3����:�fw6Q��Vn�����aĢ��|��;�F�,�	�E��=�;��������
fX~:d�/��[ �I/a}�,���TF��a_��Aڇ��Q!o9��]�l��Αޜ��0��^�F���?r)��st5_�<c��>2΀��L�b5�x��ƀ�ʐ*3�pOj]���.m�o5����C��׸�Kn��\M�,a���D.�?µ*e��a'��2]�
�F��vZ�p{���n3�8S��Z-�I�k���o�Ļ;J�;��$�V!�e&sW�;�Q�i��υ�/#*S�[�#$K�O�S����r�i=>T��LyE����k�ydB�ա�t�	��Vl��O|y�b��蚩�j��� �O�.���X��{m�@��x����*��o�?�ۅP�N�a�W�>.p��l��#LX�%&�#�u��'�L�չ#G�5�(D�̖\���1�5��i�g,�R5� �s����	oi�Cg!'�ب��h_�9�S�e]`JN�m�^�ǥ.��3�&�����Rc�a������������ǿ0��6%\�!�2�Lў#��i���{��ƆOt>C��_Έ�Efi�R�W{�4c6���m$)� :l+�o��5��lu����a�b�K ��ז[�|R#Mpj�L�ϼm�j~���'��P����wo�ڶ>��:䅍U���̈����X҆�v���G�%E8F��3݄��\�2'l���g��^$�-�7�)�5f�T����!$���6Ntb�!ɍX�`�Iq%�S$`�;�v_:�[�T�d��R.}�-��j�V��� ^���8]QP>���r��ʧ������ �"��wbؕ�r�[s��U�S-��w��#�}�]L��h�'k;,�����3��Nە&K�ф�x�f�}9V��(��� �n?��t�s۰��N?G��3W�6�펾��a^/�h��(� )����5s�����`����;�%�aod���0����W�y�ì�x-_��\P�f��X�g=�͗wB9��i��>���q���qW�ޥ�����\��'�ǀ��_�T$m7��j�(���n�[ߢg����L>��A$Zf��-Ny{9������#�YT68̮�p�.�5�r.5���`��� �f�H�p=d�B%(�Z�}�9��ese�_S�*�j�x�Ju��"�9�_�c�6��]�=m�SP �����z�5ar=]�6�VP�C��8&�i�>��v�y�Ŵ�lN�>�U�kK�}B9���a�����!�:)����_ �ծ���*ת�>F�ߒ`t/�'HW���ٟ�h3#T�R N��~���$+=n�N�Oٕ}�k�
�M���� �$N/V���]XGq�6�G�$j�� �m����4�r�x��Yc~�Em�����[<2���<����L.s�/�:Ix�=O���-G���e��0�+����?߇�(/%��U�H:M�`�^�W�j�v܆�$o.�k)���2���-�)lC�z�hy�G�P�㭉�8|��c�%��4H5�Մ��-2�s)����,�í��	k���������0>.�wpU�~MH��}�n�?�H���䙷T,��q��yCE<�qZ~��T�l�Xw���Q��]�Ks��=�GfƉv���=t#�� ���2���j*LN��5��4|��q�5(̅���8 ��ξ��늛������?�:Q@�>z4-��q�>:N7Ψ�d�8�}�����n�D��njpqy��l
A�����P�C	��V�t�"w������e����B-o��%�2%I �����%$�H|�΅��VL�"/!$��2K=E������-��'Y�c'Ԙ����n�9�)r]b����N@�L�^h��t��v߼Oǲ��I��np��Ϋ"�u���$��tG�*�2X=�D��&��D����"���B
i}Δ
4��WU?�k�6�q�_{�{��J�9��L����`�i8q���	b,Dѝ-���gc��.�k����N���A������.�5;1�XT����T����ZÐ}c�2BdJ<I��9�N���bs�MF-��8��7��R�h����7l���ZyN@�f�T`Q)�U��D౨��t�/R]4V~�TD�?g����G�&��W���N���
�xٲ9�bi˛���!J���/���v�)p��<�N���y�e�C�9��&�c�G��)��e��4f�����y�W�l�>���[	�;z�9�9i�HV��t׫qG-*����N�X���_@B�%@r>��t��yID��#̹�{� D�6Ml[0�A��؄�q��0����,��*�s-��,!�RQ]���K#,M*��c��=;�J�g��5��I�ѰxiC�x���z!zh��_��歏����F�g!
�V��O�Ŝi"ڂ�⺔ʗR2��$҈�ЊN��Dd{
�iS�e�M����WZ� �'��?���D)K QGzm/�&�<=�j�#~A��O�U4�X�5��h�{���
�^ȷ�L㌂r�Ml��g��޷�nx��8Uh���Fˢ�
�����o�\F�E�(�e j�ۋ5��f��S��/k��7���M0��7:���(���r���s	����e��9�u?�Sc�C�)5��?��7֣�>��Uj���qo��]$�c�V��v~5x��W�����%%�d{g�?;����8�w':���Y��j�ܚ��y@CK� ����T���� WW&�/�J$G��7��-#�m�����Z�2_���=��eC%o�t%_B�믔�bcB�4�C��92S-�����U%5����+?ƜdM���}R{"��ں�l��������$�("�Q^���l���5Q�wze<�<��0˙�!��N)��E�W���HP98�$Bβ'�.乞4`�Z�R�Y�"�(��U,����
ꘀ�=��K=J���&���e֤W��X��!0�J,��i���}��p|�>e&��V�J ��"�����I�)i֑cB�];)!#71UϺ9'���ư������1m#�W�^O١r�z% ?W.��:ΰȉ>e�.(��S���_}����+u���J���\[*��	ͣ)[���ƈmQ�G��/����֕J�ӈc��ǴHR���Q	��t���p���1���vi�Y�ȡ��Y70��g���y"	C�5�C���iG�X�A���s~l�z5�ZqL�qq4�D{� �Ja����sI����s���
�X��bۿН�S|�wNޜ�Ək���`�Q�,��0q.W�II���P3�F5�6��B*~֠�A�b���t�=jq9��	?��S`i�7]��,�
T�?��0w�L���f��{��:��'[��[D1EEk��s��|*y�;����럷�/R}���}L��&�¥)R��_S�����,���lj�Q Zf��+���IJ@�!���8z�Q�>��/�3�ɐ��T���UY/��kF=�˫}ڵ.�>Rɋ�ޚ����3+[�ξ�q��D[�>X��/��7�%ov)�t;<�i��*ϵ6_��uc�s�X����$K�z�s��/S+y_�I§��S!�[$�lS}�D`�o��+���"`]"+��BB��k��ȑ"�i����{'~Y~���X���2�ɠ�W��v٨�&?۱{�w��f�E�.�${s��>�<E��d� I&����!yv���3?�cq��VD�������r�ۃR.����֋aO�rz�L�E��lPi[�����R����=�#��U�]�w{C��{>˙�+E=V�FP�_l"ϐ�Չ�<@-�~yY��"#��#�h���F�^'��\9b�f��0�2K�G6+��O��'H�%w�<~|�H�&������C_\���9_�tS�]�QO�o�[^H�^�� X4@ESݘ���H0�I6G�ד�Hz/�F�d��s6��nH!*���¸Re��A���Y�_�c�`Vv��жG
���X����7��:D^y����������f�,|	�s �#�����Vϫ.�9��(�.�\�G��z�#y���4��X�� ����2`�Jɭ�E�"ة�	�b����`�Z�X����L_���������U�5�+� ,~0����!M(��ɮ�*3̾6�b������E�Jl�	`{9��y|k�4��2��]4"gF)��c���aEc��\�)�D���<0�� �Ž��^oJ
�_!�dH Ƽ�gVB��s�Y�B�0����J�}��,Lt�l����������}e�@ZόԐ��9��#m���첬�1��� >� |��B�JJ K�4!�_^/IEB�T�����}Gp���WM���z��u��M��~1��%+��N֮�$���W��r�;��3I�[M��{tWk�A��;�KPv�m��%Z���P��*���ⷚ;��ʋB&h����	E�ZP�1|�<>a�Y��xR�P��F-50���$Ȍ�_^�1��U:m�O��`�Rr��R�\��0���O"�2�L��4�]���a��w�����ChS��JK�kP�.��qw�^"����;}r����7EU)s��K#���Y��x.m���ZJ� B�E7j�keX�ߋ[٧Ѿ���,0(���d�@���G�8&:byy����ubE�4`���aü�L�v�_3o�s^EU�y��5E.ޕ oE�#�� i����jf�.D�}
E�MB �v*g�Ϋ�����i��_��W�ʬ��:�v��Y���hZ[�o8�@�ɨ������y/_�H�ނ�����r�Ȳ�&�V#[�W��_�ב�4J��Z���C
:z��#<Ƒ����t�"�7D<H�V3s���ʃC�)Ĝ�ی��B��3���E� �:��:�Ym�ׄ7;5���˯5��r�_��$���π�:{�=^E��h���N�� �S�l�:j�jU'gs��m��ԑ��I��s���9��\�O�4�#�����j��I��,�q_�C{�x-�5���n.���ͱqÀ?.�s���=�N�P� J��������C1��?if��S�;4e}��B�4����;i�8��&��Ɣ����t/3���!���1�"J�x5�k�9�m��k�$C#66��2M�%:N|saZ5�����W��&Nu"*S�2����wT��s8窶,����v�V��v���C��(S������U�X~/}\F��/�	Y���N�b�~uf��XKJ�-1�[�+2&��@:{0���Z��@���w`�Iˑ|J%a�ס�֪p�7�6�毬����W�ؽ���8�Q\�\�ㅳ��=cAwH)bs2��k]���:%��~�-}`>#��8N�}��
8�͑Df�!��
ZG��eOFRy��⛽���ȌHm�X�2�_��;G�h��r�jZ�:�G{C�,!���K�x��r��`9�^V�=�{�$h(��Њ��n,`������?�'�
 Ц�S�k��`̘1�����?�#��hVۻ���c>�3�k��)�9N�W⩧w���'�f�!�����8�u�p$n��W���9աW���#�����h��\g��N�f�j�Z���̼�&g�+(֐�2��K["��$� D�$��G�" ��;>�SL�|�G�Ւ&<3�*1�d푷>��92�熠�2sX��ϼap����6�H̞g��)��	��g�w���n�M"�g ۊ�0pz�>�����+Y�(�v�EYؓ!27�D��/�$,!���/��@��@��5(Jr��0N�d�����<��	���f��3��Ó
EX�ӹv�nVD�@�	f�OJ?������ ���v��yZ���	�b��#�8��ӫ8��nl�l��T$�O��{��ߟb�Ȍ%�2s�:���] m'c�$���V�2�3�2bLn�c��v(�qR�Q�w��#h q?L�R�G��&�E��C{����S��0����[E`%���Q��2%u�>���x��ě�s*JL{�BF�/M����%�z��2��@:o���}���rS�".h=�$��e�w�@�#A�:���ƂK�~2��f�N0��^�)T#�~Jo��F�Q��O��d���S����O�d�/��?Nɥ��x���,�Ȏ^m�y�k��t�;�*4�û�/��'�'7�՚A��x�ЭMy�X�2�!S�{P�O.�6������>�$Cc��U.2��:���ʌ�x&�˃)�]��h�@D���m��vz'���B��յ_�E��q6l$HE��84T�o���eY	(�*��bSك��:l�����2{�Ѽ-�;�_������:�F����r�__J
3#N<�MZ���9;�M����=���=[��[\��3y�l��>;Tl�gX\3`WUػ�Θ0�#$���/�r�6ںX� �c����nK�q���ݻ˸=�ΐL�w����A��E��9i8�~����Pøs��R��O��^����˦�'�X��v��Q�z{~��?6�T�!�~�����|�H'�.<&q��u|��,�^��|���2M5'��+��o}fM�|��\ޠ��]v�@c�0�ߑ�ʈ��׵Ė/�4�rp���Bb�@�����"��vk��_̖9�r.�ʪ2�}wߕH�[�yz#����6`aJ@r��A=����q�~�/-rp��+�OSc1_J��uk-k���@xc�ϙ��U���ϙ�v�2R>x��Z����Zж��R��W�B��Դ����o}җ�Ŀ�5��f+_�����m�_T�A��K.6�H����dW�a<<��<B�7�q����R��6\O���,a��O�@�f�ϊ����	j��q%�\�k勡|䵘2��%����)�o�|I���l�G�E?4s��j� 2d��u�A~�9Z���Bm�Eޮ�a�˓Kn�`�X����Q�)2ܰ	rp	���e(ˋ�}�H��KJlQ��a������� U=	2��%{�Zߛ�^ޝ^�K���*I����a%��A��u�s�	j�2�"�J�!%1�_�8����/�k�!et\�M�VZ�\d8Q��U3�X�I�dk��u3t�>��G���Qua��e��&߮d�{(_h��m���f�(-��z�塨���s�+Ցm�ӿ��%1C�G/�o績7��p�����R��r$��?��@�S#�XPL����M�|2����OA�׾ke�/ƃ0I�K%�.�:t��5ܿ ����9ͽ,��p?���AU(�BMpt�cG���5(t�Ah���7{�A���|�
�ӿ�f^L8R󻭒8*7�W�,�c����	4��?o�ץ!N�!���o�9k�B�c��]g�!�~<���9Z�sH\"�GV!�����0�`&����"��q��=��bG��	U�i�����NX�?��Wv���r�Ry���t�I�78C�걵�O�@�2�q1�,��W��_`as������-��W}㧋h�t��쏌�	r�"w�W3P��:F,8�����Y�����DRsL�����`&?V��2���f����!�
��ebNwI��᠙C��ܟ+�#�P u�+O[K3��pF�	5-�p��$�D+�ݞ����]@j�/�� ��fR���k>�\�1�q����._^�q2�ܜ�
�:_a��v�K.����`�IqY͖�?%vВ���D(�I�����9���ѡ�J4㖗��z��f��wN�C����2��Yo�S;D�$�$���	��VW7:S-( 8�':Z�% ����c�:g��S:�ӚBw�{�R`�����j�d+���d�bN�L����AJ�TS؟4H�&��Y`3
5���Ӿ<D*�6~ �{4����=��������+������^�P�������OY=o�&Z,#�i�>�ڄFB���A�SL"�Y�i9I��e���y�%���+���&*�e��5P��o��f^\�v)�X��J���B\���	�I� V [P��N���ǣ�7�2!��d0%�������d6�(�B��x�{0�+���%
�-����[��g�ʵF����w1�ɷ) 9���lD�a����&ӫ`��4|� GY16\���e�zlS��.���� �hI~��sу�ڭ�8�D �"���X#�v�E��M%9�.&�f����V�_�B�����F<�HE>Q�Gl ��Yse�Y�$��z�"��29WV��JLQ�UT���5���VK�����S��K�V���`���q��	=6��A+�&���؄ �cfM~2��}�hm�M��R�!��x����
3�W��v�6�##P���E�����d ����aPϨ
AR\ �u�8�����=ZK2s��e	Ng|�)(0�i�=B�Ӌb�n���Q��A�������\�N�1��T$'�86�����%U�����F���A��'�%&�,ԌR�ھ��plC+=(723�I��2�r��O�CI�Q�f��s�����4��V����As�~��L9U	���7D!T�uA��2t����!N�h���t�삔�*�����%&�>�P��8�:u�<^s�����.��6W��	�n�%zC�s"�t��mjS�?@��sZ�� j�4~y;t^:
��uw�����-���S'qZ8k�H��V0j)��k���I��,T��a����UQ���􃀑̮��z���S%�8��S�gp��xL�-L�'�	�Y&>�4��K	�c�����Td���.�5��+sD���YN��)�1_O;��`�G����e�Q(nw88�-6,��v��^���Y����D�i�.KsV���.��Ew)�F�޳W����v��U�9��0?��>��'p����	b�����w�Kj���L������{	���� o:�@e/o�8���0L�sZ�P��Ԋ���?���ý=����4D�=�XoyjZfW;�3�;������놑؛��
06����1���Y�Һ*n���	�N��8��r��i�5/�����Cp��˳5��"U��XϜBN
?�-!��Ջ�p{>��ijx�)>>�Z x�u��G�c<6��E�!Dz��mx{\iz6�P�A����̅X�ԇ�S���Kn~��N�0�������=�f������I]���1-UM�晪+_�p}ɗRC��*�p�J+��0��#�bkx�%�=�G�W���^u�yq3]Tq���G2��O�	1�Ǩk�u��e���ϱL���Ԡ�Y�(Ӯ^ÅH@���8�t�]�_����ʸ� F�uh8c�zÒ�±L�+Jg���'�)*���tY���3wO�^�ո������EA��T�	$�Ӑw�xn���|��[���'�~�e��o�Soqi�P�_[8=z甸Յ��x�}��d!Nk��N����NKb���ށm��	����j�h������f���T6���q���`W;.�6�c��fR�궵��ѓ��7��izc��תf>��lx��⍽`;	&��2���^a��@��$�}��h��,L�=kP_@���V��a�Ȏ7D�k��y�Dw���?1�0}�G^<�����A�	�<:b�_5����3[G�#�NB��AC*�b�6��b��H~qV����p�����?��s� ���>��s�lzH �M- �S�(�vU�:n&G���Xq����=���� �{��v19|w���51w|���@J�7N��_��v椠�s���Lx�@�[����tz�Jk�@X�����������Nv~��~����s�#mt<8�[�_�dD�R�NC��>�8A��ĳ��k�\��W�-]���x���g8���&bP��H����-a��ʧ�]���s�g>����P7_mD�Zo1����@�c�fD���ºC �5�а8���yK7c mg����m�[�>(�e�V)�:�7z�R�B��a��U1I����S��U���j�b@�w:�JF�sH��<�1��%x��5��q�8Ie��Ѐ�`d�A��d*��p߲��T�3z���4]���r�c��	;Pi��$�pnf�N{���`�=,������V{\�l���F��1�q��b���2�_Ae���l�"OnU�"]�'�����>�@_N�:<��=<�}�D
�E��驸�1�UɭD�mB:3t��b��#�[�:�O��c�c
�ʘ��R�Ճ#m�4�|(�]�Sᴒ
��FzoO���B��mWX�/&O�|�F+��0an�t:G{�̣T}�A�UdY��YG ���:;$���}K�Ce8s����ݰ�����M�3~=�V�e$��[`�u���*
���&�
�JC��g|�夼��OZ{]�-�ƹ4>c���C�-:���];U6
�5ɜ���l�-l|%��΃<��ގKΥ ���a[f@~7L���l����Oh�Z@��W��;я̡������-������B���������e�k,>r�DkH�(�����0�+���3�+Lж���d&�D8m����7��rbP��Zߟ���V��Ͻ�wɑU�-���67�{|�Y�棬8z�I~X�>'����|��hHCv1��Ă��"���`�����,XFlB��su�e���@��Tq9bfk~dտi�Fd�Ժץ���]-�ѤBH�K�ڵL�\:Y��Sw0q�vn �q�n���o��.	�O���Rh��B��%:��(�F�;�pVRq[��pB���Oj�P����&'N�]�ji�:V9�Ϸ\���Fg�U�ӠZ�(�WLƾm�����5�U�<_�<��Qι�R>Y\co�#���fr��b���qr�����
��\Q5�}���X(a�����������
h�y�.eo�Y��c@���e\T�e�]��m�j����Ո��O"fJ5ŵ����ҷcM�Q�+�q7�]��ܚS�Z��������)'㿲G�
vEti��rD/'%��
��IN��v�2Pk�_���N3�@{
Ŝ�~���� ��ƞ������V��I��չ�`=�A���@dGΤ{�em@��b��@���XCye�S�̘���ޟڶC���#4�0Xd�kg�{ r��N���A����:- ��y�P��h�������r�i�Y����G�!��&jK�S���z�7g�]Ow���4�K_�w���,�<��m��'����M�)\Q����*�sJ�9���]�ጭ&'B D��Q?��4S`�$^�x�f �i�����c��zX����b;�Al.�O9�(�0�9�b����j��jQ�}��܇1e�Ow,4�����1��+��I4����DiK���9�+�{j��6�! )��w��s��D�`���>�,cQX�K�1 z�j�.�;��M\mx� �7b�泼�hgUڣ�y�(:���oj�a�P�V��	���rV4�&l�K��֛�`�i���z��k��w!�oňT�מSd{_��B�Գ8x����9}��-j��vO�ǆ\��ٛ�J� *Z �LB��?���i�٧)$V>#�D%'�ZV^�~�{��e��d#�M>�er�R���Y�,a��eE6ҏI���������d�󇉗	+�Db��7��R��Bf�)�w�N~��L���8�o�HQ�;���CA_��(~�3��LUg��O*�����$��ˋ�F3n�k4�N�v������p��D�P�����ͯ\\ޑ���vƶYLY�����.x�S��(�*!���6sj������ �8����� }7�����?[ɿ�X�#��(�Op ,�jwRʾK�Ոj6��/
5ou��?�`y!�O;�B��N��`��'8���?`��aa�+&e��������=�ɔ
<�z;��R�8^�T�V ��D�`�dl�2`��3�'0ď>�z\M��,޴�ˎ�:��2O�o6�� _a>��I��:�)�.�_�u9�ْ-ˑ�|-���Ȩ#pqD�s������uo��*L�#����r�K���F
�9�I�}TV�}b�����;Ѭ5�0a�j������o�ՙV����[et�7��R�����P6���Qa��"F2~��8��L	���U6#�%Q8l$��	]�/�P���S�G�R!��Ʋ�DO�I���܈Tօ�Y�MJ��>�HJ�֑Q��! �Z��� ���B��!�aK�XG˰���o�Й2�ȃ��d��v5��-�����`�`V�8D^���.E.�#��z�h˟�+V$��5f�p�~����g���J2cHF�Ҥ*c�Xӱ�.�!�B���Kӵ��^e�1Vlmo`F#�����݁E�ʗ��ߨ���=����D�5�ý�Ef�.�&~��A �(af�)�Ձ=�	��}�wّ�>�uvs�.��!��lm,�`⾧��#wŶ7��n���j�}�_�۠@Iq��Oнf����!�1�X�>ڎ�;�REΗ���n$� k:�ۨ��@�+��Ps�F��k��W3���(!�R�_����>1�i���Z<��
��vqBꖎRŢW���{p�?�C��2��Ggy]�i�`�-W2�ۤ$	�@��$���ʡL>���*4C�c�Ћ�F�^�Y���Btc4	'�`fp ^m�����j^N�ȼ��a�
�@�l�C�	4ܮ�P9�)�#k�Em��f�B�S�~�sl��5c�1��t�72�n\�Ѐ^����'�p'�vr$��2�|E���	��$R�Eu�.���2��VN&ra�w�[��D�lS"�� ��h�+}�o?�v�<���*�V5�f�ꢍDj�K���d^2I�M$�UdKK1��=}��7G�j����~�Q	%r
�Y4��tQ���"���$�w��4ٻ��D1֑����D�p=bd?��ʒe�a�w�a��W*T����Ǽ�GT���gZ����)n���û�>�
qc��#��HBL����mJ.͵�'~`����u�mR���*�2j]�p�R��Y�X���@��!�?<�f�"�z�,-4e��z��̘��$א��.�����3�ߢ�v���L,�����UW
J���؀R��9/(�9	)��tT���k��F}�c"�<A�<�V���>�	�I�kn��ޞ}����c����8G!cΦΔ�E�2��H����]b��/�{�z��#��,�������g�coBY��T����w�G�:9>�=��m!G���ƱM'G�/�J�H=` ��D���cB͡.�
���g5��e���#�V��y��R��;x_��cs��z���x�@�s��g�U���)�L��~�����4=��A�{ka$P��B�y��N'_��������VQΨ�$s�F7�%)Y�b�/cp�3UQ��O�� j˭wM��G��X0$�����=>e=dN���u![�i|�6��책�g�4WG�� �Q��z���w���a�W�ƞ[��n��~���Ql? �30���{Yϔ#@;����r�Hsڣ��֍���z�WEh��6���F�Ŗ������ȒH.YA���c�+�V�yB�ZR����&���������*�;����$������c�����s.��F���kn"@��Lq
��f���@nR��6��J]וsS@yl�ʄ{x�Gq��u��ձ�Er���(O��c̪aZN
�����EEV&h z~��z�1���]^�;[L:cc)�"p��P����i��}�NS�Qg�����[W/6�E�r[H�8Kx�� D�������xT������)���3�9�M�5u��;a¹	sWY��iݙ���PM7�6efZk�*�Y����	������v��`��b�o�exܲqr>S<O�?�RPF��6q�ȁ��(�ϯ��B��[C���#o;�e��=�0�
=�JE�,ng�VS���!���'���H�'Q�e
�yme�z�f ��z�ԫ���)�G�xEj7�]+���wbx�;�oR*ˏO�jq��wz����˝��(�D;}�:W��8�F;����ҳ��~*-;���l"�jB{��)���^W�ٌț�#cx��6��7Q��ۇ�%�`��I�%��6%�<\���{Z&���)@<}E��ݷ�>I�{��#�@�<���"��R^�����Y���j�@�&﵍��J���k�za��*v=��.�2���j�m�='֜�|�ƾk��k�-V<�0Vm�չɹ��I����	�D�E7�T�bL@�D�z�,�u�>��{Dn~f�4�O���x���TCA���i= ^���\	� �45�ہ���w���EBӜ2;�FA"�w���*�6����` }L���B�Ս�"Cб���C��!��1g�.5Z�P0$����xO~�[�\��s��{h�Y/��p�j�1o�@����;��18�4�m[y������"
w^�8�<�d�ir�܈�t�5�f��rdr�uHǸ�]?5uEs��H'��!�n�īA�[��T�L,����3��;�4��Y��݃%�=e�r,�����:hI�盼q�n�|rKiXv��d��$���pmM��^J@��;���ޫ��Ţ-)�4�Sf�#9ۖ����*R4����p��8��Q Z~�9�yK����9l�ۚE���;P��ttt���ofKh⣡�G"G��h�G��x�h 2�J�(CNH�Ԗ>|�+�L�Ӛ�����+m8p��`�D.^�*����=�&���9~�*G�VX-B`\Ȣ��!Tt\˭�j��AZ*jƩ�r��>�S�,�Ly�Df���>�g��@V�_��e�-8A�$3�";ה�!�����:��8t� X�Y=v����4=H��-�U�{���o�ژ�C��|g�]ތLca�m���jbi�;�X�cѢJR��aYY��r���8���Y�f.��]��O�Bs|��3�4��6�V�?'&ݏk�'��vT0d��k�圗�UC��o��N_�(P\�ר���[^V �
4��'�� ����%0/�W��jU��]���W*I��i�B�#-�چ+�8��<�蓒��#W'�K:]�<j�D�hfH5Q��S`��a��K{���Rg���w+�9Wb����r��t4��"L���.���(s��E��9�l*�8�#��|QD��O�u�U��~r�Q4}��`��s<<w��` ��o���	�F�$�@����5�P���!�S*�{�R��7M�C��#�h���+^[Zg�F�`�+�>���N*h��{'T�e���L�w�/s@@Sl�N2&WP���!���FI5{P�/�����?����^�	vh-�s�0C×r2`�핚��^B?ƹ+2v��~v����e�/�-���(j�6��y�ZF|ƿ������ƾ/Gف!�i]�09u��I5��[�v���3B�ф>F�����#�*_b�;T{��]C�������Ea����V�G죁�}��?b��B�����\#c����T����Ps鰙5U�al�e�s�p�� ���%�$v�G�;�%�k��l\��<� y
dd+�ʇL�cn5 `�����#��Ic�ycZF���C$�+Y���'��=��֦7�1�?	�aK���P�ь�O5-U���Op q���)K�v3F�7����waMi�����7�����p��b�Yi��}�v��>s���<�#EY���O�Ԑan?�9g��o�j]�yK���T�\�����¡��U�~Ò+M&T��`!�֋*�(�0�nbS�c�hS�"^��Y���󌸰����L��!�4��@d�b+6�ۛ���R}W���^e�D$0�׀�{A�a"=����ˠ}�����H&�n���y�)=��N����<�u��1=��2ޡ[�+8>F�R���̄��ձȮY�[˓��N?����B��Nm������6�凃L��n�1�_Wb����������ֈ��"���&���p�sr�-V�S3
bV*��$-�2u���n?�I�Y0`woS��%ؚ�;\IEFV����[ȳ�m҃�'�:�,���sȫ��չ��r1����/q���ā��|�h��׆�hZz��&`_�ᄎ�F�����4�L?�Ѓ�Z�)��{=��H��-W��!���|�r�^}�f��j�*�m��( ���3�oZ�f�Y5s��3Hj*p04u=An��������8Q�B�̽��qY٧���\�9�>X@� �.@r [/�8EE�G^�NY���N����*߰���MfH ���4Hq��k���=M�F'3�i��F�"@|�TW�p�8���C��B&�fD=�?Q�K��f���Z�ý+W�0�R��7)�q��%g�$�^8E��r� 	�.��+�����9(��4��Ű�ԍb?L�EJ�����k^�Szt*�V��LP��cQ.��쓖Mߛj�{�q�~�)}q����S���]/!����))��7ot�玘�ɭ��a��\���d�a�v�>�bp�xF�vv�b��͛��38�mP��s�ؓK���)��k��f]���J Ѕ��1��4����?�v8��4H'��mqP��T��vw}�������n����dˣ���G,a���oV��xY�z������i2�l�����i�&�&+.��v@<$�o]��+p��+�Cc#������C�쬼*UY5	�1�x�6C�l	 <ׄ&���e��Hx�_�b�4xӃF�e:�ޗL��&9=t�~���_"D�"���et���0*�zy� �ޠFe��{QcC}q�����S0έv�rI�q��.Q�08A��c��a�M��qs���07��:�\MS0-U���OYb�����=f�va���G�zI]ΖAZ�gU��u��V��.@�k�	h:�L���{����C���Z^�l!KB
�6��}DDM �%�ΑU�z�4�[�J|�&qi�3�Zp>:��U��D7���KY�X�Β�=_�Oe����>�F��`}Gg7������Sf]�]�����b��B̿�x��aW��F7E��#bB��vC.ߘ �l���9�^]W����S��g��c.�cZ3<jTK]�>�씾��]^��?���n��?��hǵ�_��/+j9F�Z&��X/�g3��m����~��S7V��a	���85K�=ͦ3��o����D�He+J���n1�q^�F�&1�Uv����qㅻ�:v5uz�K��Z�آ�&���%�^�`�Si?V��3�_�+��̃w_�Y�B��ż.b ��+h.�b��i6��EKl3�*'��)ܴ�h�	�r��@�֜Ǐ�y��F��p(m�.N�3y�yUE��n�`zi��s0fzb�E/D&�1�+;X"�^�к��Y�l��~����ե���(4�/���_j�J���g7#��M�d�^@a��
l�D#�z5��d���&��I�'�:N��q���Н��\y�@�o����5Xƒ0����9�xG)��e+C>�DV1���ճ�>D��:J����dK�*jՏ(� �˖%_k(���M�t��)���U��/	�$H� ڄ�LrA��D�d}Jjr��[��?�oxf�ي�-!�_���T��v���|�ڬ��5�6��j�)X�'"x�⎿��v�Ĕ�A�C�>���y�$T�ğ�p����k� �/ϬF,~d��فU��d"��F���e�����~Z�+jJ%-�n
���,Mm�����?p1'�P
m�`姴ωk���T��-��m��y[u8��Łb�QY�y��*���:��<s�y\.��V&p�-�:��h��E-Ju����Aޛ$��ѼO��_G}<x�B.We����2�g��("*�h>t ��e�!9Z� _�]��ko/�ͫ�A��]->b������#�Y����n�����G ����~�=�p��\Q?�Z�^���J*��e�H!�v���R�y6�L(�ﾠ��'�ܴ��aV�I2k�vɤ�g���Äԣf�$�O9`���m��k�a����NyG��	�o<�r-�%�� 
x}3�c�H��-�OF��W�R]�XJs#�'�2k|oY>^��=�.]����:Ӵ�Ge���fS�ޜde�ah������+�����
��l��a<���E#� GH��	��q���D����S*g�S@�2aT� (q{v��P�������}�܊����ϯk��N [�C+9/�@��F�?X�r�����C�@a�("=����c�';�((*�O�P��.р��l�� �nԃ��pwf]���*����Eg�M��� @s������Ь�
���Efp���B�����ͭt�Qv�[�PW1F2�☇GکL��*�/�g�7�6�_ ����I��a�)�6�4}�}=)S�����G�OpZd���Q&tK�ꪷ��T�����~�p� |u�q/�<�r��֜�Q���������W���VC�	u���7�Ѭg�***M���j���3���$�w4�E�ڄ��ZHוX�f�Y�S���蕷��ͩ�G��Vvk��~J�N���� `j�)U��[��|>.�.o�kG����3�p�޽��໠�8x�@���P��t���X�r[HhƷ���]lb�2#��c�Ū��\�~�ϛ!�q >\j�59��Ӷ��'pd��0PI�ƍ_,��pj����r6y�Z� ���؞@����ͥ�s@ ��)]��� S��q�BqV�&[���'i�7U�`���Hcm�΍�j��ޡ��"hۓ���W��>B�ܐ�P,�M�P�ǉ�ߓ56���@v�{�J��/����q|�&n�
���+�[H�oi�M(����a*[̩�p�m��(�����Z��`C�=�.h�^@���k��y��w�;�dc��<���W��;��K�RT+�L-q���쪽�r�^0:�0"}��].����V��"�6�=�A��WC�x�a���Z���Z� �g­�}{7�?�7.��N>	��]�,��MjU�)݇�ce2���\��\�~�Gn��E��P+��7��G�7
�FɋS3ud�\rDm�i� 昔����߁ڤG�
&�!����o�g<<��ZB�a�P�):,Gv���;lw̑`�c�P��oFУ�[=
���V�±�+�
 �O��3��)�XA����8��;l��ԏ#�M}(��I�$8\E0�G&���'������	E�-���pkk���fC�<_s��H�$Yz8/��̹�^�s��T���Xl�� ��������q��!���.H?��%�W��f/#�im�y�Hn3Y��3lM4!��ڐ�h�z�bo����&����l�q{G����^�HV�dq���^�s�08f��Ļ�͑V������1�H���2�7��K�nei�1�]1)F��"����њ��#	�ɂ\&����<+A!���0ό�$A(�ټ������%�0�v�";�aȯbXq��^<Q�����<v<�СOZ����y?���t�C��Z�L)���A��������%�I�^AB����6�n�t+�n.I�-��A��[['*Z�r"�a\E%���{<�^�`-B ��$��EG���A�[�IK�l��Nʶ�<D Mׂ���T->��ӻ��ۣ�+g�%˅�$Ԉ���+t�k�l�ō��񕮈�g��/:C:@��,q���鍫����/��k o���mj��GR�ט�ރ���|��Uy�"2�}�W&�W�_�Oz�Э
�͎��������!�z�Ô�ci*�7��cѸ�)َK��#Ėo��`첊}�Ɂ���C��������>�4 ʡ{�2
EL\c�Y�x���C���Q�"O�p�^%Gw�R갰E�ht�s��7�����x6q\Q@���""DG�����J�p:ˀp�{� tK��5M�0�y����A���@�>�|lDd�e���_�3������FK�&�NПZ��j�8���t�M�~���a@y��~��o� �y@(�kl�f��ƣ�ysb�����:f��&Rgb�-�]�� Q�`4�No��_�%���td�������*�	�R�,�9NG��#�8���U��ş]�Xk0�l5������HU6����ȕ�TiRy�Њ�K'��J0����v�_�[?�{t#�Q$c����[۲�?Ӵ�U�4rǕ�R��}���xi��3J�z�pwW�R�W�ZZ]�P"O0Ю@�v�Q��}$k:�
0 X(g�4��o���v���p�FD��wL>��GD⅂��C�t�$��u*��߷����Z�V��[`�B+V��{�}�މz�aT�R�j>S�����y3�A3�ac��g���vgT�Oš�=N�AV�cA��(
�a4�Q~pA��� k����,E����U�Ҙ�A�O �*�g�-�UϬ��>�<����Q�geJ�@_��ۉ
Z���g"�Wnዏ�OEd�ݘ�v�ƺ{���������'4�#Pa�ͪYI��Yc^Dʤ��{C.`��wFim�<�;�����DS�u'�c&�_���;�^��d;\��i�n"���+*����@#4EMWWb�g�?��^�-��Z�Y���x�e�vW�aˤx�MOHQ��^n�\cDt�P��`����1H�	��y��j����e4���ȭ���3vț��b=�\&g�\�JP��_�Ԣ�R���_h=�����bX'3@�u,f�<��z~��y�G�~���:ӊ�jQ�/�n &Ad,�L���^
R��_�S5+F�L�'��8?p6)�;��z|�b��F=�c�j��嬏�A5 ���j9�~�T�l~N1#�#�A��+�q*�f
T��(t���Q�.���T�=<��V4��{?<� �L�Uw�+�%�0�� �"��'�H��C�IJ`	M��kr�m����~;
��a/vl
� �[��6%F4�ׁ7�"s��h�L���'����h´NXJ��Sc��:5}ELV묏��&�u��OT���r��i��q�\�돀�H�X����[� ��~ O�~�f�Xh\�7x]�;3���"��.�o]��elg络�)��$[z��V�2b����	�{}I�=�dfz�Qη�f��6���lf����̡�rj��Zb-��3ɪ���b��d�C���*h��bl��8O�!8џ��ζ��~9�������K��Z���S�� oZ�G6z�%���� ���=�y�ɿ8z�"J�:�M��V��*�-=�0J��|��H�ꁠO� z(^⹚#�m6�ن��q�!P���<ܔ�N�8�����pm�wV	L������K_�:m<_7^��&�Et�}��8|�a���o�r����R�h���S}h��O8���=��*���8C��b����?��fs,�жj|���k�7򚕤�P!��6���H�aFp��*l�Gn�y獘�e��/����[j���p#r!\PA�gc�Օ0�{��	e�>;��
�1�,��	��AςB�b+�j��+�[w�9�
�J J:	�M���X�m��%��;ҲN�̥�$C���.$�øZ/���y��7�qb8"~g��$2l�k�{��@e7,*�E�����F�.Xtx�`CAp�|����@�l����@�?�^e+N^��.�����ʣ�x$Z��0%�z�&�Trݐ4λϜ�%�����T�nڈ:{h��B��� Ư�G��|���={�m��Y�I��p�{5.|mue�p$U�� �}vT�c�z�:�2�.��]��ń��Ną�l�1yL���W�q�����8�r�� I����!6s4`BGB���,�9�D(HL���H�3]��h\~��;,0���M����ѡ׆�&c�_�{.O���oe�"2�ޤ�C����=�9�F�aD#>^���3/��[�Է6\n;ׅ�#(�pz�!凼���\5*�6�X3�:������8+���Kk{���4�ݖ:�=�Q����zw�e���f�5�T���yh0��@�F�D�iӑ�׬PU&�7����l�-��T��M��Ԉ�A���&//S�Ni\���}��Q�M��.2J.w�W�f_�`���L?�s4��[4�QdJ�&�/����m4�:l��[h���{(��T���qQ~���$G�z�o�xH:܍�(��e���q�=�3�0�4-%����\^T���ᝬ=��W���&������#�V�rv�K��7�=~Ѧ��#��mN�e,z��1y ���Z��y~��t����*b�P=��*>Z��e-E�{x���f��9
h1�qF��.��9Q�!�<��D�*����X
U�%E"��/�$I��U�#8�����@ �r�p`�)P˨���!�S�2����x�r�[�?��vQ�]��nQ�i�@��&@�sl��c�<�$�&��z��ŤQ��k��5�O(
Vn�8j��XR�⟡|����jX9��Vj�� ���5f�ɽ����%�g:�����v��́G���P�/I�q&Ϣes���p�,<�^Vr>�/��Ô]g�k���]HL7X� �g�"���0��ڪP�CQJ�N�B%��(��Ap��±|g�E����,���<D1��4/خ�m,p�חO��۞v{]9���L�FB��N�|�'����A���-#�3)��S㫸4����`�6X���`��W��U��v�68p����4	�sａ��m�Qx�:/�zVð���Q�麤�u��/vU�8ŋwI����R[f�~�ݸ�-�^���Y�y#k��1��EpIbW )S�c4�Z]+dD�P���l��zGE�t�G$ׂ���U�
~EѤ��.�Y���Ə7ޝ0�/�4�ʋ�����㑨g�%3S�ؼ_��QV4z?����ŀ�Vďf;"�#)o��&Jn��.�H�6�P^ɼ�c��ٙ��j�'$$0�H��~��XM�V 7B}Y�L�9�a�N:��c���hB���r(�8�>����G [ �(�ϛ�:M��>����w�
��q��:�x��|��sk3���c��\@�j�J'`�O���FQ�F�G�V���-I	�f:А՛K
L��b�jxԑW����TyI����<ݕ�X���yM)F�7�aAD��e�2FF�ك`_S�]�8>�)����J�wQ�J��j��}�H�w���x�)Y+u1��1Y��]��Y�̎�#���S�A��p���U(�NTY�i�Cߏ��� �)�kxp�퉸�b��`Qxa�z�uH�w�0�ۗ{����'`�.J�
E���cĨ��}.A�j��T	��ܡT�ᆝ���9�vً�'��
�����D��aj�OA����X���G�����jɂ_D'5C�pp�����)G�>쎳<��`!��>�L�y~�Sy��^b��:�(_Spvx��$�s��*�/)�d�����K˳ld�����uc��$�2�<�}%��-w�R�`i$<���&)��+R;�8]q �E;�5/���4���:͵`/�`��ye��M[W���y��F�?���w����f����g����}��>�ؘ�oM�29�r���6�-����v���E�݇���[�N9>���Fs��}*�)���[����I�9L����'1������;?�y�R	��$�i낛_�ֵ�ޕ?�Ю���P�͠ cwo3	���kp�u9�Ж�F�ݴ�X
�����>�Z����EY����+��Vp��B3�,&�Iw/OGj)�l�y�=�����D���a�*P?2F�
ϴ��/sn�LW�T��/b?zh�.|�>�Yʷ������£-̓�J��)�捀P��v���K��/�D-J�S:��o_'�솑�r�vg�l�:����in�6�=�S��u0 �!1	v���q>h�`�<�����I�n@�n��ko�ҌWƆ �o!��U�� 5ԏ��ӽ��NW:�ݢ�/���]/�`J��KiC�h?��#Sc���\v9�M(ܱ��x�y�h�<��t)�!2��}����F�O���A{�����B�n%ګ��Om�á�������Ś���#����ҦĨ�b�:~�JL�.�ʒA�*!?�Ø���ˬ��q����2-3�5��6��G�Bio���c��>�)ɋ�+3Ȯ��:��To� �n攻�.U"ߩG��H niٺ�_�H>𔬗�������$W��h~?p��p��|PS7P�aF�<r����;)�!� ��_wSiv-c���k���q�Ud�����x�P0!�������օ :�������H�M����#(eڥ��|��]��e�}o�'?�K)	�k9JcN�۟y!P�,Sk��
B~~��.�*BG��,b���U&���D�U���]�/�V�,�Q8�*�D�$P��}�����/q( ��v��.;���Ħ1�Qٛ�Nr�����^9���F���{��!���i|����<X-��ME,fǚXI��8Yꩼ�oZ�˜�]��h��͂��~��[d�G'`T��2z����[g�}�ia,Q=mh}��?��ؽ�ɣ��-���Ɖ�?c���@�P_����%�wv-Ԓ��CB�Ʌ!p�Yٓ'
�ʐV��Ӱ@!])+�W������!�A�[�o��W��ہTH��6��-Q��hۆ}��79��L�S0y�)�	�m*p��������az�ҳzj=����)�6F���$�wkλ$1^��Q\�!�]�?X��p�����s�j0����xi������I]��9���d�f�d�!ST��)wk�}�:X�P�;TOF+�P��ڬP�y4�YvX�1ͷ��ןr���X�|�iG�Q��j�0\O��K��}�/��(�s�Zpz��r�ĒUk�������A�M�É��_	s�Q��4�+.Lp`?ck���fm�����&>Ƚ�L�K����x�ߖOZ�eH�xlg�����y����b��� ǏH����u��P���}�*"6
���]�vmP`��`��uڃ�܏"�t|k�lW|_/B+��)X>��0F�E���m�ٜ�����̙�����g���s�%��W����p���gY�RŃ�z|zfK��wK��SٳQ���F|Y����.�,ܚ�Q�>"�Dݻ����8y�E�}�����@�v5�����ע��G�:	Vx�<�'��\���E{��>�����7���07�A � Tپ�Al����ꌧ� ��`��j��ʖŶ���5s�p )�cd�NG/��UɌ(�);B����]n���pc��}1˟���ݎ�Qj�0ڪ1��'�Z.��Ŗ�1�0s���;C?��x�lZu7=;ٶ/Z����T��F���jYϾ
�Xэ�K������6˱�8 ~I�� ���j;ć9���ԙ��3���s���XW"|����9kGH�5t�yy]��rs:}��.i ����\���+婯 �
x���,v�C��No�ɿ�R?sv���Ii�f@Ht��3�Uu�hi�al���+1�^���+Ŷ�Ժ�d:8G�D�"���t����q`kY�TMܡ��Uyf�<O��?�������!'��ٮ5��B=��#�Dyn;�I�B��M�|�5B��}1�� @�����-�gs![�r�ڤ@F��q����%^;��~.�{j�x Om��|8Ć���l?�5�(���BG������0eaO����W[��.=��2M�Gm�N�u�h4�e�F�Ǧ���u���$?������CWL�Ȓ�^�k��O�:-j�����޷ z��0f/��8�
�����j�,pf��ی��~�(�eՎƠ���N�-/���!��&�L�q�W�}��ݖ��������?�bٵ0r�F��l��m��`�E�
���V���r=�9�t�'wu4*ʦ���L�`
�
��7���J| �WP�1�^���l�pG��H,D�h_�9�Ǡ�ߛ���K�5{�<8*���A�s�6W�!3�>�d�0J���͗�.�hmO���.���R�
�����uF:}�է��-�y����iXI:��v�;�VʒK�ߍ����B ���L?Im[lLJewU{^�UF�C����E�|H@f�������_��g�8 ���K�AH��p�rh�2
 ��/h�p���F�w����"�tx����K�WBx�V8�;sɘ�7<�'��_��~ޟp���cG������_�O{NE�+�w�~3C������� �Q6X�A�P*�����䀇�^;�[�����erP�\�G�XK����r�c���͡ޟ��Kz��M�H&U�B�U�<��[(~�@����J%�]AUriR����y��4��(�W^�^ \uQnf������s����N5� �;�Q��B���u�)�������C~jw{�!�E>�C�ޛS��D�4n�䏳�<pAA3y%u�pDŧ]w �Q�	D�_���(�t"�X�5ط����o�~@e��7O��ԛ�T9��$�4E�9�"��ϖ;D���M[�����ėOD�}ʠ�Y�Ü�st�o��[���#[���Z��CUU���*�Hm�nm&��%��;��T�K�(<��$�E�!f�����oG?a��Nu5�5?�c����xX�Ni ����_u+�0X�N��q��<�%YC[�8a��Y�"@�����`���~mo�`("͕\�g�����^��J�5��k�[��N�dJ��,�hT����<�x�x�`�R�1RP/�O��M��iR� �@Џb����[g��N�������7����J;��r����'�-^�"o��](A{<�����H����M����Zj�3�b=N���d�O�"�U[���N�w�*��B�I5�	����L0	?�?��t#�d�Gl� ���$�yO����zv{�{�ec����[S���	��vNs���<���������'�����)�t��[J�̜y%˟H�0=Dv�JV7��@4��[p�<v=�Z:�j?�����۷�dw��8�eB�9�r�s��{�x2�=��+�Cc�����ӵ71�(�9eT��ל�'��a���h�?����S���{�:�c�r���؊�!z�m##��j�Q2���/gq���+���'ʚ+�~��~(�� y*�^��0��(�|�p�_���/O�b��g�]��;z��/�锰_J����
��'��j�k��1�lI�l��%�@�Kh��iC&�պj=��F6��-��}E�V�$���a��5)x֞_��?���1\����w�l����DLa�~��,Z�F�o�ɷA�w���UНg�}�'%�>�ɦ�jr������AD�O����#�+`��%.7��띉���2�X�9)���ڜ��e���]z"��0g��Yg�>�yYQ�����rVa���;뮵z&���'��T��0�{����V@�R��M�3lY���R�*F��d�O"��'Y��r�w�HDM��ܱ�����<7�K�`̡��.8���?�����d�Q��Y��,��/�a��P�@��rp�[�"����y]T�S�D�ɦ��EU
����,(�*ouQ;]}xI1x0@4� �dþr�S�=�W�Tl��� �o�&�p�AD��>���5A�g! �\�k�u?��:o�oh�����X��>l��#f�h��܏zQY��%�O�ƌ�c�-��)����;��¿�9\��i��C���:kN�K�a��U�
��#�����z춞L��5&�*��RL"��7>����5Iݮ�)@�; �*#Y�;�m�K�9���f���E1��;�$��G?~�6[~*���c���H�_�0c��+k�(�1��2��[*���'�RcY�JȠ��;@�Y�f|
��T;��-Fl��'7��h�;����{����n����e�'�X���m$p��H�uF��х񗧰�.�A�����B����cV��w�z�@�*	����II*=|?��s��>�^E� �GK7�"� @����e����H�A�~��4�z�E��T�-��*�E��go8�х֕����-@����g �VN��^���N,a,3�h�-�
/?r�/�ϛ��Hn��A�-�ŉ[	�g��8��#2�6q_����a��n�w���lY�>�6�~�a&Qq%���2Mۺ��x��I�7EnL�+ ����lJ�A����-%� B�k�z|s9��m1�1i���Q�<YjRO�
�1jq$E%TBxt`�p��c��TNOi_���cc�������H����=^u7��p��Z��aP��{�e�ML�������Q.����������.��f�D��Ő�D���'���q
����1�Y������n #O��(~h��w/���A���'��t�XL��j(�Vf,���^%FD�A2Jw��V�����y;|���W�?��DRlDe�oZ�1�&f�F��Ė��Z���QazK��Q{ �-��C���'%x�AO�����$X=�I��?�ֆ$ �H�ĸP��Nz��r�KiQ����-�ko��#����D�p��j��It�+��O�=�ck�(�jn�t�͋�ͬf&���h�GZ_��]a༪��/�x���̵bb��O��*�D38�8��QH0Q����7H�{��]�c�I������l(G���?/ْo�C�{r�C�����K�gc������o���D��{$u0E�����ӧ&[!���]�AGc}��">f_��^o˟���(i:�-e~B��8�N/���R�s`�}�p5�y��+K5��uO�T�>�R���u��lk܅ʘV��zgW��.L����%�㋦Ckq��s�"����i��\����њ��8���UK�7}�ݓO��-��q\�4ڳ�<2�����X�ҡIM)`hBy�>)�t�+3� D)®�zp��üsl{H�=_�v㕛WH����Xj�BK_�)�/�a�NĖW�D)�?<���$��ax�c���鬍��fd@8�-��ǶOҒ�,�i����+=���O��N1L�/��[z�:e�獒kI��s�1�5��zFt7���ړ��Or���-�d#���Sƃ��|�ٮϒ�SIFM��m�˂'�u�m���@h�����,shy�o�\?���^<>�<��;�����p�B�#��l){�@��-/Qs񎅳�P�:�vW9�t�)�=�L@9}sY���sI��n��G�p�C
ˬ_#����d�V�,^SxH[*ms����@̵	ҹ�l�xլ�QO@ڶ������r^7��A��8g*[��8Е�:�Gz$
3U����l���A�h�!���z��*�D�Jc��`X.�Q�����Y1'v����*�O�̌}��p���R��/XmL`n�2����Q���A�E��a����uh`�.������Gk({�O�y"���\�E��u��0��ѩ�}ْ�K�`\���J+3�����(Ⳡ��Zja?�f5�S� �+]����b�r��x)P~��T���'>�t{����<ҡ�[�o+R�x��\s�&̶�	0.��4i0�:�O#-+z'�����6[�b+�Q�&���s��F,�[�O�sm�:����=�?Y!�1P;!��̣��v�&^!�y#��������)k��F;�pw�0���{����~� �Y6�?��u��E._f�z�c_q�/Z���gPܾ�Zh�L�a<&���9�
����VX���G�IF�U�3�Oȉ��Lk�+�>0�Y1k��3��ٯ�fۡ�
�֋\"���q�/.Lq�u�1���*�:"�Ů~T��P��/��g��Vms�2QԄ����E���A��S���W���b��Ӕˤ�\������|#Z����2������>�]Mb�
�B?��:���G����6I�e�5!�.ʙ7���׏��Uw�a��LH��O�����@���H�:Lu���4�����^�L�tL2�s�U�>Ѓ��Z����Ssg�����Su�Z��Y��M�]�-�"����_�9J"�J�y�"����e +�yY���m��b�;R��T���	�֘��Yw�	�#='�%9�0�Ŕ�z�O��+D�%I��M}�D�M�s4+�.�J�2�/?������Jq��ß ������E�PX�o��l)N��a���7�}�B0� D�����G�Xc̴B5��ڎ�^A��ϧz�T�P�Ͱ(�MܬۈX�Z��MQ]V��<�M-�a_�U ��CK��L�A˴y��?f�=�mR��s���à��8����ܚ��hh�Y�'p�V�����[�oB&v+�
� >K�2��w��z���Ȧ����N�v�Ȕ�o>pZ7��f��� �G��f���+��h�� �C�b��.�tJ&��S�D7��PlM6��BAX�B�O|���0�E����PY	� ���X�;�S�P�T�`�6�,^�N).��xW��{��}k�m�Q3C�0��<�I�;���XJ?�-ܝ��MnTRV"0����C���I��HOXE���;�"�g_:B�6	ma� ROA�L��:w�2�Y�ȼ-�CtXb��5�p���Am��]�:t���� nׅ(#Sn��2���[��}��ށ�i��[��%ش�}9`tRڽҩ��^[ĭND�m�w�<�h�j鐚8&z�H�`-$K��D�,�P��;Ͷ��j�Ś%

��}����΄4ս��]��áS����z[<��|o�~�r����0
�T����V�R��ƣ^!�^�}��kQ�����>�c!�[7����Y����ڸ/-Kok�5�z� m�R�pr����lM�c=�-��M異p"���=��<�{�Ró�?�X��`�\�t��N�yP6�$�0%�Zr �����Zq������}L;wu�bG-�7#�y���ڀ�p�		�9g����p��� �@���<�8\pɝ���� �_x,<c"'����z�k�G�3�(�	��o�ɇk���?�����c"�����m���ӕԨ���3��k��-����E��85�9
:]����`̃���3������1�$i��\&���
%�49�]��9Α_�R�RI~N�x��oה~H�zu#�6�|a���d��������;�����FC��K��zw�)n�!�hre�~:�];����..5#h�Q����(Ŗ�	���#Ae���r/7�s��C(�<��tEu��3�tv��£uՅGzI�� ͂�LޜF@�W=&cQ���BQ�#��+�m�d�h.nSލ�L[��1݇�F6�j$�4˝V%j�s �c�������B�p��s��<Y��.�Uֆ�*	{�Cg�t���z�E��z]��t�k��g�<��{��Ƚ�4�����*:����\=t}d�;/��}�����d\bq�5��E���)  g!�<����'@��HҲI�6�w+q�$0�������K�H��W*�9���b-R�"k�З��W����wˤ���3r6\�R��y��'�gyp��q-�(��]G��3���������Ȅ�S�O�8�����I�Ƌ�U�HY$��9�9�q�ۢq�3h��+:/�4�؜�������Ug�|RԦ���%�t3f�V=��|���N���2�<�l��R�e&Kݙ�̬.ߛ���ě�w]H1�n�����pd��T�"���o�&�Uᓓ
��S`W�"��fN�IΩb�?)~P����U���JX*�+5�P�b�%�Ab��2���P��W��s9�_|��Rz����J:�IV�o�ڦb�I�oi׀�d���~v4�D��%=_-e.�b�k�Ws��3O,������d+��>a�J�j��O�"a/r����0�7�%I )q�� APtՒ�fL�#;�Á6XK�cy���)�"9�֑xc�����}
� ϭ'�]D�����ԊT����}Bh<?4L�΅�6������֋� ��C�َ�U�U�"?=�i��䬳 �Ӟ�%d�!*k���7�t���*?��n����hԥ:q����s�O�y�7$�F��������^��b�<�)HY �h@��?�< �o�Z����^[�- ��qgx�$h���Yxu��\�	�u��C@*��4B~&񊙚�K��B��+���6�B�Q���a/�;%񓐈�(Q\���4���e������{S$��W�`=AW��L2�:��z!}�(�aC�!�]��M�C-%��,I� e�_h�D���.~����T�d~�
Ұ�7�����L�7e��4S	��Ŕ�B�DRz�O��C�� �]���6��>#j \�x���yO��v?��~��pZo� :Jԭe�L>���A��CQ���b��¡I3?�^�^�������[��6Kn����z�w��Q|v"ʠ�����&ΨyZ��� ƚH�,Q�m�)��aX�����4�1J��De�9ůy���!�!��2��� �J�L�M�nZ�d��\��F��ؓN�Lq3���Dُb4��L�����v�8����<��	<z���Ǒ�+X�R�q1�iZ3�?�\,�DeF"���`��8�*����[nYN����Ad�p��߃�<��P�ؒ���#���ݷ���D0P��Z��񂆭���B"�i�.�r)7��=8�.v��sH��ʃK���jd�P��%��)�d��~=��1�I#��$2L�z�VwP�+�N$t$��>L�8k`���@R�Û��.ND�9p��i�җ��>�	�s�t~s<!m������추;�����u96��aB�^w݌��d�;�%$V�e���
c2�_�c7Öᨖ�yIp�g�j�=ؗ;o����v��	�����'SdVO���Y�丮��m�F�c7��0�z�\��+cx��o��")�H�uEַ�� h˳�x��%c��_9.�f��k�=�F5j�I^d.��ҿ�T��^p��0�6�����7�83xI~����N�Yfƀ����>���c�"���4�����'�/�U继�ۦ��B����${v0#P�Z�-��'ڷv��C��<�?�p��v%�V��K��D������Ū�� �[@_�{)��Gc��N�ҰA�c
�3�+)�k*�q�|�-�}�5ץO�m ��52��g��@��T�%
=#��Nd�@˃*=���;�~�����A|��Vt�u�{Anv�v��+4�<��Nv��gdrS�����f���[ho Uş������
ڧ5���&�5� \����!��l}8��c2��=�M����r���"�o ��â�$�ُ�I%�H�'C��!�^�_���j�w�	BY}L[�C\Kaa�b/�	Gy��G��'��P�V6�.�Ɏ]�
"���Q�[���O�[�@���rW���̜+�1�4�h���/9��/4C��'"��c�Iq�DY���0��4�J�H!��l5-/�J�x�v˔>Ƕ��3-��e���V�M�!`���1���,MWݠ��ItU�~e���wG}h�es`��ZàUrn
�!�:��V/� �Vp1����_�g���D���NA�e��g�~r+��{|��eTZ�B\����Xb�`���Z%[ݘLcjk�h v ������Ef���<��tL)���;�c^PD�aGkM<��?��.�}P�f�a*a��dZ㦬��*?�h����(�I��0_6�.�4�p��c��E�E��c��5J��Dxd�Q=�mj�W� J��)�D$�(�<�}�f!f��];$�Ń/r8�����S(�&Zw��y,Aۭ�kύ���3���,*�Y~Ϝ6cY���v˖���
/�#�����0��~#��A����<��Y�z���q�Zo쬞,��8{�t�[�E���l��I\�D|C����J�g%�P�r'V�u��y����&��:|�}�	��O��V�ˢ}q�e]���P�`�u�\����K�g5MU���գr��y�1��>p2��{Q{0wVߕl�nV�a�1&��i���]ͮ	��|HI�I�n(Y����fB��]��Mn�N��ړzF`E5����O$���T�b�DW�s_ux�_�%m��6��*��*Y��ǔ���:n�k���nZ�Z�A�w����Ij�lqK��7ǦEG�x;8��q��Wb�]W�?d��m\����h�o�B�*P�GB,Һ��T��mZ�Ck5^?�s��Q�q@���ܫ��%������&�%Jp��̆�*L���ь���Ma>�����O�`�<T
9�<S[����d(V�Y�%S�.�� <禎��-��4t/̹pH�Q:M{7%W�:>s��I��T�I��5�H��;�ɐ��É�=v�Q1ۻl#�������}W�����3���>�?��@�X=cpu:�bt���#��'�os}�
*�x�>��P����|Y$��[c�;qg�"��a�&� �g�AϾ]R�DBP�5nG�����ܗ�Lc�ñ�;�Y`�}��V.$�IK�%�◵3�2o��ڰ�\����>W�g���ۦ/�\|'�O�"�J�mV�66���9��n��0�M@���r�D�«�_��֧�X��|��e7r5��%w��[-��!�ݘa�F<����vxA-$���ju�g_��S�a�>[�.����-#RKazL��畛�\=]3l]eQ9�5?�͏�v�������7�.B�q�	�#����{��N����_�'���H��v鴷}��8��u����v�����p��׆�Q����mt���!?�����ҵ[����`�;fѓ��}�6�<�Ҿ���\��<so���jF��X��Q2��R�Dp���(^��e�M7������K���!�}���k����+�0��oHB�o0������΄9P}�h0�[�w�7����#߯wǲдV�B��ԅ�]MՊ��qR�S�a�}�4�Y ����wf�r��!K�g����d�j0؋��<x�#�s�7l �	O��RL���jhs��J&�=�[�����+e�t+/�SVx=�Y�8�g1,� Ž�*��K��$�:�kS�o�<E�V*��@6�_h|�J�fzq�)b��ˀ��B�xj���SE3�Rٴ��I#h|�����	��S���̤Ս�B��bPͲ9LJg�:� NT�y����{[߶�f�`~���t���U�A��_VV�M^�J.��~�-����_���L�B3���t�d1/p��^GՃ��,CU�>��S�|���f'B�KT������8
�,K�T�!��>J'@<�C^lN(ʹ�-3�Hp������U�L�-u�K|թ,Ȉ��֌B���/�Iݭ��c�5.�ԅ���վ��sKaATQ[io�m���D��HO�&��,�2�>���p�J��M���a�゛�'-)���U��K�f�^OHJj	���FA��f�Hvq�
�fX�.5%A�f�Gx˭76�q �*P�y �"�֊_)���Eۍ��qu5Z�Ps�)5�?�)Ӟ��^�=��b�ekZ�"�X=]�L��G�j�^�~ҍ^V:?ϸ������6�4���Dq�T۴��w��m̢I]IgZ���c�:X�8ʥ�ܧx����K;�U�F�<����UU���U[�M#4�*������B���xvUܤ�R)�=J�o̷�}-�W��qS�a	1~߆?�Q̶��oe�kA]u�G����D7�J9B~�b���sb8K�܋�GhM#Ƞ���D�i�6�|&U��㰂H��y#?��ge{�xղ�s�m��U�"ł_P���9Zսb3�l���r�ddD9�>���z�MAN\��N�&aDl������@*ܰ9Ѵ}D����`Du}�o�/�R;�0�
m�D��s���0����et�쑓�=�u,����CO��]!����7�7�_9����`�"fM���D���㷈xc����Aw�sN|ؾP4�~�H�
��1.ôX#Ƣ�x� #?�m(�uY�s�EK�f�v*q%�2"�u���&s"�Z�H��m�&Rf����縋�]W��,Br�������@/���1� I�V�Ȓ� m��h�0����?�~O��6rcd��%a�OPN[1q�O�Ȁ#��\Lz�����ֵj��l~q]�x�wPAk����ۙ�ꐏ�b����|i��x��s|����2�j����\���B8c�v�-V{���u�^)9Q�M�z�)%=�~<<��	n�ba'�Q�����]��˝�����!S�t7D���vԭ_�[�$KFѺ�d�T�lt�Ju��!�&�7J�.'����܁M�X���a*i��-MZ��m���:��w	��EN�_�9r����OO~�EA���lgH�0��J�d��ߕ�ʳ/�k�¿F���e�ȡ2.ɮ[DI^�F�)�SH���r���! ��:������?�`r�,����\��j=�-������'QrY�(� ��G;��#��D`�%�15jTv�/S����_��{����y�1��3HD&D:ۼ�X�����}k-2Q>M�"p��3�[����9+��x�Śty�K/��	#�Ѝ���ʨ�Շ����q�#hN�Yo������=^��11���!�p@pZ��ZFލU�I?,�;
J்��CK�� >�F0�B��w�U5P)gK�6���\{٤!AC��I?�R�G�իM��+��q�����A1���e�TT��P��W�V�PE8vٜ
e~�
(l,��!v���N,l(��u��v$ٺ�4a&Bj�w�^^P�x��Ə[���w�D>�}_�0/���r"�d��?��� _mY����Vͱ �����H�UD�Bu�rT���@&�cC�{����^f;�٠ qA���ea5?�D̩�B��'`Y�:�#�/�oPMN��
.�d@,��Pk�_��S7{Nx.�1W��$%�Z9��8�hpZ�ͦ=R��nӀ�c<}������RQ���e�����ԍ.��p����Ӿ��5e��4/�g�{c�Q��0��� �(�3��r�a���\�)/ݯ��]jj Єsl�0�c]��R6�s�u^،�������;���8V�{r�Pn��Z�g�`&w?��f��~'� BVr�yAN�H�<8-��aΆ��9`{���R���Ɍ��o�OoE�k�hI����kmU�AQ%�;��*�.�!>p:��Gբ⻴!�MU|���!�[V-����W{��g8�}%ӛ�_l���s�(��K� �<�a�7�ak���R�;��X��-��*v�*0�ÉB�)*ZSGj��*x���J���j@"P0UF�����Qi�z�,".c�����U�t�ћ0�*}��,v��RW��$~���t�'qO� ��2e3XļGgLu�i�Z�5lh3���6��}�R���H�j�`QI��{}R6�����{��R�'"6�O9`�Ә �M&~����xV�p3���װCr�� c���^R�w�Ltu�)�
�z[/ݬ:A]�Z�L9�l`�1�l��=F�'�t�3���� xC*%�&}c����L��H2P%=��c-I�j �����#A�6��1գ���V�����5R�/���^����!�#����Y6�z���o?sl�xj7"��=?����I�MwI��ZM��ڹ"FgJ[�w5lf%��Q��5W��=y[sd��v����n�.�����_�+�yJ@�G���!֚�P���.i	���P���}��V-e����ᾼ��a�U0�����L=���Z�<�G�/�As9~�XAT8�Pq�9g<�^S�0�E�!\��SV%��5ir*r`s����:�S�`��%��$ʏ>+�,���K�(7=%�9��=i�B�Y��$#(ۍZ��
gH�a� �o$/�[��cd��|R��F�C��i�D>'98�^
�uҨ:V�z@)'�Ӭ�s/8�'Z�^̶��� <��N���(m�q`�wQ��_�,e黠&K��n��X>p_p5�>����1 N/�5M��Z��ox��A��*i#ʹ�m/�HF2&95��*�Z��[[M92�T�������i��*�M�lj����h�a\�6�HR��PVI���`&��^�{!F_�=f�P�/�C�\��a����ߺ�oZ�x��l�pc�&7f�+�IL����x����Nb�i�2Y��-�a1����ʷ0T�g ������nm�C�GHC�r�@�)� ����dx��B��s���
�+C�\n�z�5t���p��7�B���+;����߁?+����,�@�E^E���)�E�-�Ma"�^�=<��Z%��� !d��ԧĤ�X�Vhֺ`%�Ds�HB�ޝT��f��6�����g�%1W\�=�_�x6@9\�����.\ePֿe�zI%�u�hS���G�r P�H��'+���퐡ģ�H'$0��k�o���^ؾN��oB�b��8��)
��*�sC��1��/� ��7)%O�dF�a���vW�fr-��:x�pM����7r����q#b++Q+	گ�κx�ac�� �����o���>)Ǜ��cJO�u.�X�G|�c��8�8N۩�K�v��`J����X��z]j*^�,XZ�j{��c¨�%_C|��Q�ׄ�i��q_����
��f����*��BX)ɇ�@kuz�4�no���86�����6�C��ks�r�Vn�ԩ��n/��S�k�v"���W��W��Ѥ� Aj,*:�g=�/�9�^��!L�]p�i�y�m�c��}���V��`�����k�qS�Yb_���-� 2�<ϘM���*xW�!�����PL1���؞�N$��g��t�i�]�d.�*=��*���%��᣺NA

5�Z׮ǚvHi���������Fd�:]@��H@�L��>���q��si���g�K�/�<�.*�r�C��������&�O&�4H��4���,չ�e�du��	uJ(�U'wH���CМc���jjf/["o�#��V�����m�1a
���2g����i�������\K�3)FPBmt���n�NJ�@Ό]6`��؋�4�=*��d�v��T֮���	���i��}���A�|lTg��Xx2�`n����^�ǟ�X�k�ea�	���m����gG��f��	�� \�vJ�<�r� �D1��"֞ r2��A%�[:���)������9���=�N���H�O5��ls�y��e�`��� ���4:��?V�{�	߷.=TJ�Ѣ����vB�P��Nv!��~��X��9 ��¸��س��Q�&>�N&�L>,��f����e�i��N���K
���(�FQ���_x��M�nl�I��0�r��M����SJ:W��[D��=��e��h��^z�g�ٿ��6.��B��ǝkn�vwa���!ߙ��;���=]�4~����͒��e�m�S�x:�O��<*��\�땅c�P9���ǳ�cc1�m�?h�ƛ��r�iW��%��]����S��S>�a%r�Z$�����ڳ�4|g����:��&�e�$�T-$�2r����#�D<�d�E�����2��˴�x�!��]'F��:#�t=�|m�w�$�?:6G���dU� !mБ����q�����!�՗��.i\��QZ��`��pW^/��_����x� ^.Bz,%d�U�,�H��U�@pmَe�E_6/<��f�6'�Ai�xۉ����Ï�xxM������=�QU�	���(Z�,Y`.B�5�C�PR27�(�+<��B17�U�D��">�+�z�O���k.y_5�k�!��<a]+�7�ϡ��2:�h\\�z�RW�r߫��C��N��f��xP�4aF�7Y쑏��N�m¬��i��Dn������v5�"��Gx�~�Q�&�A:����\���|9ip%#s��`�����ܔe֐�sB��fA�fM���#u@x�\���)�W;忲1�����?�Ѿ=�S��u~DPT�aM	w(#�lU��UXx�eG����DZE��"t��)4��&�t�u��B|�����5��H��x�J�H�l�>A |�����]���T�bV����T�1��Hm�5d�G� yZu*Y ���l��NR[�\�%�3����͔U����y��}GwE�ᝄ�I�C���W�L�E���ww�#}����5�w,۰��%b���9��<d��N�y�1����O�ѺamO��2��w�X��6�Ev�`lW�u]������Ҡk.3<��O������zy�C5�R}; ��t��	of����I�&0��~�?bp@��nM3,C�P�X�v� ��Ӕ5�GW�3Bz��ii��ӕ����2-+�D0�� @�k�	�c7.����H������k	y,}{�C����Bڻ���n�G/c��ޘl�q.��F�������X�gQ���]N�MaGU&w��l���47	n�9IR�VND�O{�|�}�.� x��.R��a Ex!��N;���.-��o�qj�VCɛd��QpҖt`��,��d�R�vU�+_Q(竧u�F$8�M,��/Z�QO��}�>?����y<���:�\ΣG�E%D{03�ϩGL�qs��#���O	©���b�����0���{��x_�!G����6(+nˍ���8��P����	��u��&Q�1���1`P�d�644ľ��<��}�V�^:�(�%y\ �_�k/��p~�}�u
�ý�h��9��{��w�8"�\o*���0n�a��>A G��L�2�<�d� 5���*#�j����b7:1 չ�{M�(?�zg�C�)�G�輛l
��$1��\��8<U�8�H��G�V�=��z�H�zG�p��].|k �L��m�5 �~��Y��r}S�v=�w����i4�y{Ҹib�p�U7�p�W���
�KIx$������d<�q![β�2n6p��j�\N�ŋ��꿒|�u����R5[�w�;v�~���<��a�*K�M�Y鬗w~2[���G��O.2D���*酢>1����J(�^u����7�\�se�!14!��:�NY��tq�Zw M���W�&��J��m��I���p���6	M4���҄?�\A�_0+e7n9Sw��ǫ�<�~
*�j1��0yH��)	h��Q�X���C���ک��D٩��m��|F���fgy�d�6e�nA�-s?�"
��b�s�����d``͞؛yG3SƘ�"���o1�_��e�� �f�����ᷟ�d_���3S�-s^[&�o����g?�+@�U1@0ߏt<	�rY�BtA\'eST@l U��ªκ���f8vѱC�3z.}���7�MX��y֌�@j?c�2Ӊ��# �rn��]�BLhGŠ�O���:�V�LX��$@��	T}������\��:��+�F`��&���uIY�jI&o�c`4n>���o��(�o��E[��61.L����D���-U'=M�V������J�����K��2~�E� �cQW�ձ���q�kƽ�en���Rq$Xv	�����N2d�������A��Y_I��:�i�_�� �)��0�BU�������s8�I|��A	<6׹i,	�ؓ]U%&�����1�Ju�bZƣ��醙샥���>| �;S�2���Og��\�d��}���~%k��V���T���o�����6=,-�u8q�(��.
4^m����\�����v(��N�̽��OᲰn���*�
i�p�'=�F8������e��m�趇��
��P�eY��ܯ��u���&��k���%��l܎,"A�l��"
�a�`��rh@���7'.Ǵ�(��-��̘j)ü	�]��T-AW��yw��j�. �M	K����ǝ��i�f�>��"��N;r(�z��TL(K4ܤa�e�`���7^��a�[ǌ	(S�n������z.����T��#�	0}6G��e`��H��#�ϛٍ/��
ϗ��+�rgl���PK�t�1�L�_��yd�D���>�͈@4��;)�ZAI��3�r�6�U���)t�{�¢]ĝ�jZ�l�=&g�/�8����XC��Ǩ���K�HmVt��%z���O,�}���F�I���F�O�Z�3��2cF������6-n�$N��+�{K�RF��O\e>OzS�
���=�ى)C�K��&��@�&���� L?�N��-W������9���|5p:�����Y N����%��.!��S!���*�kKvK�U<���#0�fX4�U��
Y��,p���[ͼ��g��� �L�R��� �j�7�M�b$Ĉ�7=��ԡ�f��������6H!�����J�bFcד��f�
��;&��}i�R���t���HY�d �?]q���7~�
��]�jɃ�<�>W�j���#�د�h��c�񗏟�ǘ묓�6�P�_l�`���ӥXN4Ӆ�Pu��E���9����?,��\v�2�k��5���3u��)�n��|�#P�%eDV�t�����udv������r<��jX���d Oq}�"ú��Ǚ���A>�&1Uj��}��Qy�Pz���*I������w:�w+gn�.�v��]BfE��gjn��ٓ)��ϔ���9�:�c<�ZU;ʃ(4��ׄ�U���d���Mrƣ�/k��/*3��c���=|�!�1p�K�f��"5a�	X�E��6NoP�䕿>�L�]��a�4�L��57ߛ��ߗ1�_W���>� Ke�aLc:�_���Һ@p;���#��8��[ ����z�~Y�#��,����/5���lp�s�*˼K�RU�eC���
A��dF�r{��c���j�Z��&�jb��q�4H!�
��,�g��4)��q�ʟ�u�h�r!�a�"7�p�O��C]Q�VCO�(]5�&`��F�&����l�.V]q��(����=��2�� % b�b��auJj⺘o���k ͆Lt�����?�^���1�o�lV�7�_��N�ӱVh \y3�E7yQmt��s4����U#�S<TYgak��cdg��{mR�U^�����bȅ#EX�{Bȿ�g������S�8��|�|�0K�8ۧ��Z��!�����v�-�$���yR�'������0���y4�T���W�m�b�����n�c}�Bx��7�u�Fh��	s�"�lz��$�J���.��%M0�A��s� *�!������v+�keܱ$�
$���`�P�5h8+�n l�:ކ�W�xk5B�3 �ѣ�\��;jt�ft<��eG�����Wտ�Y�S��f�H��H��a�Na�l$�/�踴��	g-:/������R};��|B�ə���3N�3����Q��{�,�)r#��k`�vٗOЖ���T�?U��O��TW\��U��_�W���Ba�bέMq��-�VT�|�|h�:� ��Olx�7ʝ��#&gŒ���/+&��y��S��o�7`��L83��ó� ����stw4i'f������hPA�-yȋ�H]OLN�O7Tõ����_Iu��u���z3r5-�"���G�P��U!Nѓ����$���;<'�!�)�Ѡ�s�:2���0,�1�����A��X��Ǜ%ÅV�<���м��Зg<�Ӥ-ܒ2I�<�33��XZXS�E�d$@5|t����P2~`�ؖ�STg�~�Ş��*�?
�m��`w)�;M�8җNR�m�u����A44g�z5��t_1O�8�L��5��َ2���d�w���x�R�0�6q���,/��+mL�u�y�w�������c���
����Ѵ�,om��M���eO���<v����Z��$�^M�06��E�[�.�qܜ6Dl�tU����J��#Q��}_㟛�
�	�.�V9ˑ%�	��k��i���u(b�ܕs b?��P