��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��t�`%�	�6g���
�%_��<§�I�j�&|E4�*����k���E����;�v>����p��: G�Wٛr��j��lHε`JB�I1�W�@Qݗ�gM�*Ɓ�����j�Y~5>Q�/-�V�E�s��T����)��H^�Nެ��l-:��%���1)*y����=7��a G��Ś*d84�:���U@Nl��,����p�uʖ�n+OT X|��۞�&Ƣ� >Aʍ5��P7��{Q>z]iS+�������6���V�h�ʼ���J�@�Ӡ>��W��b&&��khB�S�S�+�ܯ�T�ɓ0S��{e� ��"K�ct�[Ƅ�p�7�������F�s��E!{n��&#�8U?���xr=%�l��Dup��G�f�&��2978�6p#���V�N_ń?C"��~g�?9���:���a�m���Q������pa��#ߤ��j�u8~��|𺁭�Yג�>�u�Ծ=����D�ұ3\��IןS?<{�(
��>e`���fJ4FQ|�q0r�diB���s���	��B1�u`-�:���"j�.�+2��O)3|�I��𲽟�����$�V��{�T}l�2H�R���G��r~�|:R�Aə
��vȍT��\2�D�@�J�U���#����2���$�l`�Y���(�q�m�m̲[/�׃$5y����9��I���+��
��۠�2�v��� ��0��M//��hL�\��{�X���:A�#�
җ��$�̈́J�f9͜�^�d|%N��	�w�ҼѲ���<F�::�;��3�s�P�舌��2�O%$
FW�`����������S�4q�E���a�\��A��H�m٠�<�p�ZW�l#ٯ�p�Z������z�;y�Q�K�&��~ nu%θ���{F�rh����g1����.	@ʞ�����9��Wd��_�qE��zbF�p +�1<~��I�D'�s�dv|���(�}����WE��5xw�<OY!"�S�v�1S���/{R�B�!������_��
�^欶���)>Ǚ�M�RX��In�haX�7n��^�Y�,�
�����$�o��q�$	Bg,W1�R�)�M�hО`���#4[]��a�/��,�V��Z6G�ҍ�����=;��I����<\ �`�H"����T��h�w��h�Q#�y�u�c��R���G2�!2?Q�5�[I���dX�fz�I�!\�C�f�\��20�v�K��K$�uҚ��(���j�V�,$�|b�{��'Gr`r_�[Db ���8��O�znge�Q�U=��G-�3�[=-'�����c�0�YT������,�;�����8Iv��	��.��$+p��O��lR��<�p�Q�=	�Z��,&,y`�����r��=��<�R ub$G\d��圫|S��M��v9@��[�cz-zx����D�p�+b#1=�=OM���@T��>k��/��������,��"䄁���W�s�p,�[��q�`��
������Q�͚q���2�F�m�nI��;,
=,�`���C���%�q>Om �#��UL/V���P�xV�5�B���F^[K9��ȖZ��]5T��h����F��#� |�1<��ӹ��7�����0�>��N8� �����U��^B|f:~��"��ޯ6����,|
)w�))0�C���
������kxe��B�U|�no�M)���c/v��0�SG��e��+�]"-�mӸ�a��jC!IW4�^������J� x���.�#=_��X��x�,��k��0���n�abc�f��)���}�OY��NI)n��d�v�����*0�z�~cb�8�Oh7�o`r3|Z���Ax:U��T8�!����rtخ�f��h�~ u>J���J�i׋ֱ粍\ѿ��`g��+X�0�R/NW�xԮ�L��8�w}�ʙ�`!9��L���<z��/���C�e���9pW?2ߘ��a��l�'�=��ˉol!��mx���-��A"�$�����;�����S��y��xP��S|f�/����oc�[���KM�	�'�*&�����he�1��mmc^8J'�)�v����(��h����D4�����/0�l�ֹS{?R�2p�;o8e<o�~�z�R��d��V6��l{`�	���6��OV9�	Q(�A%x����(W��0��$V��b�e`�p1�lu�
�60�,M��/Qڥ,͈�g�ΦG�u_��HՅ�����j�8�*�[y����~�<C�j��:a�Xuh}���|��T�G��$��MQG�Č�A?!5\s��I��a�A8]��ݧ~�ι��ꦕ����{#d��"�h㖌)���;D-+���/��iH[�d��m8Dv��ǖ9ٻ�7A�҄�p����[���ǔ3�[}�]ƫ�5����ԟ%I�N��0:lY��B�r�)I	���ޢ���3��F����-E��(�N�,K��6B��O��&�!�g[��`�������Mw�/$Y%��}Q���!�j�2T�d���9��1t�~��o���z������¬ o�j� ��|Uf �3�YV��\aQ��HgpK�}&������X�b�P����.+�4�7	~��?�7otН��L�������36G��t�=4:�k9���c����F_���g��Κ7�H���x䧾9,
�2�F����Ky��z^���z���GW;�b[�z�R��o�?] �YK�R"�6�a��I�Rv@�[nVT���T��=BV?�'f歐�iZ%IK��OƦ�iaN��9#���4N�'�Sӆ�e�ŕjC�5{ĥ`C��7�C���ɚ]�}d�T�/�)�����6'�ۭ��o�;(��]	k'�׀%�a�*j���pc���ݝ"�o)���s�UJEX��`Ͳ����[�����۷�͜mt�V{�؊�Ɣ�
�㏬o^)�-8nQ*�Ȕ8e!^pF:za;�;#(�SjZ��E�-������Œ�&���pE:���e�wJx�����=��>�����=3j`<�3���(�F(7v[�f�w*�)�|,�/@r�5I(�!�!^�O��a)�����I���Q��C���Fn�p	x}17JF: _�s������$�7h�җ����r�?���9>۽x���:�aZ7l>���Q��E�0�����t7i/mX��_�9s�m�����
��]WF�c{�.~Bh�Y�Z�6�sgL�]-�k�}��Ǩ�F�+l��Iz�$�0.w6Q��H���gr�Z�T䨖wG����S��!?ux����|�`gS�.��:	��v�e(�$?� _�a,͜�����&}u��(�.�Հ����w�8�����S_��q�MS��>�5�ִn^i.�A+������au���nU
������2��`�\�l㦏��ى�d���[��#�ԅ�k$��#8$9��?AuYJ�E��g+;��ǌ���8�,UQ�2_dL�������5+�e�O5��l.~�;=��І���5V��%9�E%����R��2�k��Ѭ*,�Q����z�5e���+ͫb��}�����p,Th������E}�
�H:����"����q3�j=�F"<�p�?%
��D���ew3��
M��1�@K�sk������rĮ&ZZ���:s���]yW�e%&K�f�K��3��Yk��g����C�O)����ݐW��0ҏ������O�fl0ߏ]�/md]�:W�\�ʧU������e����Q�y �����c2��ZS��Ȼ�<��Tq:'�*�n$�O�I5�dm�T��R��G�v���H���,�9�Yl8��	Q�7H3�F�|�+�׭����c��t�Ig��z��	��^b�L]7i�V4> X���,�2�gK�;E��\�~��W~���"�'��bW�Z���O���e웟���SP���O�a�\���o�I�pU9!�"�7�e"�,ڬ3�^�_���z\�ytD,���Lp˩���%o#rV���h�X���^RK�����-�D������.0=�q *PN��85��e�uQO�/Q��s����E�F, ���<�c@�}�č�`EI
;�l�.��t��Q�d���(G�C��O˂�1�Ys��P,����"d�˳��.�"�k���e݁�*Ɠ�2�_r,��t4�'����=�2
�K� ��-Q��?9k����eD���O�-��9R�O�������= �s��y���I#s��:$Y�לfUYߝ��F��z��g�D�-����N�c��s�ݬB~�Qr	��ӊ	�K�X�ԟ���s�X6���R��ކ�-�j5rL�4��yUo�E'��Q����!{�Y�����s1��)���؋@&���ڝ��/F
$_��𭛄֯P��"��{�<@Ϝ��0��J:r�1�oc�~'L�=��"!@H�2 �bt�zR`�����=4���>��ly���Hk�p4����f.�����ז��s`+R�8;�t$5J��i#�)H�5���\ ��ܲq���;�/	Q�(A���ag�H򩼥���z�ڋ0ы	l�&��S�4�$��~�H
'�E-�L��vcڲ�G�By��R���Zg������]�<^+���,?|�\�1��Y=���3{��"flrRW��o��&+�ૂ̇H��o�mg?�˒TB�n��-�ݙ$cZ�����w�U�{J��k��+���r�NLw2��}�J�>C�A�^�͈ i����#�4�k�P[c�rS#�u�׀2�3p�Mۗ8�
f���[�os��&���-vb�F̉�xГ+BB��Fv�CQS�����Q1@hl�y��Z�r!I�leb�d�i=c�I{��HO�ׅcd����h(�򇂉��?���w\J�Н��{��&��T�t�NG�����ޛ.����7��-eH��s"=��h�X=&��isJ�^Ҥ��]��b:(�y�uP�9�ު�fr��=C3����d�#x;q ���%s�/>k�^���5w�{l�O/+<��75�i�|2D��u�*�z,�ǹ�u|��i�>�xyu;@�� a4�.ϐT�r�e�������w�@w|t���5�4������)����<߾-1��Y!q]�܀�=�-�}seZr+p�~m���D��N �%�SY�Yͭ5�iY�K�zg�3��v�\)g�H|9n]&��t:c$��Gu�Gk
����*$�A*�7��������ڂB��K���JC�S�"+l����2�c�L�M�a����'2l��yl�d�J���n�J"��7��_R����&!+�V����*^D~ga�����}�&?�K18��Af����/G=�GsPˮ��Lے^E֛���j2���<�I�5)����{�=wh����J`PЯ�{�;�ܞ�� �x~OjW�}/�l���_0�h���5�a�&�@NME� p�ʣi\m,�z��g"���X�ǝdZ�[ꚷ�|T��<��f��[���U�������KFg���[�YWC��e�h�hO�g:������5w���;��OHq-��W���fZ��^ SO�.2D���d?s^�`��G���S�� a�&���|�$i�T��xS:k�{e��r��$�cU���'��O%���!��I���)�=E��l�S�!9�Ek���ӷ1�mӪ,"���:�����y���ٌ�@��`��t��=^�'a���Dq�(��.�^����А����.p�U�\fΣ�+r�84B�F�A�<�W�-"&1��6����{�t�v���Y/��w.Q��Vmc~&3'�2�aT���5�5�6ŗ.��d���@�.�Q�7��.��A*����ť48�G��	��P੘.����X�v�\�M�:d��M�΄�){�c-Ur��(����Qq̣]K��Y�m�\��r.s��T(g���F&.U�D�,�ԛ\�qE��Բ^���N�Z�-����`s�"�G-,:_>���Zg��M���e�eۦy��������$L�F���r:�<����Sl%�t���~X��|���UكM��D�� ^����d�J"���j����>?�HXa�;n�Y��w��jd�d8T5�Z��A��\����������W0/�B�g����� ���W3V��*�P��5�;� CQ���������w��� *ZLE���"��B_M�V�]%JCm겻�'�rY`=�ٶ<}��o��� �	��=�B��|��>�*�)��?eH���z�[�D�A�j����>�0D浌"ЩC�AKyq�<�(�!��飵��5Jn�}��s���Q�uoV��y���X����*�>7�BUD6�1OcQ,0X5�:vZ/#\-�i�I�	��"5�L�X��j�� L�cpx��Z]���~L���2������>J��Î��z�uU{u獔zKi;b�p��a=�X��1S�\;A�(��8�L�ģ��������?�]N��sT��h�L]�أ�s����3�d�5YGQ�[�>�0�:�����E���oI�1z?��q�E@�pi����>�Fu�/�ˌb��{�F)����%�ْV깎b�̓�]|��J M��0�I!�d:9�[��~�v������ �L��e����$����e��h� �A�V�%�N�W4�}0���ݫt�U��4��PW^���O)�Ô�|xyH|Y]�5�j�������������ŋl�	���I�㊇J��R���?�^2�sC�]��)i'!������!`�9�z�v��ȥ�=ӛS��eo�+����'�Q�+x��<��2�*֐JR��c�|�ymAL�F��OL�쓄n�J���z�gP�8V[�,���%�
��rV'*���YK�Q�a�n���t]���E��Q������6��K��z���A����q��k4���SP�i?�����/ �)\U�	�3�����QޏS���ǦR����8f�-G�	��J(��b���{y����L#	+�����Hy���f����/����97����u0��9�Qke�r�̰C�|X�c���U+!,$����O���Z��.!�C�k����^�9�]���H��&.�hmRG��2'�#�a@B����?���
&b����a�n�1�;
�,gM���a�-�8��5�[�z�
�'�0�Z�hU����Z�Su:i�>)�J?|�����*��.nbxnv+;~rc�K���B�HC'(]7|��!?�f#$�m�w]����fa<�T��'���Ft$�֕n�γuJ�<��K����e����P\}?�!a��O�6��1�,f��U<�'���5�ټ\-.A��p��8�U7��F��q�UMPH��H��v�/�ߟ�)�
4��X��	'���Z__��<o��h@x��D��
��*��	�H$g�B�i<q���WV��}
�y�Wʳ�Pgr��=�QH̍5�8G�=rM�@C	P�̃���"��߸��B-�\��}�G��n��G�Zgg`7���0?���%i�z-�4�ΎNܰʐ3��b*=�튜�KfG;�������Uܾ�^�.���L����;��޲�������-���I� o�	���i7%�!b� �����5$��ƪ<Z9�+xj���ק4�S����iJ��΢��/K��	b�9	�W��jʙ[FL�o��v�0�j�d��E�*%�1i)���Z�+�]FGU��> ��I�\���nfDj��/���U[�ZD��4W�(�E��XbVT#R:ש�(������@�i��W�\u�c�� ��/ (�YȞ��8�,{��Ǹ���Ȣ��Ls�P�ܤwc�q�cL�`���&�J( A����e���E�|��O}ͷ��U͝A�`���}�V����F���.p��/ux��=�B�[ӅE�"髤�ת�Y4i[�(��	N��qp�!$/��CQ^��%x���r��y&�}|� Y������x-U����" 3Z��5ܜ���� ��T���ƽ �CǏeA��c"X�|�?��m��p�;\��cF�3���	��,�N���G�v�E����Vz�R�z)J�y��lu�EtR�xg�N�q��`�܅�����q� ܀��p�Q�,�`*�Lsf��WX��m�B�B�~�:膗x���-p�Z4��J�S!���T���6��5��ǏiZ��H掏��I����T���8��9j��tx6h��mp�|U�5�#~@Z�~�:6�0P��&C|�!������w;�dz*������T�s���{�Ԅ�#pJ1���vv�66�U�bgJ5���Dѕ�Ƶ�͢3Ƈ���L�;}�N�1�����Y�=�����K�ƭ3��:�ZH�*"7>لd�������5Ftϥ^����'!�D���Uͮ�����7��b�u��IeS�vt �I��9�ި����m4���쓦��z,�=��
��T���d+9�kװ�� ׅ"�ЛɨbZ���V$��Ȋū�I&���T[Ώ�~j�95}�W��c���}�'K�keós7[�����?��I+��������t+�P����c�'����r��1����F�� �b���ۇ+*$�Ip��%�S
���3n��*���G�'���]�=�Ͳ���m�nIQc�+��/ ��4�n���x|gh����f`�iM��A>��t�"F&�,k��]�dHE��pc��*I a:�$� �q�����aa���$��4�e�Ӈ�9�H}(�`g��{E�ZA�M�l�:�M�͖��\nM]Z�%�n,0M�<���o1�����B���#�G�wA8\N+�V��փ�����Bq�WA�F脫S:�s�%�]�9��NBds�|6uO����E�mE2�5���3G�vƊ��g'@�|2��H�׼�`�����~��h�|����6}���O�?�z��z��_�)�L?���/p�V��4΃�Ӆґc�E�o/	*�i��Mz�%������/�|,eIP�R؜��t�+�
O��R�+~�|D�����?� ��OP;��>0�iOv��U	cm�[�7�����	G�"����õ�-n�3�Ae��-����˽�#�P� +ƋJ�1~z��|IK,����Z_�M�|�����bg'q��߅0 ���!p���F��.s �"�<L�OX���G��M�y�)5�ǳH/�d���Ɍ�@0Y�K�,&a[���+�b(���4;����y΢��X}����@��=����+���1�)��%�rh�S��x����B���+H͛����BU/�-�(�H���� ��s�� ��5��2�v�n��@!t	��뉆��#�/��b���Vb��X�:��mK��}j.��, ����\ו��[���3:��Vx.��-�ƍ�04b���q8�����Yؐ�6�ω�9��zo����f��y�@�c^s��35 Ls���T ��n�B��<r܉�g���5�}���җ����J�[���H4��|��!�����x���YR�����Ta�n `��=2s�f��Ӱ�x���n ���Y��댘��w�Isr�C
��	g퓯+e9�5���w\������;��V�ɂ�Q�;���wk�)|)@%����.Y4X3 0��T]����T�� �8�^�}(?�̥���d�b�Z/42U�!kl�'bƘp�F
W���}4���\�ӵbޘ2�K����
��N�|�I�7�E3�˫h��+0������!/����L3�9���{�!*ϼ2Z�Q.�kk]�rJ5ۖ�-���-��~H�x��|�`�T:�] �O�+Z.Nr^q�i���O��$���躙m�^)����3�TZ0���;c�Ҟ��ַ]���"K���3]��9�Rp��-"N�����Ճ�--m� 4�a�۫o
ϧ��4�nK#��*,�d%�4�e�q2E� ���\��y