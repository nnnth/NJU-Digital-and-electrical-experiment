��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������Z��B��Z����eS��D���Kg��
A�N�(�a��Q�n��U��N!8ߎ`ۼ<-:[�t1 �m��PN��߭J�]�V3E@m���nf��,rﲴ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��`��(ߛ�����@�N�3��R_�}���U2*��cj���X��݊�oi�ɂxh]{}�ʊ{o|>�,�Y��8������Wf����ʥo���v�O�)���(�Jh0��n9[�LOy�]�k�c U���T6�l}�Q����9q��B�B�8vU���aVP*�� �sC��7&~P3�+zl\U*t$���"�����dF���,�����%�I�0��]����p��������і�>��l�������;%���Q�:MG�yE�nW���}4�N�c��Z	Qd�[ӛ'�������W[�K̀G���<�R2o��0ڣFĠ��[���ao3w9�G^�ã"]?�`x��4-a�)X�*�A��_[�9e�fJ|XY����R��yz��%Gw��t�뾨U�龂Cc<��A��'�0���w-4�H��P(ŊeO�i�q�}���+���γ��6�MS��-�n�z��W�[1&�+�|��*��K	
����5�H�hK#���0�;��e�͸��	�ٝ|��� U�wP�������ٕ�����w�1�?*N��6�&Uf����u�r�T'��&��֍^�h��G��9��ܰZ�kVb�� Z�V��v���;����},��,�a�wB�@��8Y�G�)A�җ�NhH/����g��i��6�$��L��w��N ��+�M�s�x�}1��i�*��]�[��;Ȯ�@:�� %h�UO/�=A@w?���^d���r"UH�r��e��D-��� ja�v�oyO�K7�+�J-lN��l�יI$�w{�ܞD�`�I�I:)W-��>�Z���1ve�PZMQok"e7{�.1w'wz���j"1]�%]�rT�&[[��B��h����Xι.�w���7��3bg�8L嵸a�tbY��Pf��rGAs(p}.e󄭝_���� {M������R`EN��kO #��sRU���C��s�d!�O��Sѩ^oӐ8�tN�Y��	T���j���p���`q6f���ݶm���G�j�U{N��N���wĠt1��y��[I$K��c�՟BJ�z�qA��y,-�y�ck�������^�u,r�L_��x4����M5���[1eP3�g�[�3�>�����cA��6��^U�ϖqt�vUy�r�O+$"���g{z�#������7����ڣ�ľA�~[�5*e���E�|0���X}ɕ@�C�5|!Q̱��j�Uu�jqN��k��Z�r47��nl����+��9l��:@qg��Gp��h�����:�o�پ>��c�����X(��)�J��Q��y1�6���Q�.3v
���'��?�Q���};p~?>���,��w/�*�he'0�`A�U�?`b3,m�ti�y��-e� �c(�}6�N����_��ldD������U��VgCr1�;�;,u�:R�����%z�?�ތ�w'E���7���(�rI�"�P��MZ�>��+4P{"yG�������Æ�ul�O��9�:c�&��&�8�0��=�t����J�����;_��_����7�{p%�r�@j���S[��A�S	���>����uh%tǓ����g�~PB-tg�+-p[i6̲��_�SZg)�/m.p$�;r�_+|Շ�	ˆ�k �H�����Q�Q2�oÃ�� 	�!��0��Ǣh�n�*\��"Zۛ�v�yѝ~�����xk�<ՙ?G�V2��������}ܰ�Y��)+c���o2�T.p�d�kY1:՚�H�J������('��;�@���H���q	������Pg0 &�ә�Ku����>������:�g�D��>��_p3O��.\�-e�Xeg�&��UC�bo�-g�v����(,o�*	�Y�$�Va\[������z��hA�&��#xQg��]�7��k�<'��#�Q�O,�����48ܭEwS�q�~z(�m�G0��B�+�;�*�s�� �5�sr�ɳ�Gz��#҇�;��A���'7� Z<;�=E��lo�4e-]��}`��O"Yъ��,��&��	!2�J���ljD�N�v�y'v}p�$��+ߙ��ɝ?�G�k�xT���(-�<6F��)L�M��=�S��.wէ|����=��}�px�9W��M#0x|���])���ju������8��]R}r̐V�v���w��>�b�f@�U�Yh���oV!��	���򦢸��+Њ��b� 8�f�����C���b��Ţm��,�-��"�#o}������IJƩ���=��M'����ީ��t�x���b��ۈj
,��=�_�l�|n����{�y�v�WAB�d.dzH��D꺄�1�up�7�a<��cr`���FC,ל;�2�9�z����NQ؊�-����d�j,f�TlP��&)q$��(�q��6�U�z�[X2DT��|7v���7�v:��q�W~E�+<��Z�|}���?B24�:�|g3��k�/(%�����d>�5���Gk谉 ����X~�����)	EWСnz��O��RN�P_Ȕ��p>4֋ؚ�����~�A<+p�Y�QE�Y�����&q����	��S�R�6Z6sG$#�
}��W�`<7�q�)� ��Tu
m8E��x{��+c*��4 �Ƥ�q��$7�|�/0�����*_���
�#��~�_�'BT���1ɝ��}��8�X(�w�b����� 6n�֘�îP�b0mO�n]�5F��X�1*�5����������W�"����5,?��D(A/nЖ���3�24>V�),�y��v� v��݀*�R(�1DZ�����Ǵ�-���x��� �ؠP���~���m-V����8v"g� �?��\E��x��8#��w��Qz}s/��0�í��=����Wzܑ;���fÐ�#A�J�?:V����Yng��g�'�֫�0-�¾�3v3�@�a��*�j�׋�~͘c�ɶ����|
ջ����2?�Ȗg_'���1f�*;��>��4zTU��QloB��Lwda>RK��ـ٫�O7��=-TA�<&�����<7��R'�#�"ם[�G�d��5���|�"^^1CW6��~�f�?sNѹ�H��`S��X��&`����m=Sg����mOk=�dg��
���;��z!K����!_Үޗ�qh�c����_Æ.p
��X�uJ�Ēb7�}��uQы����n�j�a�F>��Ʋ,X���j�haT�4��,����*8qZ�qv�;�*�ե����`V�N���7 ܝ&D�f��6������r~xK�}��ȗ���ڧ:���:|�Jt$�d�r~�9�yb[/㋕,�Y�G����$�2�����=�Ѱ| h�o�y8'�����b�)�7�<3Y��=AvQ��{��EY�_3��� �BY�ŎT�E�,۰p���$I��j�V{{������y�.���q�G��\�u�~">�p&&͊�S�c�ۘ���\�{���)�t5���T�<���=`��9�2t%�Ҏ	3R1F�;�)~x�}|��/s����g�u7򗠤�U#������]�	����ʺ�F�"T<t"�;b�^��P̠z�{���èh6Z��z���E`*�T��ݵ��	s��&G�_��N�g?M+\4��V��%�+�r�rM��! @ܚ'p��j��dpn���
�#</l{ �����Yp���Z�Z��Q@�!�OrC;%A4�2f���ʣ+�.�ɽ	+&G�vP�pb�]TioRz:��U4La}�jH8��՘���7�f)��,$[�9�r��v`�g�+��z3瞀1���f�r��rԤaΫ�۵鏟��c�	{X�K���l����o?���1z��r+In!(EE|���57I����%�j�U�m�q�<Q��al�EY��0�ը���e�|l�ڨu�Pj���0��&�C�m(k"��T>����{ e�Ta�@%Q��k�͓%�y�0��5`�ko<� �_Ii�/NU��	u��G������AP3�x��-� �o4t&��OK��[[��m���G�ۘ	1�9sd�7t�:���D($l�f���#y�(�>oj��s;�oڴ���˗*YZ&�����3R��q�ht��r�gCE��A[5�g�˱ 1�d�Vm��\��xK.�����W�\�����LRѫ�����*I�Mv_��1Ea��8梩�3{n�x5��>t��RR���3���l����~L�u�b����if�
�
���^��������͢��4���~p�������=�w���08����`4�8QC��y���̅���uϑ<<|�-J�Ԩnt!Q���an�$/1De�(�|��Ņ�]�B�;E/�-+�I��YҐ��-Bx.Z�h��zюh+i}��m ѽ�����j���v�����sm��Mۯ{bZc՗-d�
丧���V]('���>_���2�JO����s������y�\���K�+u�SR��-��诮��2��Oh���XR�\4a�S�WOLP�m)��.=N�\˚`۰/H�A��(u��W�W�#]^Ї*}j5N�/<�aN��O?��ռ<X2|�Ea#s�Ʌ�ώ`�3;H�po.����K��3��~��"C!��!��Q����R�j�;���̆2�g�(�;���Z|b���������@u��>��_��f#S]���Z�"�r�$e
�V���O�M��8�R����~���l�}
�I&��l�M"#eaK�N�,Xmp�1��W@�(����%_�0�[ha$A���Kx����������x�0�nW�'�v��Iv�TȳF�\%~~�@�n�;H��ì`]���� 6� !�&4��"i�& �ʙ�H
��'2״�XXR����h�Q���=����3hpSg.V��2�ϯh6��}�0�+&4i��@�aϿ��@F��*���=��6f�,��?��{c�5v�1}	k$3�QY�����d�M�;3��]@��f��N�����}��GN���f�%��ܳ�!6٪�q�&��0h9���]^a{���eO���vGTu!�qs��O6����%hY�~B���+V��4p+�Z	O���E�f�*���h|8L�D_�1���*�r,�uޢ�S��/��m��{���ZE.���� ��[~��!j׻a�$�9/�`�e��V��3iƂ��bJ��Lm:�7�j��V�&��G|є��3�ỡX���G�j?{�pz�Hw�*�%��8����[7")��W{�]����}�o�Ծ {:�0���Rٓ���B�^ܑ�>3�6EF"�GS�Q�b �s� �_�����n�`��ly��O��C���3�O�]�-�h��EE�#NpB}��ݵ���]� a�VD>Vǐ���v	O�%t�-U�t	�!h�S&ɌN� @�@�0/w�t!B��y�I&�}�=w�%l���k�86����H�i-���#64u��^Sh�$|OwR ؗ�y$h  Li��D'iu��6���+y an��C����s2ؾ��q�3�d�^2��iK)�*��y�X�P� �[D�t磷לq3�MN��:__�l�͘��L��K3�'�N>;͚#���Da̒�כ*f���h�WRm`)߻)ZN�FOk>�yg�l�\ŭ����e�	V�L3���@!��6$��'��=Aa	'����¹<�c���1�ʺa��2>��/��ΓC��	�,��TI9W���z*!EMf�"d�)lE)�$X�s��^`G�go�i#ÇQ2>�VUA�<��_�C9�MS"X=���R��V�B�5�w��ʷ�bK���$o��rG�-����x��"�"��pC&:�st�Xao���2l��n}��_ ^�ݨ/��/q�g����J�!�OFµ�s�w͘���F�=I���X�ѡ�]W%|8�?$��0�9'������Y��˗��H�Rӎ�P�w���\l	�m����/�����d&]6"�k��<.7P�:�м�~9�H��g��Tg�<�������b�O5$q�ѝ�u*�J�J��[ɡ�+�Ϡs�4Z��G��["D�2A���!���&�������y��
�%��ds�ui�>i,����o�\�}�UR����6bT�<��M�X���U �,_����DODq��;4�tL�FA8��eyx�	/��1�đW-<��fP��6�Ժ�d�ݐP��)Z���t�c�g@9۳p��9�>�)% &���R��������CC�vy�0��rG�Sm����(�0u��,k ��՝�Ռ�'��_�}�❈�������.�ҬC��Væ�;9@{�-�L�"KRj�ȳtmZ�� {�č���m9B��= vK�z��q�K!�>�?T���*u���;�}����G�o㡫���K~�$Swf�Cy�T��0�^u�:!�B�q�,�t_|2��]�vy�w��¾w����3��V�!�ڑ���d�3o�8� �p�a�g�UB]�D/S�距By~��r	H�����y*�k��a�3���.Ž�&�V��$��'`3 �[wS0ʓ���a��{8�qi��e5��w*+7�A�<Pw����㘎��Y`��6A�;���*�QCf$~ɹG�"��#B��y�����Z���z�W�
UXm�Q��P�0��r����E��*���h�˝��xëR��<^�p�gH�V��ѯ�T5'y1"��q���s����.��S[����'r$��|��,̾{-М&E�ND�!7�o���ak7,0���~�B���AEiQ��8�E̕mY<�c��;�P����$���*	�>�º�����A[R���/�q��P/z�ˢ&p�!�}x-�Qp�6Ⓚ�n]��k!͉]�Ҽ*�P�3/}���>-�����l�`���@����kYj�n�eEE�".�,��m�Jv,~IF+K+	����N�.�\�}��Γ�YCa��_c�z�r9E���hp� A�X$���^F6�i�o=!��TJ�%���t��Zi+St����g�!t�Am���C���4|B4m/nN��>EI�������[������T����`�Pl�%�%�:����E�������]j��vBG�c�%[ W�"��w9��������Hv̼�O���ˣ:��S8~���Mŀ|��DɅ��aq���u |����pӞS`&XvǾ�4�TMH���K1s�)�F��Hs�ҧ'�Rm����x�P�����Y���2�.������2
p��yT�O@Ƴ-7��mZ�z���U��w#�bA��7>��� �`{�
�5b�x}}�g�σ��I�{�ib0�yIx%��p��gՏ�p1��5G�(�~�Z��=�QϑsaH��B��}���3?S!�[6�������2к ����g � rꨴ��F�ן�pfi�ney���,U�z���`\{<'H�{�����@��{h����EMA��UR/�ǻ�\�ײ#�~����/=W35(S�<̫C���L��7]�V����}�H�Ǐ�=fң[�|a�Y��t+� ��.6��Q1����__L��V+�֢�=wP5�6�N�D�������ի�>Bd�I'd�I��� ߦ�۩�Z�V�g5�ek��ג����R��9���dh>�*RbP7�Ծ�2(���V/v`��q�I�@u#��P���=�ѝ��ᱷ?!T_�7���Oc�+A$��
��қPr]W��#�������->����V��J5:�+R��W7fم@!Y.�nG��}�b� ���S�!(��
��VU��k=��f5q�8���OT�2q�v�ܢx-�@9�I��މ~�ˮ����n �V=�T�a��V�h�[h����])��(�;�n�d���jN��%V��x"ÜJ�P��TBq��훍��E���н�gU�����>/��Hͨ!�3����
9��ZĨo,?�J}K�z�i�IHv��΁p��	g����w�6�'/S]cxҁ-c �|���� ��0f0yp�>Զ(UR�NZ�7�c2�^Ǳ����\�i/Wg�9����8�}e'=ܬ�Ņ��~3F������IO,����'������"�:���i�A�	��D�������?�������;ε'��2f�O�ο�h<Ie�#w�v��M��*�/<9~��:�\K� ���_-N��Dab6���w� �\�(�=���A��(�ϗ7�;�ICon�(҇p�N���H�L�.�����lu?n�m$?{K����	�t�P?rn 1�بӕxؒ����;U��K!o�$"3xYQ�$�Ef���,�C���?^��4�2-�R��}����"���֎Z|
�J�*�1�������ء�L��P�9��XV�z��`����ɸ	��3��yO��W��pa�ri�O�TC�/�/�AnUbx��[V�Y*y<Z	�y:��|"+z�a?�����Ť�H%Z�(�|"*-��(/~�K�=���^)w�#�0�yg;
%ɿU���Z�;A:���A1��+5���Q�z/��|��̟Ŀ�����a $6�Ns'���|���<pcΓ���Sm1j��.����'��C}��'|ݍ��A�i{���]�(wڈ֛�@�C�W��f�O���a=�dh^�d�c�����.NUك�P�3��9R���Q�����"�({�KwKt�ٟ��
��#��~3�}�j�VJit���n���0��[!�.��K���X�V̼�k�D��(��z��!oH����xRI*�7\��)��i��+8$�0x�[$Z��!�؄*|�I��1�9e��z�}���5�!�-���Bw*�@��/���D�P�m=�[Qk4�mU*86�p� "Ι�,�,��K���aC�����V��v-� E�w[�C����H����A~�-�om�ad;#�n�g%*R�Ro���y(
c�E�%��(y*� M2������Ů7�D�,U dY7���ԑ�?A��������l���v��;�, ������̉��̍�L����\c<�Ѓi�q� ����lvA����;�X��\9��
��Z�6/�F���c~a�pX e{�T���F����NK �?�����*�0�T^���O�N��LZ?�?�C��U1��W��6�=�%R�Y�f�|E_:��m�.�]ꌠ;(��#���H��_�˲G��8m6o$xB���3�oz���G2��^�ͥqz�Ƞ׭���u��%�!��b�ۉ�Ϳf|�+=��3_7�y��F��������fK �9���� ��_HAr��~e����N� �[�/i("dc�U%�s�R�Q1D� ��D���AE��}X������~�c%���(��L��V��{H��s���s��&�(7r�8���wkn���.�i��*�\����ӻ(dS�0�׸�I�dH��.x	��Q�y�xt
I��x��4]�#x���c�V@��s���Y�,\��(Ntw��=q���ª�\;G-�*�2����Y3(
�S���JD��)䅳&/F��ԇl�C��7�����ڐ�<�;���Aӈ1o�K�,�x�%�g�3?�r���"�d�z��n!���Oɽ	�c�E�&��b�J=VR��Q�^�k�)�f�5��ޞ�S�Z��	B��a0�6< N.�t��@��a��6z�/�����3�
�?�a��ի�Y���'j�b�)��1�B�2oX��G�y�(-�Bg�'�Ou��@�#ő+�ckm"���/C���`n@Q*&�=���UB14�gm[��8l�u���ξʸ�ybA��;?=��+g�3������7���>��[�|M�n���jc��xƽFM�]W�#�Q��&_d�� �R9��6eR�Ľ�l�.��A�Kr��FE�ӮD�)�k���A���>B '~L+����O��g��B����c��%��m�l(��|"��s����Yވ�2qX��i�,�s(�b�~���'$�Ģ�����N�"����[����*`-q���gA���	�tgw\��L-��v��P��سw6M`15Ec��j_��n�<���b
mQKR�2ປJ�Cj(��M��}����n(�(	�+;���)�UB6=	8sT8��Κu
��g���'b���W����줠���4��s	w7y���p�3�X|5�2iS�b��5K~��/���#;�"������2�m�ޘ��w�H�@��{��� �ڜD������e��P�2aVF�lZ���}%�HJ^־�mC�e����L�k�o�4ycŏ!�'�k�>�	�زߐ#B�U��~���d��k�L�X��<_ו˓�fx|�?�;����=�b�%2�l�,nO�Jk�h�3�TТl4��<�ܱ�l-;���!���o��ى�o�{6����C��i�S�e��5;O������z�B�b�g�\/�Ț�eٷ��xmh��Ř��_Ov$�U�	����ܘm�U��� 
Ix�"�s����\?F��59�`w�w��r�rC�Fc���~����_�=�;�tU09�IQu�ZCx= �kBɈ:��ڵ�#K|Ӆ $���w��2u���Ha+�s{�'wn����  GD\D�ɽ�;��,���M�&��ҕg~23!�y(��V'��ކcmf�[^�#���_稠��%)��`��� O�7�*��](�I��^o�&����Q� ���`C�:�zr�,)���O������+F���rjٷY�+�T*�-��97�t��x��:2�H���,���үd�����A�-3l?�� ���dvԒ��{.y͏�1=�+��rX|���۟]Y�گ�u�q�o?1��X���"���s抸ߦ���=�J#��Npg�������Y;ˎ`,���^�<�6S�^�}���>jsٻw���k��kx��ȭ�(�����ӿKP���)~�wq�T���l�pAi-c94�?���
�aU�Z�o}��84!�9R�!�]��:..�?�B�i��ibʻ��ِc�`���s�”�>������2��2��ɺG��'ԅ��6�:���;���F1��94�=K�Z:upXpѦ<�.-L7�F;祒-c��]܉���$}�أ%�yn�ߞf/����Kڊg�m��Eh��.����k;�O��쾇�ӡ�p[R�-� ��צ���F�f�!���A��p�|$k�>*~�]f}�E]������|�%\d���� ?�]�w��U'B�u�]2_��z��D��&����� �x�\�6g�=���T�_y:-O�&EM��V��R�����Ϡ��І�:�@:����3���I�}f����q���'�YyX�_D"�������IPԞ*�x8�)9p��ܣ��M���%)�x{K`��[
���>Ic,�m�e�hOX��#�j��n�%�40��&ohpy�Fs�>�n6�яk�|V$���ti�{��R���k�i�]��Ta�5�ݬ@79#�q�Oo�d�� 1<	���/V�hk��Hc>�T�f��n���v��A�q�
E�&G�"�6�`Iu�{=8i��e�(�>�G��\7v4����4	ݬ�)C�|�����s�Â�I�=�}�i���Z6'�XM�E�&-{o5[��>���A��;�C�m�wf��JG)U+{����	Q)�pU���ɏ��I.?����p�����q���[{���|z��u�K�oN�w=i������߫3σ/��f�Bzt�K<�Nd�}kT�SX����@���_���q헆���"89ب~p����F,�1�l�[R@mx|An{{����ZT��B�r{L�9b�`;=��t �O�c��O��e�c�u[4~�r�s_����Q-�*V����3���͟�+�O��Q�ii�	�А�����]�⤙��D�c�A���ɂ����;�v��4>��"L�:@O  ��� �$�c�q�����[<`�rCc�iϪ��u��+�Z�g�bqM��G��h�ĩ��x���ޓP��ߎHOҤKr?��Y-��Ԋ�V���/�+ҡg�R���]�
�'	Jŭ���t���Š�B6#�+�S����/4ӊE�RY�%�p�ƵU&gzY����}����DWS�|s�f�퐖�W���H3���wH❒ow�잨c�����_�}e�a������Ω�h=�rg�]�~�d��`M��!C�������y������j��^y�<}�
�Ur@"wk~X�>�x�%��Tԗ�˶� ���h��{72�m�:"��d��][p�0��B7m6����7�u�
X��|������,��L[���T�&�K,'�|�<���w8�,�NAQۛ�z.�GߜFH�׿f�<��,Vx�ݑ NswQ2����δ���Ǳ8)��Ó�p�O쳎/�h�͇B��a��˼	g��!�����'�Z�������$�71}C��\�P��sj�.�Iѐ�2&ߒҘ�s���"��`�U��[(�����5G>��螕-:�4Q��|�.B+�]���<��t��k~*���*Xd�ۧ�7T}6�§��|��Z��|���E��h����g����g�-h�+E0]6P���Ta3t�
.�u��;t�q(x!e��fY~�j�uw9bޓ}� ��R>\�d��,U���)�(o�ڝ5ݸ�)Lw$p�Z���1�iL�����X�,��ǧ�P�*���
�3�RGz9g~�|d��6	�<B"��P��ĵ6�:}{������S6�H\&Y������R�a.+�P�*޵�+�Z��sm�P�$��)�`z�a�wD��5������MX�|�o���T�5���(�1滩��݉���԰^�X���Յ�9�S�C��y��k��=H��Vأ��31���z��B!�p��f��ǜx����vz�>b�<���eh �~c�ڒ���1��?	1�#�J���[M1�̎�����A��`f\����!T�f��CX9�(���9��Ϻ-	8����*��6aW�k$�X$Z�LVN���J2���59��IB5VL���"��0�rO����tS���v�V:��z�!�O���z?���}��(&W�y}�M��>�Q\Ւ���j��m���8��0ې	��� OpF�?����y��f���+.�*E�\�B���f�]��������/���Cz�lx�ft`]z�,p�9�J��{�������]�̔��!)2D̪8�z��6>{�/)��/�NõG�^N��8��(�b �p��B�/�uѮܡ0�6' �=����|u]���ܼ�ln,��5&�i'��[�2��%n�ý%!м�t���!Ŧ��� *a7`�}�'�.�~�+C�f��g�y�֦�+���^Yt/G��B��PヸB�YIs�1j�/k�;�o!y�݂����f���-��Cy0���{ש�1hS�K��^��T����ҵ�$qۿ/W�8��c���ɶ�óQ8��I���ap���{�T�r���0�P7�b�п�����kO�KB~�*c�-�:C��yj(���W,����:`�7�m��8%��ŁYbא;V�����|-�I��F���fS�v���ow�����8�?�|��kM]�YV�Q�M�|f� 
�k��A
z�{U��^r�95E�����0�p���I�怦�+}&��
�g���w� �^�Ό.V�f_l/�*�7�*�-R;���<�tc�W�oF*���ʏԪ/t���Ð��TX�����{#�����ϒJ�z�g�hI)`�E�_��L}R�tf,K����뷤D�&������+���g0��j��~�iy�h���`��b��s�1�����튘z�ŚJ��3�\o��䥐�Y����8Y��de�S���O��b&�gKg�O����q�O]EE�.0F�3$���~v�`-�5�8 U�������%zgK�A���% qݟ9����L�����	g���b���1-Y��$��?8�����_�މr04vh+fVB�b� ��EVa���=f�A9���b��L=�;֌�6�gQt��g�ۢj$���,�,xscX��Y���L�N^����Dj�UI2���0`���Sh��:`�W�q���'�\��,�N�`� �u��"F�T޳�VƠݚ�1lя'����R[ԯ��v^nb�������DW��&���;�Z����x;��Yi��شMyE��Ĭc���b<��~7��M�V	$C�%�1ߴM�輦��4>�f&�8�(j�L���R�b��f@���mވ�D�%Z���*	  c��}}r��`x�����CA��O���ZC�_�(�֮�npw���
�9�0u�w�4�vc#c.h
"-@�hU�id�*���F�ą�e��4��6V�6%�g@�O��c:C�z�ٓO�fe+EA�\~".��f�"V)֓���z}2���tD���F��9{�#�O��@EM�����/��a�q�əs���&DL}6��;�ݍ#���(?]*��~��;3�b�E�`�(��D�׌��?e=���(���O̴ ��=aws�C����������o�,3Ӵ��wd����=Ϙ�>�W����͗�I��ٳv��;M�ф���z�@3�K��R�n�����hvB�Q�/���B&�U�4F>�C�W�ipqS����*��1���4�L�?N�sl�a:E
�]3��Z��S�s!�H�͛�H<����d}�V�>��6�Ζ�,��l�<���F���e����3Ѭ��eS�[d����z��;�^�<�,���x$MfF${_>;F���i'����r�hӹ���	��md`�>S<8��3u�Q�
ְ�A��!���u�M�f}�9��S=x���E��]a�y��J���}%<R��@��m �a��PH��h���yV����S:`�|��������v�צj�d�`7	�#����gٺ^UַHz*°�Q&8�:,-�p� Q�J�=���_��.�Ω�g���À���V��$3F��a7�&[6Kr�)�``[:�{)�x,@¯W��A=2�ޚ��H�YN�PT�ʾع��\䴄�'i�#��U�V�Ek�w�����q�����S��w�|ݳC2��cdu��3s��b]�%]6����_�3P.Q��{�M!�((&{��y9�U�l/��tO��\
4�	2��*+�)��4��kr�v�Fؤ|�L.�Uh��]�!G��g�����H��^�ѤX*Jx�m��Bwt3BDZڔ�E"�uU����纙��x�%�r��L6��W3��(�EW4�:J�K�-a�H�쭃*�Z�:�:�%�P��ysJ��`��0 �h��<�k�h����l\���_��[�l��#�� �)Y[�� ��m�W�^�b(�;GlH�y(���ڽ��L�A����������Kh�$=�����7�U�^UkJ&��#IĎ��l=	>C`mM >q��N�2a�a��4o�N��S�خ>: �3����U&O��2Q*s��\R>~�m������JU��QJT�ģ���Қ�Xj���i���
�˒F]�N��25M;2%��wE����S�x*t� <�Owip}w�{Z�~�6<�*t�߆��h,��}��1��;��k������Q<��<��f	�u�������]���&�D���e$����k�*�J����)�ܼ_�lcNq?�Lq̔�
����m���6o�1��)$@$��$� C��ޠ�9���qt衝�V�*�hHD��[�g�;K���i��g4�<,�5U��X�oS���$�[:[]�^}�/MvijC��M�?i��%��W��+��NM�)T\VD,U��Y�߷"j:�4�X��g��^��ټ裠kձ���ޯ�I#{*��!��BG�'NIeϖ�,�+�4����Y��MWF0��8�Ha�����Tg�斥��9���r3��Ɣ���Vzx^�֍r ��TGbל��P�9W���Έ����ԣ��l���ѥ/�C*�:2y�yѸ+����l��/�ޜ�W$�:��mf!��9�����v��_g���\��e�:�rS�����Wc^J@(c�j!�>�
0���跉D4�&"��ʺ���_ ��s"�)����dB\��h)N!n=5A�֫q�L��F�[S���@@D����p��(��xЕ��P�M;�p��+����+]�;���E��.ʰ[a���vދ�>$�z��h�O}Ak�i�Lz���l���ںl�͘x��OHSP�y�K��}V�::�	���
�7�[�֒u��oĨ�O(fQ�������9���-�_1���p̬\�JK��˯�;0���>�!� 5���!��$�6�1��n�|,m�x<���A������@6��{�zT�J��'����w�R�S��8�P���ofP�F`�*�rV ��^! ��ؗ�� M��g��W�Ђ� ��V�L�Q�ء* �/9����x�z�/Q:�	��#�"����­�>H�?�3����]������p��S����i�Ab��pw�˅���S.WbG���&�	P��i-�J�׋���Z�Ͳ<����Vl���;X�|�� Yl���
��߆���r��QE%��(�,�G� ıfXL���O��!�##1|�j�-�}QBp��I�v-{��@��ͅ��:S.e0b����D�47�}������8���ba���V�h��~���$7`>��4�P�x^%T��$�+�S��V�BQ{�+j��w`�O���k� �������w�zZrs�q��7�S	Ͳg�^��5�Hw�u-��b�7N�7�чxaH�x����"7��_pV�h�p��4q�2������[����{=�O
��ֈy����]Qc��A�,�>f��ѫ%Cr��-� ���FJ$���>���ꞅ}ܻ_�&xJ<�Ņ�{����h�]�q��4p��dr�zy�菓�s�e�F���&C9��q��Exl�����O4ݬ��i5҉��M��P�Y"(��g���ivY ���2��֪�L��H�2Kf�W��N�.�q�6�ʷ��us�<�%vB(��%;y�>v]q�1��=�`�4`�G뛻�����F��G�G��%�5X�����}��p+���v�s�	(��O�󇄏�����I"
n7<s.q	D�`�aR���ް�� ���V\~��\�.hmх)Q�d�>Wt�?{��a�@�>?@ܧݑ\o�^���ɞ����$K�t��τ�R���3i%�韅�Ⱍ�ڢ��~����j��x*�f-E�P���_���>ev����]�_C���OD�+�?�Ɗ�
�]'���	���`o����r!��.�?-��PK��?E%����HJ�3)�T����vy�vĘ0&�2���~�>�zb��OI��XYys�ID�W���L�A|&X�[���>9Ǔh��+���Y�%��I�ڀ�N�P�$	���u�$��o�a��Z.l)i�a+�Mʽ����bE�ƽF�M�ୁ� ��;���v��S�ΨVJh��b�����g�@�+L��(am�v��l�{��D�~@��kDOо��fH��YB�O����w�ZLf�H���i�"�����W�k�C°"�w��{�d"<��� 2[H�r|u7r6�3��}��k�|�>�(�"����@�'�! �Q1��)�GTh(��Y�-�S5ffT	�hT��� ������#��H�.q�,��H{t�:����-�n�2��{Q�	ϗ����hO�n&!�9jv�9N�e�r���Y�+r@	@2���!�ct��^�{W�h��Mb�ڥQ-�jBZ�=	OD��1�WBC0��n6%����S���|�`a�����i!��eD}��k|t�~�"�S����M�8�����e�NS����S����i�z���6ƴ�6g��~�E�U�ˑ����r�ש1M�y�@�G�`�f4v�K�$�S�[��A��r=wP�.��ฑ�pV�M�3�=�cn��̜�(R�O=�A]Кf�ҩ����ۄk�U����I)���g�	���lmZ����;SX�i��DzϾK�'�@Y���0Z�� ���j �8���}�����C�L�.�ΞCgУt����a3�@���H��7K�V�s�� !�"�8��TZ��U�@�ŋQ�\�SR�� Vu��Y=�ӏT�f�_�Lf�<)���o���u,�048�	����{��P&�����S�� 3Q���X���Y4s>�su�3�@�Jd�|��e2�L�� {��?K��G��F�Fs��S�%�.�]kА�� �c����
u��j��Ŗ���0d��paXG$@j(�N���ZV<G�4$"�BtL\���9��<�8���1�X�Ff��L����B�Ad%P�}6��(<Z�o���.�ǾJ����7��r6�n;��Zܟs��E��N��qu1�p�ڠ�<YPԅ���R�)�}Iv�%��~��nd\��L6& !U6IȧZ~�-Y�l`ެ��j�oK.R	���z=&��T1�YQ����^�"�C輋C����	�B6����h�s�^�wǷ�v�qYI��L����/I��؛�r@��x���lmx�Q� zW�c}C�uN��\>:x���d��S�;��g���ܺ-U/����a��@���L�2JvMF>6"���/�=:=���f	ZY3;n�15 ����d)ʄ�:<M���iUt���ztV9O���}-����}� � sN�!���#]����-
��r*�,�
��)� �6��:�Y�J�W�!���->"3D^��=��5�h2�=Pe8���Ҍ�Z��m�����0�!rL��>�ɓ��a牂l,���#��D��0Gͱ�[p�Hk�CN��'I�� y'6�Sp�����4���6x.��	�v%n �����.����P�qݻ�ux�'N9������qpl:�	A2���y"ZS���uI��"�OL��������좺��ϹxA'� Gxl���e�F�3���&dT�.;����t�+i�$JN�4=j�'���ԕ3�E ����r�O�^j"fI�ێpͨ �v��ևV�Ļ#hL��k:�bMO���Z|�)WGEs)5c���E�vVA��f����۩��7>��KS��g*�����Td�fVYBb�{(#��O��VL�v��G,`�!���U �)��J�=T��:zW�	Y�R�uNJ���ZSqF͖�*?�Ct�
��y���HKV�jF�g��#y�jwfd�=�!A6�2b�Dx|;a�$�U�&ru�Z�t@���3�"�k�>�N�P�Ks�	��p[�Bw��܅��;�~��W�T���c~a�S+��M��n�am�C��������a�����RZ�;M��|ׅin��Vx�$	�Zz#��e���[a��#~g��;sh�V��]�a�x.f�a���'tP�g�M���Ó�,�}}"��{��&�����O ����0��U��UE�)Z|�����A��A=���A��Y���V�W�ђ�"�������9��^@�.��?qlL�R��m�@�+�\څ�e6r�m" K2�����1�šT,ƀ��t���I�4�y�a��ʁ����k3�\N����MP���b������F׼�m���!�����[jߺ<�R���ކ��b ��0� ��Zk���� �Y����њ�9��k1���|�F�|M�4pw�P�'�`X��/�zt���hT=p<�a��ScR;U�8�IA��C?��
�mԦ��JO��qd-�څ�p�0U��j�ZnU�{\�V����pe+�VQ�T��Y��;Ys��	���Ԡx�'��H^yϤ}�%�*/���q�p����bq�u�^Ё�_�@�p������|���p[,Ĳ��ړڈ�1�~P�F�^��KӊG�-��&����Vɟ�^�u<oRс�(x��#N�RY�`3P,T�(�[	�W����긟ίh~�#ߌ�ʇ��)�̉l?h�-ʅ'��ܔ�y�[#��&q�����6p@��M<CYl���,�K�п��4����$p�)22:�����
WMW��
���1�ګ�(���&�	Qʆ��]��{�o.�mղ����w�%P[`Dr�9 ��g ����
�J���a�msBj�A�g��Цx��	�a�䉻z��s`�g?�1��a��Ou=I\���7�Q���=x8�9K�k}�l�G�5G�M".
5Mf���{8���A�D����E%�5w\Rw!�If2������9�#&n��l��JnUJ0"�؛c
���W��iK(W�-?o�����g��d�����9I�e�"1�@�+���s�.���:�G0i�j~'ݣ��-����y��� �q���f���Z�^�W�Z�^����w���]�(��]�.�5otB�n�!�fպY�r�+ρ$ξz�]!z��ɔ��+���E*�8$�cIg���'1vsgw:�'�f )!���K���������%���]W�E ��ثS/X������,`��<�<V��7l��4�>��YMIgr���̶�q���dj��!�py�qi��6w������.uZY\M)���W�k->�@�Ĵ��gm���z���/}��9������}�z�ԪVd�t�,)��u `2y����{�d�w`�y��	}��<<&W���m	�^��E3j?�bJAwR���`�ɔ!m�^�w���{H�+���©1GC�r�L.��\��;q�cHFF8���m�M��EZ�p�*�w�d���o���қ̬�4s��q�l,����%_y�"ջ�pr����0�)�����p�8M��D���؜���k��s#ѧ�A��w0����[�����|���q�%Y���]b��Z�ATV���a�����(Ve|�U7�[I�;�b�z.�F���ܧ,L��(�j�r'�n=j�=�Y����5�b��܍Q�,cc�Om��������O=���L׼
��γ_�M��*.?6#9Dڑ������~lb�3�/�B��z���T΁�*�N�'�Ծ^�#m�l��
�P*,�m���=�c�oF;>��&7JGxn���/�x�x�U��p�I��ӌL�O�$������D<yGv.�0��"aXP�H�pz�j`9�N,��k[���=ofK6Mݡ��	�iV��mq����n� !18UD�K�Pȏv2����5	R&_賐�)T4��T��VY\��8�n���|�4��/��z��pR�Ӥ�V]��0wHp��n�Z�N�,��b�
 ��k5@�m؁�7�l[�)��������E��o�k�-�~��8@��I�ס_1��>������(�棽
zn��&�el?c���y\�G}t�@`|}�T�+\�
��H�c�B#��B ]C�+ �9.���%"��D���h^�8��^O�~"�wJ1�O��`��U�����YWT��'�
:�Eĕ�j'�
2�J�`
��'�Qr��N8�-Vl:	�!/��-t@�E}������Ҽ�3�sb"�~[���b�bE�\��aq�>(�@��k��ǥ�� '�o����B�,������Oi�u�ћ|3�rf�ɣ��2z��3��aO�����%M%.<0��i��+��O�a<d�w��w��LS��qƄQ�1w�N($%;U� ̙U��j����� ���b��+�}P����k	���5)�3�3k�Bt)g����UBі��6�j4Q1��{~2Y�|�7�Q�����鎇����iY�|�'P�MhV�xvh+����ɋ�����Sd-]Gغ�9��{�<�����qx�IG��M�����I���J}ܸ6��w��iBD������_̄5��N�g�ϯ1��3O��(��T�[L	��i��z .�O�X��@vP>ATo`C�t�S1�:�=7l�s3ʚ�'��"~g�P$۟�s#W� ��d�:D�]�̝�ϑ�?rja7z���7��;ѯ�p`��	�����B�r�c���p0�����d�詖���Q��'k�u)d*I�	`e@8��η�_��H�8O��y`\�{ա9w��8G!9@h68[|!8 uj�Z�(�cf,)��4@P2,ጒ�K<���3BH��n^��A��i)���@���,�x���[�۟��۔����[���d
i�C��~@�b܅5)��j0�����;y��6M-�Z-ǋg�Bȯ!��#l%�� �.y������
\@�H��t�B�f��9���F�����9{q�@6+n$��i]RWc�^��h�_�D� �ow{��ح%�U�^Z+��)׌�!���~g�#�?�lH9��l��!��,��Pr P,���KR%R�0�A7�Ebf�Ю��h /檵��(4O����Z�lβ�?Zl��|���6-׽E��ZB��)��O�3H��<�Zyح�CX�;��?�K���U���ojԗ���J�f�jdKt�:�������DSk6�Z�4��r+�F��J�<����ҽ������U4�yJ֮�g���Ys��sP	��3��R���dy~�u�L�v��ҭ
�����B��ƕq{���`�B��M��J(���)�J�A],�Wv��C�/\�[�]�4�gX��? 7H���$�p�(��}QS��Nf���-���w�vX)�A���U��~͙���z��;�з1� r�[)c�r�`5g�a���_ڢK"*l1O�lr�lU�����%|ܑ�)�"���6�������~@�B�m�E�3!�-�/��@��;%���D"
D��jz6|�ߐ�;
�cZ�0�����y]���D0Y]�#���($�C��R N�_�E��fG4ᛗ�-���� �ÿ4A�BQă�'�'�5�E�A�O�Ο��7�4X��d_���-u!��zu���ko��
�1�+��u�j%K���E��y�{�����*�'SB�ɽw�)+��o���5��a�/�q�Їq��E��ɹK��P���b�m<��-���ZC�/'\�eJ���W�p0��T?��M�.SunF�y�?��tbi	����q�/Β���p񼠨Ǒ(*]ʠd���&�N1��T�}�2{>̿,�7���M�,|��`wj�T��э?����o�FsX/	6￦��۳�\�p�]A�f�@�S="��[��.�7$��MҌq�� C/E�%�Qg�o~Β&�!\��6i�+B�w������PɌ��C�x�}�o �e^p\�ho�+�(����6= �0��d��`��^����%��Bq�rr��B�+0?��⥎��H��#���l\7M����w��#��K��[C�|�����s���Ҕ�=��>��jE�7����-~�}��:={���:&��Y_�ɩW��ɜ(�^�F]!�)�	��>�b���=_2�����������AD�k�x^�N+}��]&'	�/���㉮ �UO|�B���e8U��S���xsE���W�w����"�K�_+ �!�����F�L*�ز�X��+٣�d�m�wf�����C`Q@~N���߇��^�v�N����M�0[^{6ʺu�ba�o������C4�^�o�����ٝ�*��$>섵�%���m�د�/�������0�Iޚj5Xlڳ�,B���	��)O��W m�ޖ�f0�sHz'vV�O�|A���J~���V7+ӡ������X?C��=�J��p�-�i�sj:T׻��כ�9�hT�(��T��JkUB��Lȁ�r#��Þv'0$��=��Q$�|�!)��P�J�e�>%΃"��<"]�-���G0���cJ�tQ<C��./7�q��޻�tq�l>y�l���CL+i��$��GaF���P�G��/n��j���a]#UB�X2�v}�,�T�
6��6z�,+���{���"���~�1�zp9.���Z��vʅ�26`{��ץeb�������2��Wȣ�����B'Sd\��NΡpc:b�c3X���{8��Q�T������W�6Ad2����s*-)����l������:D���m{�Z���,ھhN�2� ��\���N����s]$��b���.�Y� ȩ�4���U%�,o�)�tf'��.EV����
I���,'.�x�I]�@�z�t?7�8�,u�(uPK�A�`�D�އ�Ɂ컪�)^��T{� N��%�L����l�A�V��x4!���$��6��ks	���p#.b�5ImO��p���ZN�R���B�Y)ǃs?��@1V$�Ό`د=�K�&ғ����o��2;ݓ�����z�[��FWH  ��+��2_�(�]�L97�T߾�9��^��X�>�2�L�6a���D��.	R�G�K%�e�Ck��mB+>9>�ЁAE��k�$m�u��]�b�ׯ��.I���Z�*�<�v�� U�V�a�Uae)@�ގ��1��^��ċ ���Zq�#Ұ�G���N���:Z�^W$�UxaN�<#<��ŝՙ6��X��72��΁�E"�@����*P�����a��?�3�@�o˚яW�`��p�F�.�2�cy�(�O������6iG�G��ق�L�/)�_|����ew.N�\�í�%�bn,����%}�$��r�Dž_�R�|Q��<��_�E�5{$��;�6��-9\��~���uӨq��MWy�-�:���A�.�6 hx�!K+P��������r����Ąu�����s��>2
lA!c�_T��V�����Iy6�&�WDa��V6%#���EC�����'x�I���*��'e��kYC�Y߮�B�L{���_j�bG.}4�+n��-@ޅ��W�f�e�w4�/ԏ#|,�By�R���w����/�
�u@
��Bv��8<kd���o9����ĺ%��h�I&��W�W:�8�t�C��%i�w�z��f"v�7Gb3�8��`��Y'��h^1s(H��:d�\�_h��L��hq%��ߌ�DmZ�r�o�G?i�v.P��\|�o�*K�������Ӊ.2lp*W����K����|r���>+��w6�k�t$r�� ��u��#�^䘍Lh�B��$�ҀH^"`?E����p}%2�����@�̵���u�I�������}!���ݴ�5s�O���}�C}.��};�ot��j�RB�x�[�(y�ݙ�~E���D�J��3��^KS���<��P���=��صm�8՗�4_��(l��z��`VT�2g
����(s�R�eeGf	�,��C�%,�yئ��܈T�eF|h�>��T�L�l`��4sT�t�|�~'U`���!�0w�"�a��8C��b.2d�$a���A4cKL���i`�c־�(8,e1Tl��;�4`��+ˀ:0z:(�q?��O����$���^g�>H��6N�����,��ˋ�-���5P�N5F��u0�/BL�����Q��&nfPR�1�}��� 1�YH�?W�U��g�R��h]�y�A��VW2����K�|�cl誯��zN�m?do��/���a�����z�un$��ꋀO�v.sS�5E��Z�������_�Q�����F\����0m�[ԓ�A�FgZ�yY�&]eArF�"�[Ϭ*����|_^YʘgNA���o�_´g�[k�x�Ο�w�¡��GC��[ƀ_�a�̚;��p��C��m�nC�L`���JM.��6�+o�E�aҽ+Eׂ��sŔk0�Cs�[#�{X��Rq��r]�����m��9��2oZ����҇LN�S5�`^�!�m�N-5���`c�R\�H:l��ԍA�pd[���A��	�s qe��]8i܄9X��I�ꊫ�+�%@4�{G:���1��*��4����8�,i~&�9R��(������%p|5� Ŀ�����C��vvӤ5IDp)t�Ԇa��r�y��39���q�z�mg����B�M����	��B'�Fo�Y%��R�E%^}�����!��cz��c1^���m\O�����?Y>4�B������W��˲t�5Ѩ�2D�r�"�K
<W���-�	��/g��n��s�ɣ�|V��"61CRPy��A��_�%*|+/����/��|f���x�(N�K�ږ����1���O��J� r@N؆� ���!��Tw.�0B �圻G-������'o[C�x$�y`2#W<A����|g5K��iuULzc��¨����s�&��m���!���Z����3a�m��ש9(L
u�޼~��1�F��Kxn�u����!�(bN�n��r����7@қ��r �١�-� Vul�`L�@�x8hb:pnȳ����O�+$�������f��{;����b�����g��\��5���a ��`݀�Igݱ���%�ܱ�x/�q`0��s	v����Kl@/���'e�=���cKg��(��.�,D������,ѷ�n���G���E)�}/�>ܱW$��/V7�ܐ�I���d�DLJ��Wg�8�nR[�����ċ�:���pL
n$cԿ��@C�U��P+��Z bLN�*>k��ۜӂ�{6;�qu�\ �Ŀ$)���l;�$l�%4	���.^ɓߪ��)Z-Sg:���^jG^��'p�M�NW�S��g[�pA�:�V(�&�x�h�K!IY4�(���TfD���ƵC�ݹ�;��g�)�6�a����+���I9R6��!,�.��T������~=H��Q'�{p�
	�P��I�5��f>�[�rw�Oӭ��omV
�P5�ټ��O���.<`��l�y�<@_;��P�#U��:������"��N�$�sE�)S�y$%Y9�
A�*tV�t���oô[6~8���X��0�:F=��6'$ZG#��T`����e��Z���y>���h;7�^ϳ�g���q��)����[x�2���G�N]��s�>Xw\���ܔ٨A�yջ�qV�Z�Dz1u.��157L��'(s�5Sw���S� ���i����JDt�_#b�8!��w�>]�N�W&{9�
�NK7�-��b�!)X��H7��=n5 m�sºv�/�����X?)���A��ƙ��:�>=�9+R����3hd,�{.Ld�H��p�d�
K��NN�޶r��v�Ֆ��
�n�}s"�O"���v���Ȥ՞7�(OU�0�c����y�c�)�s�XTKiɇ�Ie��֤��~��_H3~�ہ�0����5��]F�ȯ�`"��5�S�Cq�	`�����3[��:�AF�� p�q]�&�sb5���)��nP��_���B��r7J���[q��$�D�ݣ4�&�>�@�_��V��b�Jp����{eRH;�\@ g'Y��@Cq���J�?���v�T����P�^.$r�)��P��:pd!����]�2P���}fi�f;���eۓ$#���8c���Q�S��>ZW�/��ghW��=�_q&���m/����T;\KvD����^�������2Yo��]q|�άz ���-�����Q{.�����vH5�@��qC:Ε�#�g���-M�\���G����N�B�Ŷ`���* ��8&g�4�����\��Rr����f�W6kPhơ (G��qvG���X�a��.�-|�U�y��'��Ż���L�fS#̺�$��Z�����O���{{� '}kr������5����R?4�wn=��兖zbP�P�IH�^A��Ϸ}����4��
/ʤ�0��܉j��@+"s�u0�r}��?njUi��by�NѸqsN�T�������tt��S�ؾ�5�^�?�1FO6�U��F�d��"B�����	|0='�*�	"��e�~3 �~;���dFwϜ��K��-��W��������lF�MN��cM��G� �C�Pm�����s�W5y�����}�:Lzr�X������^�O���������!w:�L�ǩ�B�%!A#�ҡ����E'���rW�oK��ZK�����Ⱦ��; ��T�9z��3DVJk~za�Ie��$� ާZ��*�h��^�� JV���؀B+;J�P�*x�BKGe�P��?*�5�4G�g�AA��LW��L�׌"hr]O`4���noگ����,���v�.����ZRz���/�.��ϬI����4n�lk}��s��P�(l���5f+(x�cy{l�ZJ[��\���*3�].�*j;~:s:��� }^���Sy��YB8k����W�Kj�4E��[%3��${\���DL���j�J�u���r��4�<�K�;�ʔ�0�у�;_r`���M��e1�8��ń��rƾ�����y��C�^�X���2��5�2�=xrLvkܻ-g]�g)6�w�$-N/�j���<Z�N������X�a�j��݃X�$��H�O6���0�F�_����ԧ�S}dہM
'qW��9�j'�y>W�)����7��KXי.��jd0a�r�Ls��^ph٪�X�ŵ[��= �G�̙
`R��su3��=ϋ3��D��n���J?�O���bv�� =�Je���/����=��Y��rsJYF0�ͣ&��M�Kg�˭N2��X�&���u��g �E�� �:�D���X|U]����Piw��
��8Cg�UWţoW@@��P���W��>�%A�mtg�p�R���Z�a�r##i�hG����=�H�nH�4�b��%���6���V��\i2�>g��	�����Ӡܾ�ɺp�y��n�:��]`���a�v�0���ؿ-��|� �����-�6h�f��/�����1�fs؁ó��I;w+���[@����ADa������z�ۥ� ����%J4�ճ��� ���w�AT��<n&��UCu�E��n��?����Ne;�;r�! u�.�W�#��Bq�fl��:�	��"�>͚�������
�=S��p � �������{ǮNc��x��o��{��C�y�ٔ��mE)��ݢ&�P~�y���[�/M�-�ʳ֟���v�ALh�h���'�zx�����[� ��S�p]��{��L��Lr=r�#�Q��y��rJ�[Z�O%Y��J��Zݸv/���u+�j�:�V����9'%5dkq!a��_�pae�~t}w"m\��� �
T4�������	���-4��	�u�\g��`m��Ki������զ/��t��&����[�P�G���sLM��0��#e�U�GJ�Z�]} �1�:��KG���CM�Y�g3,�.YzͤU`Ӌhu�������&*  ��z�5�����|U�e�陁�g��0��+[:�IY'2N���;%��=��:���%b���A��#�`�vt����-�M��%�$�p�D*Ѭ�[�����@ξ�4�@��rFN���&{�CK�oD�Cu��43�D�v�Y_6���壜/��u����s���_|=����R��`T�z�^����}]HW(���`1O�]9U]��-��]d@<�7�l�դ:�73�k�TƑ��z����9�6�I�i:|�����Wu�i�uF9M���/�j�B�Uҵ~�z�)C��[��G7��nI�����Hz#���0C��
������tV���������,4��v7��Y����<!Z�-s"����o`e�������\9U�g��v����~����� i
%!�X�;u�*0��oCD�2��Le �O�<������Vݶ9�v���њ���aE�HQ�T����wOE]d��_]Y�{��c���/��fvH~]����-ƌHT5�"O����������q^@zX��X�'��\�	:#ƚb��}���b���)!D_���p]f_�`w &·8Y:�����E������2J�(g����G���%��P�:���a�'L��[�������T����1[r'���`��@�K"ˢt��g^$)`ʡ�W�+)9��A����s��ʼ�ѻ+k,����f\�����$�́)�������ʯ�x"p+�<z��Zb�r���$t�#gIk������7,�����d��~A��}���$��BÈ({�"��.EBg�匲����:~�4"�B�S�J.}��S��M��Fc�Om���[��5�9Z\��������~�;h�/��C"H�26�n�);�����|�Q2���zt*n2�`*�"�|��pÑ�����TP�(%���H4���o�殺��7�f��@���ӅL
� ��e{Ś<mǧ+v�G�"5���p��/0���'�W�e�\a��{@����� ��ة}C��V���K�d^�����n�?�%'����\8~��afϕK&���Ri�J?+�2]n$V*�
=lևȥ�>ש5b�<��7���pU����Ӭ�i���:��.Vxp&[����"h�L0z��K�}�?�;z��vq��t/�C.�T��&�����(��f��t��"�̌)����*x\/(�W	u�l8!�.ٸ3T��L-y�2�C"R�tgz�#F�ȞΚ�)����n$���ʉ���v�y�d_��τ5oX�)�A�?�h_����7)&���N�����DQ��Z�&�3�]p�,����Y5�]�"����W���Պ��f���E�6@1�`�	�D|���1;j���\�(�m�<���Z5�y�.�g�g�r97�s���i�m��UC��J�pKj*��\�V����C���Ys�ˌ��<���j �L�\�kp\l�
�ܦ
*lM��>}����&>5�f�k������h�j�I��&�昌y�s����0�j/wZ'�!Zx����D�����C{QS� +G%~�d�V�B�5�5Ye���~�۠�i����ĺ`��]�9�O��Vބ�MY����L�,N�>̟�R���z_������-]�<�@� S>	Z�W8$�[!�H��:@�Z��+�2�봓L���9�`m�k:^_�(�+�Nc;}An+J�� �id3�T�����t��>�ig_6`��p�$b�~,k�����u�M �Y���H`s56c�;�x���
U��_�m�{����3I<`qOTgv(����u��2��n8�4 /;[��8m�������+?AZ)���G����ZM�z��Da�|�06���Q�����A5�Y�[���� �翂�Y��O��8(���_�-�% ���z�-�Y?Ŋ�뽵Ȍ��a�Q�z�:?�Ϻ����'@�(v2���(���SvӤ�81�O`���tr�b�k��+���>:����4v����g2.;��x�I�O��U�|$`T�2\ bS�Z$J��ף*�xx3�~#��5u�o��o��ner�zW�𹤛'C����Q� �pn���<�_Y'�ӈ9w@��B����B��[��l2}�S&C����Kw2s19�w�R�*��#�W.�-
����0�N�-+��(���ЎҞ.ײ�q�����y}#��qR��2�����zRu>����ـu��~�u��<>P��������U� N�H���%ٴ�WA��K��/�/�� �3�dݠ(�5�^4	i�W����"��y|��ȵՓ*Uz��i)A������c�� �q�Wwz��#�0J��1_�Y��c��w�9�qMF�Sk��0K@��*��?_��%̺ۃ�v1 տ��đ%O���{����E�����h�����؝q�]�F�>24��o�H���Ӄ��j|���1�z�A�2ZV�a�d�%��X��k���^h��S8y��M�SnQ.GeU5�xX��8�qD��i\�4�R���7�!$'��h��i�э�I~H���*p�yڦ�X�,�(�$ �?�p�����\��6-����� �(�W�`�1$�4�0��&8���cI�_4��f`m�X��|
_E|�F1Z{}#��[���j���P�v%�t_���\n�sm�����̾����c�p�),���Ѧ��_� }s�W����ڎnO�1�DͼlA�q���D^����mA8�~�*�d�W��c$��M�~XYΪ�Z5����gҮ�獗��"�9Zd n�N�-oJ�Ӗ�h�B<!����V7(��ڳ��p�\�8�{'�b�^ �
w_I&��
�L=�+Nʕm�@�/�g���|���,.����l��ʹKbX��>e���s��o������A��>Kp��[īi�yzS ]�cI�>nX�x�rG�3�N�����f����?�]Y9#dCԧBw�/�@�C��%�����:'	�)ߪ���D��01ڞb_�X�⩀Zn;��*�N���O5�,�V�����'�����ۋ�낪�s����嬁N ����������L�Ui��l�`�� �^<�����������������j{�_���^���Ҟ�ܞ1Ҫ�k��V����؟��GK�G ��u��Jj|K�t͑J4Q�&ż��d8C#401�
ިT9՚.���]�qsl.��F�b&/�ݠ�o�eQV�>�1�K@�F�Y-�RL��4�_e,�0��5hpOx�����˔���!,���{k���̩X�	T�-��x����]Y?�
��@�~y�'�Xޗ���n���N7�L+���L=DP��.B}�Ds.�����0a�WH�Q�4
X�O�ٌ�m39��*���;{?FAA&�A�W��ptd�|M"����Y}�#��UB�G��2QSP~�P����5#��p�Љ�]�Nt_�5�y�� ��Q�c ��~�R��������[A�GV�����,O���g��V��}2�#�2�MX�I��p�(����*��x��U$�i��uQ� $O�n��iY9��4pu���Jw�~�c� i�!�ʒ�<���>���7�Y�є�]��D���E%�U��wX8�����N�̥���9)�����Ĩ ?���ٙi)�d�����?� V7��hd�}yҏ���NQQH՘'X��W�<�����>����AyV��܀�}�*q/g``	�6i.�(�2�.{�#�i�R�O;�?���-�,0F�B�;���
�<��m�:9Q[���>�Ցj��F�W�o��D�i���sl����f�?_���$B��gE�;��'�rl�9�0t�?���'	��h�Ś�6��T�����	 ��扳�`�KF�֌�m\h������39E��k|��f׶i��{����`��Gk�ɿ4�U�<��s;vV<ض�S4.�=Z��V�;���6�v�|��k@WU��L�(U�Z��[�zO�4"U�E�ߌ,RF0Z�5X瑣�yؔ�{'>|n&@��C�oYb��@����6^VI�j��#��3jų'�U�Q�x	CN�E��:C�&�����"�	�l���+�5�<Bŀ��v�^��|��L��?��h i�#e��å�áy��4����Ⱦ�#�K}(�+�B�q�n��# n��7�o�i7ƙ�0�E��3��x������?�za@��ZW��ڇ�/Lj)ű���P�LG��^v�����P��G�ٌx����M;�t���-�Ұ��( o�H��z-���w�����fߟ�#U��i���$���{��j�i�P�@�4��pYs/��V��D1FҘL���C&M4�a�kc�F�-����*��θ.�E�6M!���A>U;�c��^8������=���kBϫ��%R�����
X#��p_�Y��P�U&�Q7>�ft�WMn�XbD�&&B`>�U��V��ᾦ��:���B#�����f�����-���h�� vM7�0�!��K�N�p���!f�A-鐨�si�sڠߣF���B���*EP�0�Z��< ���[{ҖhڴU*�D��{�uF�&��Kj��7`V�w��%A-�-��A����5����3"�A�+��827vKDL�Cd��P«U���̸����)�O��V�Bf�]�=�g�1y-�i��Ƭ̈���Yv�To�j��̖~�.\�`(���9�X���p8I��H5�����Ke��y-�U�����=)�dHЎ�D���z�נ����r�z��s�0#;H�$PHm�f.��6��Y��Z�+���<�q7��-q`O-~\g-���i*>#ES���P��n�@��=�UZ%�� b��p	/���Gx�tG��7O��c�<-����a��FSM�Y��ͼ���=[����Gf���w�W�-Ej�r�{�@�S�>���A�{{Ǜ���}?��	p�Хxp$K�% RQ��K_F�o��(n1������l�֢<���k@���s��RWo�v���9r�
/�#ޙ�Yzz̬2� V���b����t��A�銗��cg�H�2����0r�)��������5�����#P���q�t"���NX�\�±~1=����{%~���YP�'ί:����l Y��9�j��U�0Ĩ7��'�n �w�I>�s�XU��1�Bt��0ls�ٻ�02"j�B�v2q{w"���9�|9R\z�c=Ē(O-e�&��Jz5N�~�z��Ϡ����t�;��Ds��,��Ɩ�6�x'6�MTo��Lp:r��4]gg&{�����#;�s,d��޶�Kwː�8�Q�uw���BS#�����p�b�������m<�dF�_JJ��8��NS0���*%�7!�����x�=�Μ���p���4, k��!���k;�MFX�<��}s��2#����N��>����R؃I���4y�����e�����͐��SH�����S+�{�n��UQ�
�@ا�y���-�;Ź6�c�٤ 7d�5u����u+k/�����AU����Ų��K���K�>�ȦMPe�V/�/����X������6�kAn��KU6q*�#d@�����K�Rs�5��"��.��ÀX�	��ޱ36���_��[Jך��>�����ZG�7���`.-�gA�4�]oz`E�d�o���\�B��0�p�L7B0������������wKz�"&j��_"�}�6�>?�8h�n�Vf��4Wާ7��{|5��^�����Re������m������$6���cX�HX�A��������(���q��{�{�%I����f�%��|����ǄP7����1d[
�W��'>z������+���]d��c�1�9���a��k=�qp��wI`p&c	U)��ym�e4�=C�37ǣ�7�o���4lQ��#^>�L�%�^Z,35�=�DG���3Ƚ:j�ˤ�vL��Ds˴�q\�E�ź
v�dғE{z��_2r���xYS�{ $��e�6�f����d#jժ��V{5z�d�AY� c���{]���Ml�t�ɠ��n�]�8�zb�nk����'������������^j�q���5K� ,+�
u�fL#�\����2'�9ۤ��w�0���_���,�au�6�r�� C��uWc�V�
�'��=Z5/���H��:�#�4�� �]V�'�^2���k�l�	ڰc�=c	���W��j_�g���X�K��X�*{���ߟݲ���P3�@��gMſ��)�@�S�PT�	gX���k���KG̩�p�{\=�`k�q�;�#���^�����i���	�!��i˻l��n�yY����y/��:�I�ȉ|J�jѨR��4���h6'�i�.n5���$Z�{�EpY�����h�$��5,>��&�������#�r?�X���FU����Ő98�UU
���z^ƴlL��Q|�8~~�<D��	9$0r^�)[�ݤ��L�	0f���&3d������ -���7���݌
4�ע��b,v���!�xK)te���[��ǀ��aҙ������<4���[j���>���_~�C7��� 2�A�(�z��>D@_@Y����raZ���o+�z��t�L��DK3àx�o<s��Sp��(fr�̈́�S���]z�d��g'������q�!/SV��v��:(,��e\����׿�{z��4�L�7� 2��P�z�c��:^���@~�����u��s���6��'�x,��Q7��M�k;�%�d#�2��J&L��]���A�I�
7���JRO�d=-�e��/�ư*/�Gk��璒�잩�Մ��[�V��>��g���v�R'�
����@�(�Ն���F����@���zj���8��U�u� ��Y�G^U 0�&����:K�7�%'��~�2=��I����/i٣���U��tY�̍��lg����R!sE�=~.���xP����3B�gN�.�8ܐ�.��!1��?��XN�+)b6Lє:��� &j�h�)��W�Uq|$�c�-���ƫ)��������`|;x�t����g��V��$ѭup��`_�b���K���WLIF�S�mzG+��#)��&Rg[/�F�E�2"���$U}󬆘�1���ʥKʂ
-F�6��W.�\�Ph,c�.ߝ�ܮ2��5�x���%�(֮�`��v�t�w���:\rI�2xK�.�0�3�pZ�p&�ٹ��� �}��mL���E+̔�Q���.�u;F
��) �$ú�������GF�?m�y�M�˽є�d]��a�?�"F��=4��L�H4Dk:���ԅ�N��K�G���y5D�򂄙�b�#T������=A/g%�P��8����n`d,��l��E�RV]����]�n���94�v|A�\	��@c�L�Lz���3a�U�1��pP�ܹ�}��h��C��ANu$�I���VB Em5^���K=L�"���E΃پU�����:)��n� h��i��8�oL�����.�E+f���Q.s���Ñ&_�^~��'�TP���l�:M��ֿ����$Dyn'�,�K���*�v8p	Dg���)%��Ĕ������4�;�P��ȗ_,�R��$,�
����5X�k̗��6�Y�##�4���i�q�_�T2��UtB�A0h�����t��6�(�����`6\mB��W0�b4�< %;PĻ��ɍc���A��K��sc�eu���j:+����
_A��K#���B�oqO��^�'<����T�'�����3L�����vr�A5���p�B�����Sb�B�u��趐�/��ձ-r�'=퍴a}ݟWn281�NӤ���7惺��ri��/{oO���a���kG9B#�a�dz�"C�#���x�[�d��F�7��B
`q�A�T#`�YʰL���:R�1��=���:ybۏ��O�7C���K7�"���+�r�a'���w�\~>�����M�>t��l��{i����!�}��y!㨽���g��-�NSHr� ��haQ8�M����M�|����1%�o���(*a��
�*Hs��a��s�+�SeS��jؼz���S�c�w�&Z���D�B��H�>�b>ѹ����	9h^-;u��d�/.�iDw�")Q��t�R8���["JCᗦطe(�ɾ�h�ԇI��k�C��&d��|����n[���w�>�7��j��-��w�2�-��U�78�{7DO����˩�wŜ�p�v�W��-��44�~B;F��( �1��:4t��3���*�ve����:c��F��m��,6�ᰮ��jj�Q���z^�̝,�����m��ک��Q��޶*��"Zg8�����,���et�?��U�����GJ5�&R�,