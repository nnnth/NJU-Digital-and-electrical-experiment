��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��tt��R�d��(� ��,Tzd}I(oCS��L�2�_�
�M�B\ɋO\1�o כ�_E�O6�{�.�_� h�.K_��Q!�WE5 � 	7�����5k�n�����(`��>2o[I�.��U�l�8��{�E�;����f�~�:&I[ē��5�p�9t��@N[����J�xE4��z�3�HHTC���zbH9����L1Z��}�G��04F�i�x�sK�[�"��<�3=�=+�[ � �T��G���	��eR�K�@��R	^樜?�<UR�qc��`<�8N25��z����1ޒ�utΩ6��Z���?����1{_v�З�͝0?G�bupx�Z����n֔z��F�V�s��D�� \��u����K�z��`�����>j/l8>@!l=��ľX��@]��{%����2�lA; J�r���Gk�$܏n�n"����LT��"S�W�E�La���qgn�2�p��bZ?�zh�����'?V�F�Q��8���7�ʑ;�bR�J�D�^ (��O��EY8� v�?K�{5��C�*�yL�Ƕ��ȧ�kC��&rt���Ƕ8���Ǥu�D����$|��5�)F���>�i��VAӖ�[RBC'z�����q��̀<?����D�օP�����k�����l#>M�`�P��� ���.Lwd�n<�������'�۹=+�}�uNs7S�CݮDFS����^�e��_&����uR/�+Cͱ(Rψ��"��T��̦X���̵Hn��ɔ��g���'���^;��y�-�eY���k1)�,T3�Ж�P����<�4�f*����Lq�S�x�(q����A1�s�	�j��tT|�_�%�I�t�GA��,W;���v�=�='Z�g�i\�}�:RW�I���%�����N-X���ȝ��LY��Z�@ �<�w���tA���C.��Y�����RX_�H� ��k]B�v��k��|�@M��Q�nWD��܄�ZE����D���\�`���TE���^`���+�j�+�pVH�bu>���"܋<��>(-�[D㓕[�2Ù�nG���e+�C���C��9_'0s�G˓��@���,��>�µh� z�/��["��V�لH:�T�$\�Ź���������R��c�ó���Rjڼ+���� .i��EO�Q޿�����H0�� @d@��ML��$f'K��o��7��9)���]�(2�Y���3d���+���y,���靶s�!)�� RP �<1X�����Ќ<\�wgwثU{ΩL̋�U�E��?�^7��Nq�ؓ��=�������y�z
�p.�+�wR�T��ݲ ���y�R�f���<۽�9*�����Pj�h� ���K��"Ձ�G'��6�'QL7om�	�V�9)p8�)\���-���_��9W͗�)T?VL�ά�+���H�.����G�%��tw�(�F�:J+I3%�ʁ���6$jY��rC�����������^4�Ć'�;����L�^J�q��"A�v��*�c�UDo�v�k]�|,&m���S���(��k*>� ��>���q ���HV5
�jz�	F�N�|�B4]�1�r�9Q�{�N&�x��a�"�����x �	;]�+bL�ı��AU<�䖹9���7P�"�b���J�7st*S��S+���D�����*��O���ZXohӭ@C����ԺB�~Z�:�$z5Kԍ뇫�i���W��C���Ё!k��ӂ��y�$9�/!b"�>ܰ��c�e�p�v��Wg��M��Gdt�@�����(����P�"�ta��t����O�r^�:��ۯ�ۑ�N6ړ���	T����U���'{⼜̇q>��"������r�Q�K�������d%���b�m~�������o�WJ>���|R-olw��_����CZ�p��ʸ\��T�i�e�H����w6���H�ى?��A(�2"����{�,XG**��DvRxC����Ú����lS[[���瑊���h�ȷ��L���e�R��x�'?1Ah`����jGGrNS��͍��e-��m,���&]��4�u��b��A���r�ȼ��E���Z���Ċi���n�W�H�=w�
�6-�/V���Kn6���s��|��~�-�2���#=�	k�>���l���Zϵ)kHj=}���-��.�7LG_�0yU��ޢP�1�p���&�<���(�d�C�nM�anr�T��DO-ǣqI�������+i�s�����A�i8�('H��l�,a�י�*3� �sE��(
i
wɐ�� ,���s�/�3���s0"Q��y��E/���MhS̪M�t���~�rU�g(: ӫ�ѯ���+��F1_Au�����Y�p�}*�v2�h�/=`�F��"Sq�$�%I#56��9Sl���ϸ��<CUh5�*q��֙���j�s��n������rTΓL����e�pX�7 ��떇�/bQ7B4d�����OLu^����f(�Fb<F�!>/šǕ��� Пu6	�<.t�F���V�uP���XM֙݈�/*ۺ(�ĊTI�n8}�
��#D�������$��ߛ7P�Y�R����*���튽��N���fT�b�CX�����i�n8xj�I����jrO�u���9�˵gz����9��
g�J��