��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��pi���Y�)h� +Dp�zXU��<<�w��w�� �d���NF��Jٯ>��u� �z`�h�v΋�N�u�ߘ�@��G��_���Q�H��G��C�A�褆�=�I��b��vK.���1���=،��CɶpU)�.��2ӆ�`���*�.�L^����5h�!�>�|�4ޝ�t�؊�U�MRJ.9Q��(�%{���I�¼BB�^s�
�i�%g`��Q�H�����M�1Ix��ɪ�Ok*�Y ��4�-w��y��[Y^\��*Nٰ$�y���R)	f�ǡ={�"zc$>f\� �^KH(�fC���\�|�&�c��yh�4`���U5J�k���?���&�C�J%۱k$֥
��j�4`�)��:����#_Rɧ�J,�@���T�bqkn�;d?�Q;}� ����d6��$S�z�ʉ]�:2���>y��iZ�k'p�#���e'Vb���9��#%�"h&��a/�&s3LſN�DҩA,灃ʦ�A�N`i�SjY�4�:�·�P���2g<U{GVq��,�2���wxUw�����d��K�#�ca���`�`�j�:���F>�#��@�N��T1��~���.�8jJR�,"���?+���Y�/g��hQňv���Y��r��Ij�?�����R/������O���X�7�i�?����KԘe#�@�Hq~��V�W�+��<�}��;��LM�t��]<�dY:<c����	;� ���`M��]`�R�ɍ�"Q��G/����߸Jw����-�1���'W�9G�WD�3�@�<]UP�t�D��(R�)���N�$�Q֠u�b
r��R+���P4��P���Mgܐ
;�:\k����3����C�g�.���j����p-�w����ѝ{�>&�����G��0�{H�ԉF��:�B#�f��,ꇧ�
�(D_Ш׶�τU��9j>�)Y}}�yճ?&y]��p�c7)�f�QE��-L�7֧��/��Q����-���$
2�?�ZaF���J@���i�>K3��g�5�A~��%$�Lؑ�C�t��R�I�\e�,�w���ٲ��#I�81�s�$�[���ˊ;^}R��K�>�gb��lG ����n�`?��g�qMQ	H����SE�vւ���^2U*��u��i����A$�=��A��r�_���E���L��!��	^�J����=эp�UK�O&7��24�)E��\�/=���hJ�淾�2���4!t.��%]��J�U+�,m��c�^�q���d�`�x���f� �a����%*��T���B"8��o��A�5��vC���n�{�߸)�b��Gf����[K,���w��������w�%IQE.~	/\�ӆE8��!kW|�D��� �v6���������*]l�'��U�h7���9�*^��^ɝ N$>$M�HѠ��g[���g��6&�� %�B._��ꅡu�ۥ	-8�WcD4H�L�o����C�31�}5Tk���W0�0W�z0/Yc:耻d,J��T�'��Nc��@I���IoQ)p�-�������5�i��O���-���ڳҙ�:��,���w�-<��aP�Ղ ��G
��*[9��f��	�qh�U{C�mFϱ$桲�&ݚ7�8}�����蘟wߥ9�~Vb�ceG��me�'�N>S{!g��Xƚ�a�G���|Bp��?C=��{�� �F��M���6r�:b=�皡��Lk ]�J�=p9�7���߱Ϛ�i���ݘ�@/�3�f�m ��7�;��+����=�����KP˛⪇T�1u(^n�����0zp�;JK����
�t:�Ĩ���^6����i�+h�Aԯ>\�"%0���^��-�V���ۃ|�VR吔t���I��S�L,B�2�9���l�q >G��D�8}���_N�y��M�G-�D����q�P�nb���>a8��s�L�����/*'�x\i��X;���=f6�ؗg��Ҩԯ���j�����6�9.��
#ϥDa�Z�g��9#g��C�)$vx�X�y���#�X���(?��ĲZ/
��TEE���������lO�;t+����j�\H$���V�n�Gb��d$�e���'�4��f�{{�b�G�J��,hn�^���1�Q���U�4\^\�q@�S� WX����b�ԑ	���fjl��/IW60쑶-�<�`]�3��H���������:�Q���4��GL5s�
R�=J&H1`-��T&ŋ��ؠ�E6�Ʉsm�������X��<��r�d��&�/�o�\����x�;��� :�V%���Y.mq������^���5^{)a�0bC���N�r���|�j�-p����+�:?c��`��Gmj��h(�|0��L=l?�I�@�v-ގ�~}��:�h�]�օ:�]@jh��k2�o�*�i��3R���w�W�zTE�p �i�@5�D�_��@=M������LI�2��{	��c�'Է!]/�c�_���.E��� �y_��{
j��rl1U��S��:+A������,�CQ/�ަ�X, ,~���.�+��Z��9��boL�.�|74ڸ�):��L�i�O(�*���A�_���o,�_X�G�k�}K�$cM�������6�đk�֩����Ʃ}��!tĈ�і��x:�o=�X&���e��R/�Ɨ�҉gď��c�B*i搯�垕3�DT�?�R�&hiI��ز�e�b�h��h�4o�����a�z�ˢa��XJ��	��nH2	����c�z" Ӌn�[�ҍhE]<�N� -�t��/�/�M�|��8�*�'	����
˓���x��'{E�i��N1#I��n"�XN��0�}g�œG�����x�5�W�hK�(.Wz�,��&̱�r
����
@[+q;*�8��uߡRO#�S�"�-�v�Ia���t�6�짆>���9�A}�=�1��P��)��u��|���j���,Y��:�%�o� n�#�~b�yp޶B,m�<�m�0x���V�40�H(d�e�2a�I�-�]����􆦗͒80�'��tF�%xxv��K�&�����Fx����p�ۅ�2���O$d=krwh��G�2�� P��%����v��ڡލ�����z���#y*�����)O�����2��w��fƵ� ��uy�S-ij�����G����=�3Q�� ����}/Wn��t�O
z���ۃ�gULY�GC��o@�	ݛ�;I�����2�d>�.O�Fd����`Q^�GG������D�_�E�Ӎ��S�%ի9�V��bÖ�� P����������P;�������(�x��o��	��$��#�n=l�ۄy1�n��+_���sMR�&� �x��"�ѓ-�:G�8R�-�X[�PW��w�s��7��?'m#���졡�j7��\8����;WI��K��3�>��sU�v����a������¸�*��o�&36t]!�i���V|A�����[q�KN�ͧ�s��H�ȄF�_���:��8S�9�W_F�9e
�J�*�Cf��▃L�Uֲ��*_EYS�e���=�:�`ۓ����y�g�+�d_�N�	`�ȯDq=ؐE�ҟI�qx��q/��G̀��w3-����>�7��$u����'	P�JD���8�H��h����W�%d�����[P8���8~�d.�OwH���v�)�Oe�`cz��d&v �'���\m�������k��OE����G�����F�}oG�"�2o�	�| q��k��O�S���n
�'�~�P��9\��(�+��w.�Tb��"�����Psۭ��}�e��+�c!p
>y����9�l�f�m��/��k�b�:!=���^s�F�j[5�"D�2���]+x���� �v`�anڙ��%���������,����������ݒ�r��v�OE�)�B��Y&XT�y�שf�]�'�J�a^�,�c�m��s�����.��c�Fn<ݜ5pe-.�Էr��g���'b��9G�Jy��2*�26�[��Е`�u��'ħ�}WuG����)�	��N��~�{w���h>H�~B;���WѢ�����UF���hΟ�|��; sߠ�^�?P[I�̮�ϱ��T�=��&Jl7�){B�H���k?��*�&�����G��9H)�;�����Į��	����qC�e̓Z��w�4����	�&)�S�=P®�6T�ɑ�߷�7w�x?���;~��:�,�Q4CJ
&r04���D��I3T�rk?JX���&��v���Q�;����x��,�@��n��#
Wf�!NUc8�\�e���=�����5�Nڜ:�#��*��ޤ��D�X�ap�{���<�������z�tsQ���8��m�f�<ܮV�	/�I�f��t=�.�2�j���!oP���8><']+���\�$��6R0���RK�M��	�}E�+�3���Ҍ�x��,�B�E��;\x��!�Fz��W4���5�ԭ;K�j��-;��H�jH�A�r!�4�������/�F�U��#��+Y,hr������
�2�⫾Z�)�Z^�v�  ��]�:gs��z2�!Q��\���[�_�>�ք���B�&�uQ񤎈��J����� O|�a ����;h9��!5���^��*�繳��ڙ����ß��T����H����	�2W�/���6ai�柎�/��[Qw5ă���0]��ԣ��<�r{���Jt*�h]}R���m��E��b�����.5r&��Ë�%����<�5�Lm��ƅ)�Pl"v���k.�V�������s)\k||���H���pL��������kAy�n9�� ��xh��������j�8u
���TERC�w��CXz(��:�Z���`��z�"�4?MJ��@�����W&1�wH�X��QTu}��Z������[ L
7t������̬�yZðc���Fx��|�:7�����
gH.�u�B���ݪG���9�Mg��i�3Ǖ���H��nJ���tk���B���[�:g7#�\Mfm;�\+lm�d��BΚ�+Z���z
�}kd��4���3��g���|�:��6a��)�����J����ETĚ�9��9�$ԼD��ݛ��9/��Z������nQ^�:G�����{zș%{܈�{�]�UE^G��m��=�-�]���<Czfʸ�-�A!:�ʙ1�S�[���%E��AVE(����t �7��W�P�*�L�H���4Yƴ��j��/0���ne>�f�єV��m���+�-TՋ���h�Cx�2�(D�0*>� �|IB�4�!�z
����2��#�!�(�s�a���'�8�81�JY�06^��D�a�%B��j��f����5�n�7�nE�-�Xc �Q�?��Nv��N���.�c+���ז�;"7�-�$:�p����u�`��d�rC�-�m��ٲ[a��9L %�HN�ܴ4k�4���K��~�K�	����R�$hP|$�Ğ�i����ƇE�%��侨�m�f��cR�"˶�v�lz�av�y�#�)�: �����'�+i���1�Xh[L=+T������J���9�W+
>/��2¶'�.h���@�Kl��}�|��.\�+��9�R.F�7�L$�R�t��`�Ny)�r��Yz�R�{�$�gXkP�u�R��?��m[�枤���)!�(9b�sS��T<?@���E@6�9�ņL^ �k���y��:ގ7A�ͥ���ҭQ$u����!���؀�}�
�0S�'WQ�m�fM�W�[������U�3��Y���`Xd���"�����N����567�S ���=�O��W��yD�L�~���v��u\����WQq�Di�L��[�6ft�0�oS�6t� ����1^��w�c���(�?[m�n]$2�O�����{��	�{0g
�־��3�na�k�"

�go-|VK�cm�O?��HýA\��n.�+�Nsy�E�����W�T�̾mjg��[�����K�B}����7|��#T�q�����O �40T����,��4�"�Z�6x�i�g
��_F�Y,���6	n�gS0ل���r*�K����,�e���^��j*���D�����!�ksJQ6�3KB-,�!���h��g�i]��RI��2�Vhd��evn�P�T�aa<��N���e'r�b2X�����(o7�x�إ�Hd,� �E�|A*��Pپi�KSmгȕ��l�\�W����kR����/�D�{���Ȱ�y�N%��ʴϭL�eKt»�9R.��ړ<�^�N��+ě|V �׶n��P�z9n[;�*ǖ�V3�ɍ��^��;7�BIP�o��7��B'�ڋ ��8�C;I,Mp�6�S`)Jw��z�:��U՛��W��p^���Y���;��u�)��bN�+��l�EF�g�ԏ8h��2Fi!FĮG�CM��^��6�
m��3��!z^y��(��0僫�C�`�4�v���x���n|�X�F�XU}bq���M�>������y�JX58�Z�/�,�\n�\
̅�f@E?
5�8�>l�:[U���H��(6��~rzI&�r�݉�i4��P�/�&`���4]�3i1�z*�\vB���34r�^bD�����Crh$1�ʹ�ȸY0�6Cj�]e��/��x�P��xx���H��Ѵ�^e�_ 
��ln��}B[�^"�s7&��,l%]N���F��_�/
���&�]�`㾣n�H�Hyv��w��.�#B�P�r�p� ��N,5֗����s$8ִ���a� ��	�￾HbU%�IC�.�u�%��@�F�jb:��.��}���M��1˗+q�a�L*z���#�R1V�|!O;��ַJc���J�J��]��&V��H��b���B�G���*���K�:%�E�(�9��B�=�?n5������P^�����c��Q�W��b��lpTrG�7�C�ܩ�`7�15ho�A�ȼ�����r�73{��O����Ĳ=I���Y���[�+�KĈM9NP �Fc���xƅ �0G��#�s��lx�@��9�@�S$�iw����1�����)b�l|Ic�oӞ�.�����V�;����Kg����58�ցQ�4+3/��/��~�H,�O�`��d5�����y�7�m�Ϝ��~{�cO�".�r�r'Ε}�V�b�泚�o��pz�È�R3���%��+>ه���x��}��O���ӱ���L�)���g��D>أ�mգ�|�{o�U�}bQP��������rG�bn(%��/ښ)�яA�<���Jr�2mӱ��[I(��!����'�ݚ�R/����*��<~��
�Rc��R�T�)vkY�?��t(4#?��~rǯ�,4����#�@�L�&>��W/-��jش��I���e�ew�/v��� ?�O���� 6��hC!� ��c!Xr�v��ubX4���	\�$2͇�i��-,dGIB�n�X���Bϫ!�]�E^q.ާ)u?V�Y^�.�W+jҪD��γo!r,�	j��{��q�b�m��`�PQ,��`!����	�۸��6a�f�\]����X!V��u��H�L����P-�ތC�q.:+�/����=�H=��{O},]|���u&��������Y�'�l�Dc�ФI�9�!�ݽ0�ޢ�ʈ�P����Y��&�GXՕi:��@���M=k��U^��(��K�8f<L	��P��eg��PV��;�t��A�1����\=E�4I����̽H��2ɰ����mY������b�[�+ޥ�Y#�EX��]�H�3�xR:� f%/Qٲ^���"K�����#�/b"����x	���m�V�>�����a������E��I1�#?O�[�̺����>+�}�r���������hj����R�t�~S-i�m�Ԝ����'#���2gK����`�p5!~ǘ'З�:�g�8��n��`�;��6�[��=|ʀQr�Q��8��-+zH�H���z�h�8�Ⱥ����{���Pԟ�kۆa��+$ѻf{�����p���V�i���+!X�pru2�G.�>\&�ù���]f,o�	�aK��M�^���x�ސz�\'�#g�:�}ӵK:��Q�AW���̗���BD<�s]��v0ߵ~���bpM*31v�qΤR��0a�����U��Z{�쵥�G����Gc���l4�������Q�0����B����A�����n�!]֗�����a� N3U���aߺQ�ZEb�v���߳s�?z,�	�$�r0�4e{��j�����j��_�$�Z6�R��a���+Q�z��'����4n��%EK�G	Xt�F����d����k�Z����GQ�������6%7�� ���2�l��5sz�v�I��©�ؙV~e?2%l��\s���,v� <fmHu3P��'���c��t��k=-|���8Bz�8�;�Ζp'R ��d=�U��WmXj�������ׁ#���C�e�)!����B�b]�#�G�t�+�.�7�~^IC�zp.xiک3)��h����t�KL_Ⳗ�N[P��,�dK��W_��H��	6�r
�jK�ε�"�̽�  .��X���3`��=Wеn��2,�WF�GT!�cz���q<���H��UjE���OF��u��J�����+�T�ͶtYz����Z%���#'\��J�����}X��|Zq03�Y\����G_�%���I4�$둾[��$w5� '=_����"N��ܷ��$m��ӝ˙Lm�4uJ��<W.v��:!���;D�c���?p~�R�X_0ٌ���(�w��e1C�������er�A+�V\q�fI�/�v$Z�3���q�F%a),��G�h����b��y�N�	�hV�"���W\��0a�w��-^)���Y�	����;��3U�QTp��~4&�r|:���L���I�@z��v�S��rg�#�Ф���1~��X�TpR4��:��<&�	���[ģ&�Z_��^�z���g���Y����] ��*K]����kt�06�p�H�;Oyh�C��K�psu���G��/W��)U�w|���of�Ë)�ZK��j�.��`C���V)�]rB�[�%>�M̌p�}LL��L���!U(�z��;�$-�	���pdٽ��C1?0�l����Y��/O�y1Dmީ�F�uMx����ГMB+�B�q��X'�lx=��X8!��;P|=lu%�r���=��$^i&l��	
Qh�CuR�2�1	W��9r���Q�i�?a{O�����6��.���9X�籨���UL���>�q^�_��	�,$U��7\" ���*���K��e\�F�R�A+��w+g�t�r^��8b�1B�������֕{�9-��?��~�ڡ�1�륖h�?JՒ�a������H�j��$.*�7��&ל�b�9�YO������n�����{��=`N�Gi���,�-?��)i�P�6��Q�����V=�e"kƵn�K� L3G@J�1��m�{^�+��=%|���Ħ��o!Y:5Ë�9�Q5�mt����0��7J���0��B�f�;��@�	���\Ѫ-�8�L/։�ڼ^�I_� t�P��ae��1jZ�O�SV|$��O��ؕ�cd#9��L@_�8��J�~����^�2������R��Ov1��D&�CY�^!6�o�T���Vt)�9(|��אO%���דejfrS	%:�����"�'/Z��"q�NMJyz��z=���@2���+Eіg캸����B�@��u��;�m���Fq��x��]@��r-�u5v�2� N���+�|m��:���������g􂮁�KaL�T�,[�����PE���A<cJ�\߫f�ڍ�e���!�şQe�'�L8L��;"b�(��n�ߕj5|��$�zV��
��}k��]8:���~x2���Jw�Ho�Lu�X�s/0i���p�4��.sW�~֦xA�q$��?���905������+x�Ds�%�?�ZIt�D�(�O��י�V�u��Ii��B;5	���D
��Šm��K_&,C��;8��%��<�r�"�L_fho��?�o��Sb�6�/�?�v��7wu*��ë�<=����8o�`f� ���+kD�"���v�ƻ���h�����b�sC��o۝x.�T�؏g���/u/)����a*�b���� �z|��g1Z�y7�2�@��n�M_j<����ק��l���Iܱ��Z��ytv�O�$��K��+`���o	'���f@�� ���)0l����~Z2��_,v�l���H@����V�~R��E��DWq���{�$��AC��I�������2?L�I1���*�DPؠ�!��31�#$�0i�����v4]�7ہ�E	J�c��ej�Z�_��Y��͂�;��U�F0k�C��d��6c��"iâ�O�b���	&e�6J�6COP_�H��>m	c���m&6�3:����C�F�7)�;��a.���&7 @���������|~bj��d�5d���+W|����{����T�mä�,PW�w�q�+�ʜ�z���o/��}d��tY#%*���(	-�^��>!J^���)��BTN����e3ޏ�9�_Z�E�R�V���^�zԒ���hfQG��v?�Oq������:k��U*1�iҴ@~9:��-��T��a�LK�d�ߥa?��8�i��2���N��+.��)`S~kw�[=��
ԍQR2��D�������7�>�Z_�h���� ��ѐxءb(�m��k`�J�*(7���겼��q��A��_e��`�0�vy��,�VnG�`H�٠༼X����9�f˗��1�Q�_���$�h	��X���'�$�����-o��(ץ�Rڕ9�����E0�B�g�\4_^���_s��5(���
�f��ܤ�$�9"^B�>AQ�A��<��$����Q��y��&�`{�bPP�5�ԛW�`����G��{�2��o�D�ז>��N} )�F.ו7��?9��"���f�5��<��+p��X���ϒ�~С��qp��՜��2�,Co�����������vk���V�����
�rs�c��r�ٻ����?ߡM*��� ىaF~bQ!b�l�'�o&�����\+[JI����<+��ʂ��zLB���O�6'��� �\��g�z��Z%S�9� W���跅Rw���g�Bx��gTۻ#D��Gz�MO�l* 隚?���2&a\�{�03T���W3�OE.����R��cE�ף@ߒy���X�j���ѣ��*>��ߟ�' �x�t8 8;�y�o�ֽ�p��Ǚ�$���Ę@��C?��U������R�Q�&�O��i��OY\ĕ��Z6��O������s� r�D��eR(�<�r����h�c��i꾧���������=�ƮPn>��J�%;2X�����R�K�Z��Q��޾���
�@��v^��U{)t����W�#����uf��X��� �6�"�.҄��/Vǻ�E�����}T�>׏���+���{U�sG�1xB�q1�E�EN_rDϥ,�X�(9����!���\���?;]�"Q�� g�v^�!K�L�tkN.V�Y(��v*D��ߐ�7�Q��Ё��-��$���w[3{��n��)3G��|�њӈ�LA�}�G���@iM��|�)ǟ�l���@}������4�D�K�zݨb[h�v
ɋ�;�����V��.L��8�<���_���1�=1D7/S�810¼�G�Į������U���X�f	��Y����_����,p�Ty�;=�{^� �	��������Lx�_�a�tA��ʂ��0�^D?�D|��y�ƚ"wB�.\�RΛ���x��mσ��i� ��糑��K�����x9
�?�]��!��r�f��n��͈8��xh�Cd]�\9W�YkG�S�G�����,�d�[QS��|�UaJPU�r���R�_�c��yd�z������H.�g��8�w�A[|����p'��2�7[Ὶ��ӣ��'����H��|��Q?���� �H�w��"c�\�&