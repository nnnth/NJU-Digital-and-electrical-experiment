��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�E3�hoA�zFҿT毉Ua��|���~��r�*�F��7>��������K=UP�=l>b�\*B�E���3�^��m�(�G�wI��AP�%�-�|�a8=�JS�o��4��L�	�kϏ��:���G�tA	B�l5;cǡ�t7΂Q�@q�H�ښc�6�l��Y������$Nԕ9�2���(�/;ʠ*�M�.�+b�+K�}6TM�� ���������t��>�z�J�.��2t�����z��]eܖ0ڻ
3z�g�>џ|
� U��C���Z�ސ'oEF?��zy��іX�!y�Y;�uf�Q�2�X�6J���ƥ�.�J0^�w6��7:�&D{�����1V:���*�Q;�̕�Q8��U#ݕ��u���]^Iă��?E�j����:l�120��NT��D�'���A髄f����@,<�%�x��S/4̶:"��+r�!s$D��ѡ9%,�'�CR|7 �\xG�5P�V�s ��V� �/�	ec�}��ye#�$pOn�����l�*uK���C��]U ���@����:�9r�h�z�2��� a|��~��iw���]�c�'�%6��
�9�������H	�KQ��ުĊɰ��[T���=�O~��"���c��Ni�;��?��A2�~r������;{v�����H�v������MjV8�%�����HG�ԛ�]�~lL���M':���t�PBE\F��j����Wg�I^R���R]����A����m���{A�ȴ���UX+D"K��J���>k�Xޔ��X���o* /2��V5�^{aʼ�&P*�Z�T��'`�e�_��n�ӡ�yJ�
�/(����a92��n�^p�JP�d��E� x�����ao+z�B({��.�rG��V�7�8��]mB8�?����;��-�O
m����d�)	�&��V*�y�2b�Z����"��c��K�l�a����Q���D������>�_mZ�D���l,ޡ�-4b��%vh�EW�7�Fi6
z� �&���\��qf�0Or)�-NҮ�ȇ�X��B�$T�Qd�l�d�\���z��rif���2Ljmͥ�=I��rro�LC�ɊB	��PԞ��1>�b�@���{�qN����$֫�R'���6'�ȈzwLR��̱�l�d/��x���%�A�1W�8N�,�ĜW��eJE�H�R���P�R��a�u,T+�� �S��M"��!���M��>"5�3+���J��{�b���d�y ���R��x�f �	�f�R����E�u�0S����T�\!_�'���疪�W�˒���(�^hs�+q�t��EM��!ej�������N��A�Z�I}�U������˗j��E8����>�|&MYZ#�h����Q�t��«Ƶ�5U��v}kFm\���6/TF=5P��3����Z��̨3��j)�� �?e�U� ���"��O٤�w��|�����JJ����w0���-kn6����j��L��c5��;���^@��<K���ޡɇ@���������F+ba�~�������������ι��G4i�U��Ru.�$�p_�d��,�:`��|NY-��⳨a�xx@�+����}�b�<�ξ2T�z�~���h��
T�%Ə(��)��z�3�ǡ$�-n/�~�Hx�$�W�+���eu��ӗ��k�g����OB8<��R�qWtSs���[��B�'Tģ�6�Q�3��i�m��ga��!ij��9����2Y܋.����`T�S��׋<Hj�Z䯩槸��
|\�H�댤��@�wf�Lnۘ����U`.�L��а��&<�w��e�x��+��{���=���s����|��=�W�B�C��F�5�3C�&�������X]��q9j�z|�$��$��'O$b��Ϫz,�g�,;:(�*H�&���_�U�L�<SPH�`�C؄�'5�w�-%��~�sq�Ɉ�����}5����fߒ� ��WU'\���,���F��H��1����o�"���)���&��@���B!ƴ���N������aMb�{�@�pʣ�/��h5�#�"��}��V���,��A�%-����~/�.��Ƨ��ҏ��i�_ڱ�8ɀ������Z����Q�Љ��]�@�=��������K>	H+�7���9k�Y���8��F�"�)5$����h玚�N@��NYX5���!J�k�s�։�h��B0��3����ü���2r �Z]M�p�x���C���~��ڼe"�)o}K��~%�??�
���w#���C}�n=��o��l��>ˢ����(���k��t9˕P~ρ�i_$�������W�� ;=�"�a$7��-�2��t���A�?�ƈzy�\[ƻUtBI� ��J�a���nW�3�1qc�����S�`2�(1���WP���t�x)lK�+����ɋz�R�p3$�W-���B,��c�����`l06>�����ܧ��*āF\�c�h���=A�4+D����9 kV#J_�wH�)���UNF�̥(���K� [�3D��U>!'�k�iP�mw�4"ω�k��0#����Й�辅�Yz�����Ϟ��g���#y#atY�����k�ƛ���f��@9�-�I�Aq�����)�e��"��R(���G�i�bL�8��c����m��+���n�1�C^d�g7�g�#���8��"��Y~�@<`�v�Q��ܹ�p�O<=�%?>puF;��ş�)���V��V��|�%�`�dNd��D39k�K'�ȭ}��,*�HA�����6�P�sQH��r�<F�m$�o/6��Fa`¬р%��s/�=kk7���~&��*g�R��ڬ�Ar7Ni��y���#`%c{v%]sT��	�l��w�V!��oL��`�SG�f�#7����Zv���"gȆz����ܱ����WO�Jk������ ��(���l4�R�U�Ns�N�+�b�[|��jz������g�����>���fңu����)�Hxq��*�˲�N�� ��4��<XO�>��6��"��e�Ǵ6*���n���6���k.��ӟ_���!'ǅ��y��xA`}��	 ��RԄ/�e��?�\b(0���&�����8$S*3����jj§ߟ4ǀ���q��?p`ү?���V;����Eó��*�u@\M}����7����'LY5�kx,�P#I�	�����ѬY�%?�?�����r�߮)]�o(62bъt̐�n$�`����S �g� |46{��ȳ<�&\__~� &GmoͬL	T���s8�V��R����ruu�P5�7�i%"6�����d8���ɤeʓ��.��=�K��^t���s�HQq���D��B��V5��ۏ-�e���Ln�_7��ҳ�ks���t���Y8��=ˏ�.�<i��XXv���Y�Y�w+�=���h0}����/�l1E�P#Ь�rt.��&TS#ֲ��Ϧ����oH[\f��3[g���9)ж�e������n��m�}}���IϢ5G�-U�Wz�VJ��N\.Z������٘VI�wڃMb�OJ*~��/�As��먪��;�X8O����&�>�!�a��K�2���z������ا�������x�oL�o"�E%ā�����ڗ:��>��cilA��N�~��1O���C�ܨ�p�dHcW��>ҲQ=�"����0�����m��-��Y~���p�C8�9U���W��	��t�{8DER&��HLw3Ũ}�=fU�
r��	�;���2�81�n�ɪB�_�r��;y?�qI����D��݈���GMB68ZS��� �(J�d��}'����%b��Ս5t���D�N�ߠ�-ÈEfވ�Lh?ŭ�a%��5?)���b)F�
Дx_8���eM�&o�ſ#^��k�^;��&���Oy�s�9#��e����ϨL���q�,+C���ɣAȦ�����Jhy��r����e���K��p�G����!A���Z�yu�V�V�EsMT���� p+&ݕb~�B�0sX����&0�S�`�y���n����h䬇�қ;��Mn���U6���L��V�����"�e.P3#vgxs�Ģt:�|B�4��3�2�5�}�J��-?��\� IYR"/֦���)�N��\������O=7�>&-W�G�T����02q��=(��#b��Jܵ7"h6e�BS/�!`���~e�
��祰�c�'�L���)�qt������z}h�q?��'I`�����\"ijsCP�n@"s�%�V�8�f0�u:C�G����"-�DE�����y6�q��_�=���`�'�2	��f��i^E�Ĵ>H	nՎGe�XR��UI��5�_J�a�_���KƠ�iwA�G2�4#*��1�n�������D��,�\T�ߞD(��~$B�1����IX���4		B�r�\�(����顅�?�����Ƭ��Jð�����ǀJB
��t�p^f�r����G1�ޒ�Ʉ/�@[�[���g-���.��b�&�8���G��7�G3��X��Ya��#�n@���<���%��Y�j�cq�JTdG)����P^�M�mJu1���*�J���a���P���R����b�H��G��7d�I]�_�	,�{xd��J����+oE֣X�E���%�ɶHR���/���(4O~��z�8�t� �Q4 �Ԡw��}`Z`�\���+�[�@�\�~��u��'%x2�<L�8V���]�T��Ǚ`����&���� �u󽈤��i�-S�Fv��#HӼ�ְL:X�l��_ �96d��">:��vZ���Z�r����R�'��>cj � ����)ǃ�/?�����J_F���z�'~�)��tZ�A�a�c�i�<�^!O��zUJ�G���S��f��f:�>MZ�^kn�C&Q��*s��uD��uIwʕ�u�s-͇���
�� �RB�`S5>5��_'A%X�*R�*���N�pb���K��:u���i9��D2��X�%�c�ib=m_�G�Ji�-n�=n����V�W7�aWY"��f���
k:1%P�?�B�n�?��a��Ɲ�Jf rG'FI�|ׂo����I���gL�k.t�Ga�l�^��c�,ˣnk̅�͉M�'�u�{�o\��Xg"���V�/*�9�Qy�?(��=]����d��Y�9?P�Q�C@	��N+��7#n]�_ƄVq<ic�-��5e�'��(����v����AM�W� ��o����@����{#�&Qn�DA?q��M�$���9N�A�v��b�><OY%�{X�<zW��6��; �h�۝���I�6����A�v�=�}�q��a
ij"B��"�~{��dB�'j8�u�ÿ��ԯ8 ����hW��h~<<�գ��
,�jFх�ڕm�+�F\ݵ�!�%	�҃��:mŜ�?�M ݩ��i()
+�}�ډ�8��N�Z��f�� ����j��W~fsI����|�4���gI͂��'����N4��C��OP�����ԕ�g��ɏ.�׻�C�9�yE�� ����`��_g��%�Ov<,�k�r�T��A��[�o��GB��-f�1mɛ��1zN��gͧ�a���������ћL���'��63�*�2/����T��iI���*��]i�ȯeW;�m�ƀ���Sc 
�<�9��s,�r�%��U�z`}z������O�x�1q󩝶.�2�,[���N��� ��!�tD���z��.QKI��;ȃ��5�����i�Z����ќ�־v(�E�:r�ĠE�vK��D0w���Tw���$:�!���n����A�@��-�a��k��l2��K�zd�������9Z?*��I]��y/��е��<�pp�"/����nᤫ�9��4{HĶ	�5(��5�sّ#��F�	Y�{�O��\��#�*7��j����6���F*C�}r���;s�H����U?c��峃��ׅ�d;ע߃�M���(��&�P?t��X�,�{�z���e)�+`��'-E��"^E�gC�♯�d���W��x��N�l�̴��f��X�>/���vK���1"��uQG��n֖��.'�+T�P�F��4FN��-r�F{h�����9��tJg&�oY�� I�eI�k5��ӎ����!(�ˉ�@�;KB����[?�gNХUK��{��ma��'�_.R�"1�y��p��2W~������n�r��it�s�J9.6s�nV��M%e��ߟPG��BY}�C���������'���eJ&�w�4|���v���_=�w�et��X+;�]�DJ��=�7H��x�b���/O���qu����e�X��X�GO��Cf*.���|BFk���KjE�я�8�~$�p�S�^��s!.(�b���,#d��k1�� 
Ϙ�cd[�D:}Se2���e��	�R �T����(�\�-�=jM�Sj_R[�S��wM����<E鬳�����@��mT���DKB�Ơ�M�:^a�:_���>sn�=L��3�M���톭�o�]'�N�����Cyb��y(��H֏�a��=	m�zc4�R����~q�'��73�.c+|���%�f3��K�h�����������.q�֚\��@,����}2.����4�@b�ކ�4���`z�z�}��W#�֐Ck���i��U���m2�@b�0�ͼ1&
@�a>�[)��4�	� 7G�����]�?�f�2�D�,�1��� @y�X��)?�����b���r��\e^F9OK�ÉZD�M�Uvĩ\���6�O�3�l����s�^�S�v�Z	�)���q�m���$Ul~Z|쇌��!�3�~��+9��
����֢�t�����v����6­������Ф-�d�#���l}�[�0�+���Q��C1���ò�5Q��<�.Gy뢑��B���R'O����������I3ިP�v��v�U�(͟u��7c��m:gr�[q���=3ʁ�g�����p��qB�܁�s���l�/�Gcrwhn��k�h+��,!b�K=ڃΔNy��puǛ�7��)Jf�U.ha��:�����������z�Pb.�J;�2mL*ud����d`h���.տ��ûҨ�j�v2Ɍ	��9�yD�h�o��E��é��S��u�Xʸ�|���o�ӝ�G�u/��==S��f��B��BP������!�q!�����A7E�0��ؒ��q���N�]�+b��5��N�����Ә�Z�t^om���P[�� �j+��R�	�m\� M~�Y�J�_
��A��tSJ@�������ס7���e�|�����Q�ʼ����i��kBe�L�����������������H����=;�<V��tZ�&�yP|��/]����%���@��b�����Η�5�$���54��H�iw��Ԝ_�%.�$8�2�Z�G�l��[Tt�&U0���W�{Wl��M�y�Gܪ	Z?�24�@�J��(��hh}�U��gD��ԯ���wf`�H������[f��-%����`�v�h�;+�L)8������6��o��n{�kSArC��a�ި/���%n�����Eb&���?=����лhϏ�B1+��Z��p�j1�jD�u �{U�G=Zr�u���6rWtMd1:i��.���;+��uq.��;(]�Y;��ӹ�ɇ5�]�֟
�Y��Ęq.�[i�0UF����V+���]Bo����Wo�4X�-J
I��8�=R���rG�����obG���f��㏽Ԣh�X�7�&�,��7���xYdbo���B�W�"C5.,O�� ��g�O��%KZ��nI�W���V�=Z7L�m���藧��X�)�B�7��z*�(�J0�_B�s�1Kv�9aG��{���P��3p��)d��<�c8�c��zR-9��t-�SRZ�]L�턇�h�2G��Rd|2��N���z�chh�l���:��v�	���������rg����e��:ׂM��^��7�I�Ϳ�k`pm��J9�y�b��b���s���ņ��1*Rȝ� ��!�� F�)�1�[߹�[����\����I��L���2
6:�i�v&#�H`���X�V)�:�껻�G�s �)�O��� R
J��<4�Ϻ4ય���#A�������p�7��8p�fW�R p�$�=`�]'pǷ2�h��|��G7�&Vz|%߾h���l��#�Y��H���y�DE��	�U��u�A�\�C�߂�6�"�x.蕳"�ִP�;]��N-ƌ%1���m ��X�T�x�0��P8��uR'awtEM#�i]�(s�GL��%�ܕ'qP��t�i��5sSG]�����0�M܍���3����.K�@�� ۽����?��h;Ц7�k��Y8E�X�t-^��p�*�1�"��۱�+JD c���_IC�HP�<K������mU��
K�����FD����&�0��D��2��!3�w8N��$;hq�X���S[hu:��J��U4�i&Rn����&�k��c��.!a�Ǯ�T��vr�3��kAb�"�0b1.x�!� �u'Ο���ab5[�TZ��P��i���S�.*./b�����W= �kޫf�����;<?^�Z��5v�� ��ڤE�c+�.����/����r�����{</4	�רU=����SF�W�ŅG��R�6�w~���z	�B�ܿ�f4W�k�7�2}ؠbi�j�BB���S3��5��jE�ŖX�v�����
0x,��6�M�w{�8%e{ �N��s��"	��ɛ��~U��fc�_�2Zv�I�+ ����t�f���Ky�����Ĕ�	D�K���t
k�:YZ��\���}�B%ֳ�O'y�v��OSz��_�����;?�,�*ю�cGR�u����m�m,HQ�*�,��8���CeeL}�x'�={ �mXX�bH^~fR��y�S��[{ ��"'���cLUvE�Pv�0,����$�!1��	��Y�t�Q*`%-�o�<Fa��c����C�O��+f�hk���_M8Q�O�߿�.i{�r�| �B;��h�r(L�B�c-�%��Oi
R���_]�@vR�\�i4#�k3vG�4Ֆ�N`�$#AS�۱�n��:��6q��w�e�ťs9C����G8N6+Z�������}�K��\�'�x]
:z.� ���5��d��x��6G6j�:�n6K(�^A��?�z# T(�u�cb$��b���#J��Skõ�b�[��8��<C���NZ?즇!~��q�uÚ;Fr��6�ZL�!���=�c��]�Ne�A�H��&lpe�~�J�Wv�-(إ���!��
*�*�������>ǩFD��L���HGkނڹɑ}�tg��54���e��ߴE���F�]��C!sv1�ܯ#`3��i;�%3���
���`�]N�0�y=��$:eE
W/�S^%v7ώ+l�w	+�b=��ܠ�[���$��#  �`�E2�S���`�P�4�_ U�ʀ�uv$�'�>Y�y/2����T,ĥ��7�b��ʘ�|Ec�I��A�J��r�m3��ζ�kƚ�5��ρw�G�C�J@"W@1�%�1�5?9]��	����1�}#&3�	�B#����q.���|ʨ]���-���؁F�_�k��wR�c<(�����(\K�5�C[.۲��h��~�'����'����K�%i6aБ�siF�}j�6i��"���М�����@g���"��v�95A�e�H'��^g�d�W�m$y��=����B�{߶2QD�k����-�6��"{`
�����ˑ��( v������ |ˤ+E�����,}�C�:5w��z2�G�j��<xp�>;��Ӫ�i'gL��L�R�(������\���,����p{>�����&����;$��1Ñ�|%���}�����4:'��3v��5���x�)�{�w'lE�q��^^���A�uGZ��@ڍG�5!7)5D�� Xv)��&ucBa}0 �iF�rn�	�����~�9A��Ϧ��K������asq�/*�,�p��p`��P�D��e���q��_5�-���
r..�+]5�눔ꌕ �,���q9W���1�f��22����-�NU�\U�YL��i���Fk�B߾�Vz(_=�	0!u{1�>�RT��Ë́|-c�گ���2�������f�' ,������X���9W�!����6���|����C�����QA�B�:#���{7#?P����)�M�%�&�?����E������bo��ʟ|-.�BtT�?~w���)����Ä����>��g�0��J;�Fz-��>�dC5�g�̗tb��m� ǎ���!�8�i��0κ�{R
8��g:����3n����#A��,����:�@��ˤ:2�������X����c��a��|���t*9,���W=I�7��^5�Y>[=z\�C��*GF�C�i9x aCĎ����1m����>�b!��S��,D���h�I1�y�0�E�J�a�F<f��$�L�zť�x��;t�6����P��p��`gr�_�H^K��,i��V����D�		�v" eD�3Nә>{S^�]{�����"�+
{���6�ry���6���9X�.6\�����t$$]
u�n�I?�ŗDAYR*$+��ϫ��:y ����D��QG��\m�@#Ɉ�U���D�	QʼQ2�3����}�IZ>n8�`��Y'�ů��%|�/U�(`,�� ��?����Q�>9���kSO��L��?$<��y}��E$���[�D�QƧ\@1n*=�����W[@ƣ��8�+���4uh!f��i)��D=[�MJ3z�T�V�BcW$Ɍ��|��ޤ�������5I��|%�+΄7R��BRzT+cX�l�|��z����QB�`��e��$;�Vy���q��?.��=�Ź��K��Ɯ?��*�W��B�ʰI��4�np�&v^��=�g���;��l��\���w���f���rhL�v�a�1	�[�K޲v�adx��u��@*|Ր��R�* �Ȱk˭�����l�n�"F����t�<��zN���3=�Z�u�1#�2����hr�������0E��T�Tނ��M^z�b��>����G���M����-��i;lߪa^���V�;6���9i���w�@����C���_J<~���[8�M��*/Lȷ�*S��w�u�?Y����=P	#J��fY�������O�w޾�7�Vʠ�D8x�Uv��{���GxQ���iBH-.H�`j��^͑/1~S��*�[,Vk\�-%��4A3ERd����
�}�(��<a�t �ߧ��	�T���J��'� ����;����&?@�/o^�� �+��u����U���Ff��&~AݹhP6�h�-49�|r�@�dt;v)��ߢ	�T�F�7��V�ӡ�;��&^���{�j�=��㔉��]/�h��gl_;2�d�/M۶��bS'���u��� #P���(V���a��p���܁Z��g*X Ё�lӊC�ǉ	yШK����%	i��;�|v0��O�<&�؇)�2If\O���j���a)5�R���k�9D70��?
���"ױ���"�� �8���r����a�m!�k\?�ͳ��P��CP��q�+2ͤ\o��������E *�\R.�y��b��؇������_7�0a;��������e��z�K�1?�r����'��@�c~������$в�:��Ks�ri-��UC���V�Y��m��	a|�bs	�����Q�������ޱ�d�_x�9��49���M�w���t�#ݢ\�(����`oP~�(�%t��ȵ�:V!n*��gH$g����Τ�I�t�a �\�vw6��e�Q�zc�F
ԝ+��r���(�-�F6�E��sF�#��k�ǿ���=��Ja�4�v�F���Y[l�ݘ
�,����to���y� ��$�,��������V�s.g�C�ۿs���Y��`�W?s��4o��)ʻ�9� ��O��v�/�@sF�'�*lC��}�`�g�p'�^6�(��FD	��zjK�j�P^8����?��B���f	*O��2�w�i� ]1P�2�qP�U�=75��P�8}	e�-��ޠ���9�h9
�دE�p���_���s��A	�u ��^�Z�Y�Ü���!V �t���1,��'�F���s�'���cD���4��t/�6x{��0��O4��f�a�^�		��A���#��8T 3��7�(��l�~9�3�1�������B�Җ��Ǯ_h��VEǡq4��F�NM�	�oEe��%wT�@�"�F�Ȯ�]�qzz�8�6䛐�ۉ*�Π��%�To�0�i+uD>l�KSO���iF@�+�~Vu7��2q��>U��#�)�G�#H(g���;��E���a��`M޲
Vf�c�'%i����z���J�L&�`t�뫹�]~PKD��4M���x�=W��K�4܂��)dJ�x@#�PO�9mD�4K�S	d� �i�cɎ�=�x��J�0�6�Ҭ�M1��w2�8%n��N�I�ʢ����sJ�0�"2�ݑ����� ����x$��-��AL���Ĉ4�Tn�9���hbֈ�#[P��3�) ���A&g��w�o�@&�u������&���<�I�Ku�)���O�F�d-
?��c�1	?6�v�9��uF�Xq��b��f^m���S�A(Y��,Kw�o"�ӼrB7[��WBE'�w�%��t�� ��&���8��C����dL�����1"DR��F�y��X戌+�w|n��jZ���y���� R�:���'y5ߟh%0�`N~PtJ�0�"��j������pG3����/�̣]�*�� ���������bR�_f�b�;f��eӗ����Q��wO'"B��Y�Ʒʑ�A���>Kz�>8�a6�P`��	j�}�FVA��a;P]RgS�b���U�! �M�+�����pX)
r������p
^ۈؾ
���c��tMC�� �.�W�g��5�F[B�������q$����I���D���*SU!�d�ѡ��}x�om9�,_�q�p(��q�����"v<���$���[d��B&�ȇ�	�ջ�_�<M��A�g*��J��Y���1���q�
��J�O�0�����;R�w��%0v��P��q�|��є�s���N2�:ye��[mG��01B?V�~J:Ӧ�q�z�h|7|Qq�7aЇ�sM��.R:���I셏���
;�_j�3Y'�N�sG������G:s����Ɵ�n_*#����@G�:�i!N(G�o�5�N���b�h���-����Cq�W1�t �8��=�tF6j��z!lt��Kr�����A�Ã�u�0��dq6(��E�j����t+	��2�FJEy�9���0F%��E=$��q���)���j1�~״��&��]�o���I��N��~#�w��M�^�������DW�(o�3雙IT~�_%*�����Q.A��$ �Xi�7��uf{�X�����xp0k!:���,���Fr������"�BBx���){:o��q:bm�������j�	�t-_��s&��Qi'6b!�yk�y�ӫL�xt��+��ߌ��3�P�*�Gڸ@aErF*e$߻�M!�߀
�fUg-�G#L��C�2��6}�. L�tO/��U=����Wn�,a�z<m5�{�S��+��j摇[�TlY���ӷ�!�[O�Y�n^9j�l���k���p��IlZ�(y��
��E��Ɛ,1j��Tz���u��(fͪ�o00J���L9�/F2�:K���߲�rj$@P�Er��Z�"���Xh���b�'g�f��}� �z����FDX�hN�T=�����)�*T���?  �P�G�m����K?���?m=�ȋ9D�-���k�v/����,}iQhZo}�!�]/;�+\��|ͽ��w�=׎bF�Jwls�rQ�I+.�
1��CSKaq�@��qu��\e�`�S�y��n�"%���)�=��H��w�2!���MF�{��T��E� A�N�����)i�s��������1�2������+��!&� ׉wN���쥾�o����޴4����O7P�Љ?w)�$� �m�%��4��_p���]l
~/:�4�Td���u.DiZ^ 1'˯ɼlBB;xn���C�_���VK�7:ᒌ&��>{�Һ����N��J�{�fZґ=fm�S���鄃�l��R��ܣ��%��T�3H��J�\C���Ը��$���L��X��B�^b	J}�/jȂ����r�YaH���@~�4Ϳ��R��yw]�0ͅ[���&v�Ya��6nT�qlC�����"o@1à�(&i�Y�0��+�J���oa4�2�Բ8
NJ|�ĴJa���+���'m��Pa?a*��U�^Z�^c����>��&S�|x�����y�ɋl3�G
M����Ъ�����ɘHl-��ch�e����'v��E[�9��tEe��&�y>|Ŧ�򌉕�{A2�]6M��s���:�S�$�0Q��꙾�Dq}�YGO��U#�]�J%~�K��4���\BH��IZ�6���K8�Y�t}����Ƶ�����o�,y�VZ~3>O�J�8�M�ܺ���#�i��B�~a����1A,ވ�(ky��I��O� O�PS�gfUQ>kۥ��@��ς���鯖��0�u�
��h�>��'aD5X=U�%����1�-���w|k� d��A��f��+����AGp`�ֳJ�E��p$4긹ÎPXڸW����֯�H�1�C�A�n~G������j��7�4�Ħ�������s9�7��ί�#�@G?)��ڲ�L<���ف�;�x/\%^����n�FZ��ɺ1(�f�CຝO5�Q�d}�a�8�}O��$K������,�B���'i����sSϟjgx�����_��9XX�ANT~���
�f�1�}�%�a
4�B���V�ʄM;���j�`����K��s�0˝�>G3gi�����4�(������{��	ų(.��fN�ޑ���Ok�����6�V�}H"-ŝ1TF��H6��u�_h��}��n��<6=�����$CW�΁�WuSG9�P�;�Ⱥ�}T�㩭�G�/q��SK(��0$�*�)���V�
!R���Ł1n!�x�u꿰t?��6IWj���i[���J��>T���ф�T�D@k'� �0���I�S��Y�-: �R�@0�ا�O�FN�6�[�pquH�l�,�}��Ծ�]%�"�f�~^����e�S���"�fk��-9,����S�d�+C��|�]K?��2�fG	(7�(V.��3�dɗ|~�0��VkSZhsHR�R�xS5����9:��^Q�FL�� V�1�WpLM�~�1���>����/TK2C�57��(y�װ��h���*N�|}@:6�Zt?��=^&h��nr���Δ�[X$�ȼ��
��Jw��ࢳWL�B&��)�j\0�į�P�j�\<���9�'��&��2��j��!�����'+I�x�H!DE���M�]aA��_�@i���pqw� �E�8��BnOӷLZ}�Ro߳+�B����$��w[I&V�Ne��6C�-1��o�+b`X�;�0���\��դ�O���m�F��#L����k���E��׌�u���这�]��m6_�r��nP#�����o���"����4<�*>\�ӯ.TN-<�M��[q�n|zd����S��"�-�ه>�_��������)h��J��vqa�gG]}:����*�՞�Lmk�����@i_2��Y-� ����`�:����c����ⴶ�Bi'������p��R*�������g>$o����NB����M%��Q��n�_J:��2�$��a�r��}1�v�
T����&/cӠH�C���!�a�z� �K�{�����xK�*��5w
��`�k/�PY��mO�:e���>;�.�o�	�KE��t��<��\%y��>� c#�	�υ��P�aX�΍m��v9�y��Z;���fm늮W���y���s)��>��+F����_nu+�(g)�ȥ�d˂��Ou&��TH�*�H���-IfI)v�4r��:E���`w'8�{]��˂<����R����o	L+��kbf���*|��Ei�4��<$��l����jz���w�-	+������ܧ�8\�o�P�c�/71���D� �4�E�]�� ���&vZj$��Ω������`\G���}���S~��
��cHqݜXC�l~���`���QZ�ݒ�����w3�2x� ���3pC�����������CX3��V���e[�(���|N\��za0���}��f^�3�T8���>-��B�wT��0���k�ˎ<��bQ`B5�ɀ����S���bs�32C�,���~Mg�l�����O�dj/���\�:�_��<�[�
]�xR��$Z�2����� ]��cՅ���Yjs2������׳�'�]��;8�)`�J0�8���ctr}ό���Lky��u����QѬ��j�h�T�8o���~���Ftբ��r��ϗ�W��׊ru��y��SxT�([d����Ķ��Nvĵcf�Uؙ�(ڽ�z�Iϣw���L�\J�
��L+&�h��<5(�HO�Ǟ��!t�#��DHM��A��;�,0�~�e�|B0��v��,]캶�\�-"�[{��ߜ��<��o\�$@y#�c�*1H3NQ����+%��"��>:t�T�H���0�+�M�(��Qi#Qi�(-�7�6���pC�b��4ї۬���.����-i~'Z#�/��o��~�Z)���1߯��y�j��"yJ�!Zfh`7��w�ܟ�(^���5Q�i�r��)�c�R6����@՛iB[��`�NaދD4��޿^�o3X�������.��8D R8�y<X4B�.�״����z�Ȳ� hC�$v�(�����w�����6Q���A�U0D�d���Ewax����Ȝ�%'�BC�ڻ��	}=�#I��R��=T��v`�l���/���݈��ؾ�Zz)�H��/��0�����GJ�ͣ����4%��[/ℹ�M�e����~T��T31��zX;\Z0g����Y�p����@�n�"��To�#�� �-�r	]�_�`f=K�&���;��="�;���L��ݾ�
D��n���ڭ�����<���H\=b�r����g?5�c9��z�p�dU��֭�z��"gX�cs��H������3�K�*f�J�=��\�S�A{k���L�y0�H1��5°�h����3Êp�І�� ���C�����g�w�^��e�B@7������Ҋ�
�n*�hϼ��2���y
}-���l�>"� ��ٱDk���L��U��O�
O�hޝP��^q��v��v�k}Z�e~�<C�L��9�9{'=5�����'����H�O/K}�A��9�/~�dY���{��p�n�IC�//�Q�鹺|����b�E����䩶��0K�蜣���gtGB�HXn5�6U�T�&7�{x����R�T��V�_�au�|�b��{��t�E�<
�T�]F�՟@��XD���/�{���9	9��ͨ��ҕOt���( g*�Ȳ멢4��
�:=����b(�ˍ�O��������kD�Ϗ�����U����8�GR�f׊T��;~-��q<���k�c��1Q��]�V,���>Mo�b��H�[�A�l�M�
A� �.n>Ӫ�cX�����	-	lj��rݜ/����R�o�E� �oӳ��Ʊ��Z:1�%�d|���l�����y�������r�.�>�N�?$� ��PɃ 9֨*dX���0�͹��� ��� ��a�#!��ҔI���y�N�E����e�C0R�Y��ּ��� ^D�m]��=?l�j�B
��Q�}"G����i$�X*�v�Ns����[x~.[x�aV�j����y���˟ĦY�b�d�� �6@W1�ژY+��?�T����uOUC����AcCI�5f_m����&vJ���^�<�ltBq�ӄ��j��h���s�3�*_la3q1�,�������:��!�
f�W���nD���������jl�cS�|^A1���彎��Ja�"��Rʊ�xՋ���i���F7L��Nþ��sr�����L����y���h�����rc�����O`h�c�q��T�F��,[8X�d�ȡ>���,%}iH%������',��T�+a�����1g�����b�1Ȼ5Mů6��i���	EN��k�G����M83j3	�?�>�t�*H���M*]���~;���5/�
 �5�4Q��M$�����:�>�&�N�1���Y�K}c�;�eN&?�YF˳G9��Vn8��C.����&H�X�!�4�缴j�K��@���8���K�a�'�7���s����T������NQ��E��@Ψ��_۲~�Ֆk�˲�>0A��J�h�k(���Wo���ZY�M�=�q�]�����_5��]���*\6�%g:Q�2�	E��#��'+9>`�����~=*h�^gD�XdwLN
4#��8c�cĊ����ku�x��j�ri�8�6/��V�R���BC@�~F{a��2��ka>N����!Z�k}Y���B[�$�#feڄ���_(��$h������n���dx?�+�j�W�PFJ��[�[��Q��qf)hf��j�k��흈��Ic!'�4���IN��oE9��cy� �1���;�Bx�����P6�-���jl/d�Ҭ<�� ,�~�����D�w�W������?�om� AI�Q"9W זl�����+/��"ik:�(�[������Ч*͘6�8�",VX+�#@�]ᚈA$�V,6�H��t.(�X��5l� �(�ԇ{.��e<g�qjPP�Ǹ:�#����Y�%��C���z�,F�s�S��髴dQZ��GK�U�k_�`8d5��ij�˥�Lø�:RN활� �O9>�����P�6,,�}j��i�W�3t1���#�1�sȻ 0�����B2td@��Ӡ��IV�����%�G�+��� ;��SY�x^;�R`�$�U��]L�PpZ���мG�鮯p?�s�����06�A*���q��B��9%�b����G��F1l�Я���t7^��U�8)��Xc(1g^��RO��#�/�G��w�&�
R��ï���;l�B%r����H����_2��S� �M]���$pq�D��s�#�4J�bO���ile�SwZCXm�p��<ET�!R�ۀJ0X<����,��))[�]$��C�&�?�Wz*���7o���O)v4*΄������bo�N�o���yy�Gܴ��Q�;�E��֊|�b8�D���k���E��A^�4�$��C��
h�y����l;x	]1�������2 A�|vTl���AI}.7�o8�f���,w��@�uFNIL���3�=[�/2e�3C�!D3�8�׬}G���l����3����ޫ>�9���i�N�.�����f��S��%�=��ms��v�\�@�ZŉS�%-�H�����s�$y���@{ˎ>�[��nY9�a�k w5�<�QB�C;Q>lZ��O�w�&h�~�0X�#��*�ld�B����F��+%E5�DP��m�.\-�n���ӽ�]3�0	�>F.̍x+�����ܕ���{���Hf ��m��$�K�p��;������lP;����%.�M�o�n�7֗˓n ��LcRh* }�y|�iK�da�I*�z�1__#?�jf�U)�f�QNg1j��.���`=����2T�� ۠Z�v�cwp_�<fK���Q�� �t�5o}]Cyc{sP�TE���U� ��C'�] ;��ա@md�ߤ��$>"%a~w"m�Ĉ�Qc��k���Zƛ�����C>-m��5N>nu�@�� �e�z/���,�㨢Q�_ey���y0ן�6���^�f���>5j�����t�@Jp��`H�$ ���1���N���]#�kb�sBB����2:�CU�k��,��M72h��F�H����W+���N?���Ǻ�����%"�5���ԟ�B2��mk��B�L;{4��v�UX�_(^X��)s4�J,�ᄫ0Kr�CI"�YL/'5�}�\dLi�iPv�D�E%����㰟�imԭ�����M0C�J�R��P�ct$�ߜ7��=Vk:f@�!Pn��2�5oT����Ε��hV3�����H
@Lx|T���<�'������<+^c�-��)��O|������6j���˭�b��/_��
��5׾�ש����,�'zM��j)G�Y�1��-i��4d�7~V�=��uΉ,�<컆E�����C�Q$��)M/`��|P��}����N�9�5�rD~�5r�V[i�3�d�X�<�$~�M�(Ȳ�u>˘��\P�cN�(�bX_a�)O����t2"��U-Jb�Z �/�§�������o2��%W�e�Mq�.�6I<F���%�u��'N3�:�(�dh����QS���q)C��%��yY��U�l�o:�BӶu�@J��4�,-Q�TU�Cl�mC�D����i�S�Hy���b���&i��g?81�^�'f�q.���ɯlQ�ߘ�!�2� <���K�Y!����-5@�r�|��4_�O��*�RW$ʜgkZpT���L�l���>d�īi��R}"U��;ϔ�?���G�+��;�~��`�ު���d�sݿ��Paa[��>����<������Q�S�!��	)!��Զ�D��r�D�2΃����.�G�;&�����B?� Q%	�q��Yc��	���{��q���Thl���);�)�އ�Ĉc[��C���� 1������m��J���).c	ln-��C��ض��:�ܽFr�M�A�k2�E{�f]�ơ���S����#Z��A7	S�M�FCF��`�#N���3��c�HJ�}�b{{U��k����!ڏ#Z�JI �:����`~8�䴮�8¯A��%�yY�D����k~t���������j���FO�����$���f	;�s�� ϴ�_�*�ܯ�����꾮���y`$	y�2���
Ģk +� �R�I�ۄ�,��f[�b/3U���6)Ox<L���W�c]����F�)c���ূZB����Q�'ț�ZM�<2m��t_��l��!�4��-�B�O�2ݿe��Ci�)w�K�L�m@�:ξ�3F# ��t4y��Ֆl}ɚ��������O�(&���1��oղ�]��Z���YYM�6iR3W��d��?�V���oGiwO�c�'"���}x���ڥ����ﴗʨ�J�(�-v���e��vmsb�=��=���xy�̱)�0Y-_kMxjQ;�xq�d�Fj_T՝�_�O�.�yA����/����}S��2����o�˓��9���$�'e�wwJgi۞�0��q���62���z�V��\#M�e�N�,��~ږ83���,Ti�ݭ[��xu�>�i��u��і��`��t(��zI��Ɩ���>�+���q�a�T���>(��'X�W��JA?�"HU�W!}��#��1��k�UL�/�xr�J�y�>�����0���{N0#ͧv��hF�"�ȼL�_=�Zۜ;"��/�(��}��n�S��"��4%��ѡ�8��7���Pj&�%�K��Y��Ikޜ}YB?T�א��`#mdI+��oZWf Ye*�?������|��_�#���l<Р�������ѧsh�S�ñw�fB2j>Un%��H`�!��R������=	�ߚѭ.;�H&��z_�'��� ����u�yN��-WRV���#Z�/`Knp~�~�];Ru�*�R�[` -�L�yg �|�Ey��_����[���c
�"����陦0��Ȼ�O��Fm�q{�O��x3�՟t�G��^� �l���Z�^%εT%;�b��[���5�.jF*W�p��� �g_lf��2@��ΨGT	@8
ܕE�v/˿3�K�yn��B�P�PB><�����J-=:��re�H9�>�_�1) �jO��i�L�{�<�B*�����@���҇��t\q^��*�|,�st�ɠ�92v��rUD�IG��k��3��C�5�����սk�l�s�ȗ�e���uqǱұ@�|�#F��q{�L7Y@�Olxr$���`��xG�K�V;�.�X%���թ��lϜj����ɢ�ց�\Q�lE?J�̢�?�kc��h�*Z(',k��I�3��� �˿uƐ���B!��7s����o⭻�u������w��g.Եj"��FG��D�&�.CIX؛��S�5F+n��kϫ��B�B0�Q^�����;�6�*���W���YƖr�2-��7���C�`��9׉S�=��,�ϸ���[.��b^0tp�@8�~�G�9���q�R:1l[�`s�R+
�io|���L>wʔX&ʂ�Гϯ�n�ƿ��MfH�a��Uo8��Po�ݢ~�	�i�����vb��<���\�m�A�[)�BB�l"�	��ԙ�+z���M���2�ތ"}��G}F`@��:c}P�f/���F�_\��|j��{����ˡŰ�4K#� ������5n6=�����4yBY{��鏭�|ؼ�T��S��1�#���e�Q̮R��7�M��B�C�k����)+�a {�B�h���	��ֽX �R��Y��~/6)�4$�ג�x�R�(���0dg��#A�I�Ye��B�u�����{6�ڣO�gܒnh�e����%J�Gm�2�����r�j�bWQq�^�s��^�����s�VUԳ	����ϙBm��&�����	�_Ƌ�$�|����ZC{	��j�.7 �<3f��X�5�[=�|�r��P�NE4v�U����Ca����n����Z�i��gN��;E�\R6.��>�w��s+V�Gk���5<3������{9L+��3'<H�X�7$Y�I[�)Q]T�MʎO�/�	(�x-OM��3���]����� a���|Yu;]�$���ЂF�������h�	�.rh�Z�w��,yb�裞8�]S�٧�wE��@j[K"����6��ʿs��~k��>����F�,H\p���ܶ�	���*Ͻb���ׯ�ȏZ��o���Of�*9J��Iº���H�x�s^����蓗ӡ�]Y�XP��w���'\����d����9���	�b���F+���:f��fR�r��P�vjO�&�P�/\�[g�G���zy>�Q1'h2�iľ%��o�'�z=�e	L}'57��-�����a��E�����r%���{~���D��]eK����^��dz�4J�BB��bV�;!A��@��ӥ;�u�g4D$1k*ɒz)���Aά!PrX�ϑ�6u�̤w+2 �!�Z�&��z<t3�}KP;�iX�(krȭ#���j��M��A�*f�����K)�(��=�|V!q�t��B��y��De\� Y9��۟D*M[���
��MP��}���^�kD��v#�Z�Fn�F)L��zl�C!vJ�v�ۭU/�[�J5��3�>������>����CH�Xw<�{{M�o��Z��߂�����̪�Qͻ8��l�=�|�8u�-N����b%��.�dkL�5�p���)w05��J�6�����T�M����k��(eUo���ˬz���C7�U2>.{�č+��{�mX�"&��:nt�!���;��(�4h?q���Y��
�9kjt���T�>�ȤE��*;8� |�j��a��l
�Y"gC���K�"ZH!K,���G_�,Za��Y������/唧�HtL%%=��GTaͼ�p#+/�� 4(�19�!i^0L7P�'�g�C$�9?�
��e��v�[F��(�`u��w>!arm�;���Y���ġ�S��,{=k��t7d��bi�L��n�r�|�f(ֈ�PrI�ĺ��� e���;�'��ߨ��󠡚# 2B"�w\�+�nT�.���|�?te{M"N��^ ��MM�Ue��1ӑ��P���pEj�I)�?� #e�$U��V�K���s)D���s�7�{��%L$�iYJ���b����]��'��z&�@�Rz��A�>q:s�%�����z_�V!a�F�Oe�tV9)#��-�c�Pɧ�!w�Ӟ��͝���@wP��])���;e�������۴�����mzoz琛�m��t���K0\]�&ʢ���!Ig���7� I;;W?�%Xm�	�Q%D�(@��k�)���Ǩ�A�B���}����X��H��t#'mnH�</��6�'e^�����~��Иj�lF5< ����wFDk����N8Z��d��mDr1ù&ڳR,�r�)����M��ڳ I!�������N�6�
q|�1;N��%)�$
�N�}�z����(hB�� �d���#	1��ۧ�������Vy�J���kg��ө|%#v:���x&��������h�����4R��0�qT���?���#��j=��.��וDR��ֻ.nm�b��u�s�t��C�.��������-ۿ�<w�Q��ep7��˰�e�5qg3Ub镂���?@p<Cg��1�3�!�X����6��|(�!��+v��v���t���2nF�>���0ܛ���3�����y9�+�����Ѱ�b��S�O�i�G�����}��V�̞�/�5�x0�b'���{I��\�\���CS��B�����<E�/z"�+KL����S#��S������D*�Nt3@��i�J;�^���W#���y`>�t#x_"hx�Q;K�l뽋X�0q������OU������H<q�^�#�K7�Z���,��.X�� _1?�?� �W�$���T�m�J�E��,�g��i�s y##Q��Yõ	��3n��!��/mፁ��ob�� �9���]5g�5*)7-���*#��C��J��S�$�1���^�����ce�(����C�#��V`�*�r����{�a�^T?�1ۗszȱ�0ۆ�r�NC`���߽u㥞���θ�^�o|G���Z��6��Q�(�袷X�:9ʱ�4E�zS>�YPE<��z�W54��
+T�پj�wy�di�K}��C��F+��D��d��d3<��	}CCji���v��M�A�%�ټ�_�� Q����x?���3�e�(���>f��?˱7��
�Y��?���t�,�9l�^�. <�jQ��h���$Y@5}�O�� ?{FB����E��+ȵ��ݲg�&p"*w-�S��e���:Y�z��W��/K����i1���6�������5@J���ݢTpt c�Zy��/������mb/�Xf�$躱��X6o��1X�M�ۨR��C��?؝`L��&�~*Z�Ѽ+s�ͺ�ll�Q=g3â���U�}���m�CxS��˝\{^G׋RNq�(�~��s���g�S%�N�XoOB+iU�o�߲I�_���U�ʢ<���5�(�����h�9Д~�]I2����b)3�����V�T������~�!Kv���]!��m�3�y�J�G8�d���t�@�U�}y:v�����s�Vx21�gu�lRݾ}&]��5e�L��(M#A�R��|�`�8���}����3���ﰛs�+'_�K�%��?��������ʶ�G�s�ȶ�A�G@P^�L�i����t���89�/����b�
7R{\�i�k�y���R��$�:_b��i�T��V�Y�f�h��U�	F�&(�x��c�0Cc7~�Æ����lĈ�O�N����vi����c��#)�k��p�/b~U�ѣU#GUA��G������j�n���%��Э��h�x���a*5�,ӫZ����1�߫�$�e���[�]�S�M9�%���J�q�[�iO+e�!v���ԇ���;�����rl���bIҹB��^Ӆ��D�k-��Dݞ�
ɑc��r�(�/l�+F�Դ*e�h['i���e˽Vu��(OmG�D��har�d+�2���������!?���1f	G�����)���yS�R�F���"l���d�ˉ��^�"�6�Ģqt$kx�hn<բ��B�K�
̉��r%;�癳�s�B���{�J8��sP~�8�� �~��K��@�����D������V-T)t��
����,�j	�"�\�8�Nm�=���ڌVjҟ�$�7������;�kX��Y��gb�����齶xn�E�v`"�6�z-L�U��v��T������P>Ү�M���e�,�C�&5�{\��-�/�=?��(��9~��?����X*BQx-�;6W�Hә�K�==||���tl�/�	8-a&۞,M$��ñ����N�������x���9�Kc5�d��Ͳ1˽a��8�R3V�-��!���ƀRp�T�pc����b|<N�8��$����h�V:�@�$m��u�ji���!G��a��V
�'aU#@r���j������K�� �*�Wiv�����ر�	�� Q��\OBҿ_�%A\��U�;z_�(D<;?
���5b����ّP&���XOV�fܞ_K��O" 3��Qx���<�̞���zH��3Ĭ�k��{wX�V���h��CF���1;�{�C�%��L'��Ahd�^i
R�-�T�e"[���z��"��h1اKG��D�ּ��SvMU�?�Λh1@���3�Xt���ڧ��}�IqV�8ʁ�u���M{��5x�F�aQt�ef�3>WW�6we���ǻ�_=L��wr��Nɀ��R�>�M�îo�%n����t[�i^v��>�Pؘ��R�Fk��d�4ېEgu#��b������O��`o��vb���o�	�����q�"��$��]-AP�!pi�_�1�2�M�Ȕ��'|owz�G�s5W��� #� �HHc����
L?��(� �b!��)΁A�J�۽��$����7�h{TV�)"���a��s*R/DYƇ,�Y�z`�A�O'����$#i���}�~���t���� x�+�;r\ra��E��g�E�76�ꖙIY��ptnw#}ڗ�8/,N�$�Rq;9�¾���3Y���"B8"V���OG���S����h`�ZDe�CRB� �T��@��1�a.
�9�[U�3�^���o�7o�'-(���|�A��M� Ӹ�s�4K屨�w�k�S��&d��S$/��L�~�U��v~=���[���sC_�X�A���.<[9|G3��y��}�bEb��PR��%��y1��h���Dk#��m��̖&~��*���>sƘQ a ��1�@BB���oW��_���s/W�L�2*���	R�J� �ꎜM~�M�'�#����H#�$�m<��"vSZS$_�#l Q�+�R2�AsLhY��sM�#3�7^�zU4�"���y�.-ɰ�[�f{g���K(�aυ �`W�6
��=0X_ᙫ� yD^����
�
] Ƚ���Մ��}ӂ���h��Se�Ht>IO��U�ɯµ���b��(���\��L �ʊb����dJ��,������R\���ȿ��cb)�.}��+��o�u�JN�O��J}��F�����o�\�>+I\P�G=�jm��?x%á���+N2�ڿs���)�P|̃{����A��|���.ov��I]�D����~^��g�u~9��}��t�skv�N������b��6S%4׻�@����%�~��ӎ��=qv:�5Lܣ�����N�]#�x�`hɐ���G}>Z��]�(Y�Bv�J���%�UG`�Z�|�?ڣ�=��w!��d	tdYB�D���H\�5AJ3�{��Ո��U�۫G`jGY�4:���.{����)����v&�*�>o��86o�\���1}�f�1k�� �82�Z�zj`vۖ�'�A��@�i�!,�Q�P������*=R��ƾA���=v]T%��t�be�/*n�%Mƚ�{�ժ�C�t�ċ�f^�	J��D������Y��#��`z��]�D����	��s��9#�s�C$����(˺Y��y���6�J����SF�!���"}�b�<��Kv��K��~Iۖy}�qsxGD�v"��lO�_�J�귅P�3�L�~�w{q�7�	����9r9���1AU��Ppr�p`�I�W}�ܛ���hߧ��q�]Vn���a����iGo@֘����)C���H�����܄����k
�P�a��U|3��|��ͨ�R� W��Y��r�3O�&��Ұ ]�L�����F��QH1l���\I��4�����`]������\G_�7��P���Sئ&��N(�y�)G[��b�)c�a�5����r\+�,��!�oZO_��.��@��U]z���&N^��u��D�Ex�v�z��2���e^J�vF�N6�C6�����Q6���(�yf+�֢�|� ��	�y&ۆ1������]���
�p�����x>�aX�K��'�s"ұ�"i����U(���8����ʾc*#MD����8N)+�����"r�5���.�B|��Û�ڣ%Y{Fdv��"-�� ���rB�
� ��=��xP0'�urL�=f=u�N��W\-�6����v��J§�c��S��Sv/=�tE�E�נ�3eս���0���X�_��e+C,�2�5#�NRp��Ke���jm�s����#���Z�+�re�H����Ӱ�vF�w�`�A@۫�<���S4�iL��6��C���`�߈Y>���a_C<
����$gZU�YN�� M*�߳v��QDn�S~��C��G�" *,qKQ����侐�PR�ln�ۀl�Dl�k���o�����l������S(T@�u��?F��w5�#������#=�%V�,��� @T�J������X�k3�Fn���^+
�4�&��>4y���v)������l�=��M	�l^�L$yE�:����u�`|��FC� 4�$�8h2��>���0�%��/��j����퓂��3�ڈPQ���Q���!α)�Il�\|���\"3=�k^Y��"C6@��}��.f���� �x-�h%�Oʎ��sV�_]jo���z�]���$
�VR�	>!�G���_z
k�g��G��Т��y�[�n�`չ�V�]X�y�������vʹ1�C��H�T��|`���;{lr�z�f0������5qlإ���|�t�c�5�	yR-�C��2R�]��e��Y�>1/Wn��>���R�:|��F�P�~�ĝțat�;�im7s1��⃌ӓZ'�8�8������ނ\��������~:unX��s�Ky�b;�$�U�L��Jiq+����T)Bva�O�N�[�cn�qy��݄O|d}Z�fk��<Fy��*��R����,=�r?��Y�q�����,�%.0ߪ6x't�Z&��r%�Uj@�#4^Zn�W`��ϸ�g�������1���bCy2^-ڡ2y.�v�Q��6��5C2Ϭ�|�p��z��r�Ne��`}=_�` �H�TS��������	P��e���b�`t���S(���E�G����\�V�h��+�<ѓ�=�tyH��Ѧe��2�n -��M��-`T#��ɛs u�R�i�&��[�b�`Al�s�Z�����C����s4�ܠ<��o$����r7��7ĎN��̧��{X^*�n��č�\V��-���K�ԖZy���ǧ�3"���;i�������
�uWJx�'C0��e{ЈV�Q���W"�&TR���M�s堃��E]����?���BH�.��Ƥ��V��-Ql��?�����/�wx<��;�'R�d�	B����B˧0:�'����9{"?�9m�ml"�X���,!��t<n�wq*� =�X��7
B<o�]
ZIRc��3Z�c�H����χ�ީ.A}ܗ�>��eO�DF0�@�Mٮ4�A��:�������kC����X5�w�Ac���ŗ�9\��e�}��;뗻 ��l<j�σ>)��A��D��Ne���)}ͷ��}}�7(q~��Z·nV4Q�XL��%�!��"�|+4h������L�W��E� �ǫH�fQ�i�\teȂƜ��%��-O�W�̃o��V����so���q	�E��]Ƭ�%�P g~�u��@��;���f�hpΙ���#�P����niP�h$�G�Y'��#��kd-��A ����5E��O&���R���Z�p�v���Ԙ�0}H��ͻ�X#�8�pU�c��O��lGÌ�QVz����o᧮@�nКxE<KT��3�~P�]�m�db8K��o�r�3�j�C����p��K+�Ds�-.�2N��T�%��n���S����̣+��#zv�p�L�S'�u����qΤ�Ԡ��s���Ou�\�Y)���
���9��Up�fJE_�Lf�R�^��+�1ȤwM�Q�v�V���|ރ<z\��[a�(G8�œN��� J�z�:�KX>MOة�B�I��o�~�FT�AoI�*���Z+tlݼ3H�3A߆�ܣL�rS07������ �v�}��˶�m�Tܭ��;�l�n�� ƺ�n��C�㧎�}q�s8�I�܈��>���������n��#§���� �3�8���$ �FAlW%ata٫d�i3��U�S'��7��,~�}���s%�+��	��{�5�U3�'��H'َB������_2���HTԤ�4�LAD��U,�(��D�����_����C�S�rH� ���æ����8�C�>�=^�N�PFAd�p���+2�Ӛ8nb]v�Ub(�À�2p����2�w �R�0O�@���|�ȐS��r��w���;�?�ʍ�
\�P\*L��_��}&��� |�P���&<�?�N��A������vq��>p����٩�����A*g(��eZ�e{�]K�e�_5��&��w�|���;�z�姀�5 ���PT�Z��Hu:T8����]sN�B�}���!��͢��N�,�܉�E�/$6�<xI��#�G��U��evi��ʝa�&E1=��L����2��H:���M�>�d�8�g��ՠ[>=�ˊ�����2@���^���J[̬��0�7ɨ������4���#�@sr��k�g�,$3"v\tX�q��M���iJ:�e���c�Sz?R<|fR�7'�`��Lu�~�G"N���w��xW�DD�pu�ދ�֡��3��L��V>Qx��)�O6'� ����0�	fo��j�$/0S.K�%�V @e=��P�/K+hy�&?<)�Np����UY����i7@���?;���N��{�d����c]�B����H�c����6ǫ�`n}k�M.�w��^�1��!����ۦ�8�Kl�zf���ו�c*��1p����s}�Ԗ���8g��1p�Z:y��:�M_��a�ʅ!Xl�̼PX�C)�����÷�Sf~O�\�c�S��'���Y.�+G�)Q�s��bd�p
b�`]!��R�}M	�6V������"Ku���Lq�Q�!kQzl4#�[DY�2��:���pܤ�0ì�K���H�h*vڊ�v�h���߾utI:�-)�#�g͋��*���*�<[��]?�ڠ]�w�$�5�B��Z���OJ��gp!�<�W�V4��U ��CK����i�%�>-v��*�����Ը��A<�[e��p�O��"N��j��U�~�&�̰�����߅D���*/`��E���#�	��Θ���U���cY�*z��F���Pe�5�}oq�wh�.�_W@��wˑ\HV,�{��(���A�	D^v -(Z1iQ����x�=W.�N������z]�ϗ��T3� �g):>갈P��b���R�؆�o0�`��S���Gx�",��;����oX�cO�E
���gZzڳ�Rm�K��R�[x��*�S����N �׏t��[N�Zq�Ȉ�.��.�7w��e8��Z�:�P������M�J�=���f.�h��ۦ<�֞ E��P��r��(��{�����Vӓ
��{�Z�	�X�X�N�l��HB���Z���n����<�p#����o��r�gUW���Is���H)3������0l��2q�����~�#_3?C
�;�(���R�����QiZ�;�t�8�w�/1jc5D���̪�.���6ڷ�?kT�/� =�%x�I�ׄN� Θv ��
3�[���vƓz�S��L�6�Z�D��(.�����fx�2�$�FP��=/�H{��Iy�S�����N�jO�
����Y�3J!�<k넘6��11�e����qfpQʎ3ݾ�7��@�� '�xm��mb�~yl�0&I�l��Ƈ,h�'�Z{���Mb���Ǌ�Ġ]���a���q@  �Sf�F�57��i�5)���%?Pp�?w�f���j��P�y� Ϊ�=(/Зǌf"�d}|�*�/�"�R�p]�ٟFl�zE֥�d�^�t#^�/h9�����ĸ�Q�NUfQ@Qv�gA�� ��^-�3�_⡠� �[CC�E�:��7x�� 06�t�	�M)���[��"��k|���sEd|�𐈃�KJ�|�^��D�����|��`��e��-�1hнC���ρ2��~�����3���ûr�"�#�rN*�.IC�~֎��PO�/���^�vsܡ�G�uO�(X�:�U�`�h�&ۃ�T]� ��0҆'��|kx5 z$�.���̣�L\˟�y�* �:�����~����,4��5	Bn��~M��{�(�ë�_S=���I&��2�NC�fG�^7yr���{{xד&�_c{�!��*�
.Kb�]P��AC�8a�p^*:l�<۟0������t�A�UU�ӝ���t��á������$;̵��Pq���O#Is>��Ē�[��dK�N7�;͘�����{?Me����~���`�AN�PmZ����`C��t�H93m���WK����MG�瞕�i��~���	(R!����$�_����,�:ya��K[�]�]���ȹ�����q[FV�c�@Rw��f.��F�T�����,�Qt,�^E�A�&��"T���)��}���֭Xyg��#eu^�����˶P�sq/KC̤��i)bK��>�Rѧ�,�R%�6��B��\_�����P�5��LU&6���'^2A� �����X��zn].�s-̈����9�F��sn! *�����ku��t�5p�,�Q�͘_qy�V�":m/��!3���%s�HuMBO 9Y�ʆ��� �_�@�o��5E.�n���m�=%#�cVM�6=	NȪ�M�N�l����a?o}N��=���7H�k�"�x�w��������~N�Z��+���-��H
0�W �#�J�ӤC� Tu��3u[uЕDDW*ڴ�� '��!lC�����+_ Q�V1��YY����=��͖0�o��F��\�<��L��P{��
*��ؽy����A�0��g�a�Uf������L�e�b��=�$|��zzD4��#���i�l#!��aq�'�;�"f���HJ��H �����9�Fo0�tb0���W.��t�A6K->G�nX�=*�n��o�����GJ����-i�ѫ�	�+��B�����v7�M{L0X��&2����	Ą�Q &ǎD8츚҉� �� ��2�Z72K����
��^8�I�$�0��#0Q�E���2*��=`	@��S�Ng���s>�A)U���R��	8s]��I����ס��?F�h�?­��pB޵S@
-"p��[���%���.�E-�4کѤ5@��7J���3r�	G���C�N�R�a�#��d��m�T�IJ�����E,�x�b�$��}���P�����$*+��##�Oۮ���=21٨AH��Qc�������ҁ�܇�qx��.Ru��ua�Y�%��5Qwm`dK����!-3"�h�� �F_��t�F;���s����̝��0�!����䠷�:����V�mr�;XTߡ��Y�\s�5���9/�'ęZ�L��F4�[}�:{y���V��mZ�D���.��V�B�׎���ތ���`W#�鄄��̃��tگ�'��349�MB�ex�t7]���Y��|��~C���T�c�E{.{Xp�:\b�y2]u1�� |���l*6�\-x��
=�C+yX&�c����/?t��]�f��^�_;�eP��'�C5�`/Ga�f���]��R����R Ҏ�cGA��j�
�	��4V�e��O
�W�襁�W|�ի[�C��= �Z��#ř>fD�$C�D�Z�|���(��̺������,(x���=%%ѝ��/��N[}�o�y�BBD�cϫΗ��k(��� B�`m���^e�O��|d	#*G�KIHŌ�~�QPJ�9Xy%K"�WH�7x��dr�i��+�۟IG�j7��Op��)��2��O�Ǒ���n+ֲl��N��b M&� 2��W�Vjbwٯ�����^,�.�^h��xR5#?pR��W�k !Zt����;z�nP��Y=۬䅭vL"��i���~��ɞ�^��p��u���?�w�Yi��P-�%�X�ag����^��$M�Zh9-�R�}��/��˨��@{�e-׺b���L�&(���v�mw�:`@	�q����h�(���-�U�X��"*'�%ڍa /�fT��\kFF0*��ȱ�$&�1y�,�Z���k�e���P1/1ٚ�ZE�D��S�G�����t+��'�yC~sPW�{�+��hP�v�l<���2�Z���bw��RɕJ����ex8�r:�����-��5C��g�#H;3Uk{8��W�I������u8���U�Ao?U6^5@ -�>��`�/�Ahf_
R%��x�	+�%f��{uЌ�2�����iC�����I�b�2g��A��o�I\s~=-.
��ͩ�H��8L��&�E�"���m��� i1(�"N^*Z߸Z���ƶ@��g���3^1`��:�ܼ����!\1���[�u�I|s
=����x�n�:aa�i V;k��z'����jWN�qM!�O2i �I�A�V2� T?�s�9�w��'ji�#Db�,�(�kB_�.�!ʔ��RY�l��y�'�oB�\��\�+Ȩ�vk��p���p��V/�c��W@j��#����P�1Tz���2���]��sBf,���T�E<�$���}Ȃ�C��3v�&R�XQ1o��Z,|�W&����2�?S�=�$1���E8���N6����Acb�:9k13�2+�c����ڋl�<-�(R����Q�ϭc����`�<a��B�c����� � �.͔��*4c�:����Pd-QDu;i\s��=�sh�Ol.b��� ������e�q�@�T�,�A*?�S;���d-���V�q�o�HWaM���9؃?�M��׫o�����]�<��Ԛ�<�#�-��޼7��$��t�C�Gr݅9A���Qw�|�Zׇ'��~<�!0�qq)�C��*Tܳ��*���m�i����7KF�
5�Krp�aF��.A�j��M�c�&�-\ʊ��P�bb�e�v�d�V᧖�Y*ye�y�p�	m�U	�^u{E��LGdLs��̬e��DU��)�
n3F��+Ҡ{@��(K��Cu�2	7��,�o03@o8��3wR��-�E�m�n���4�?�����WSY\��^�؝�ѻY���Gϲg>O6Z>Nx���X�D�ݦ��rvB;�ɕ��4�^-��-�C��+xg�mئ��Ӵ����@��\��tO"u>)\-�z@_��
�ݻJz����6�^��T��ŷ������'�9�Tx����JQ}��JTYBDB T��8�Q
6����C�p0\x"xdVO��*z;.2<f<.ɬsp�u���t��,iXӲ�"� �J�g��צ�ͳM����ݞ)���O�ɶm#��-�Bk�;Y<#�QK{�f��8�I��-Z@��w�Z��ԡa�pxz�ON?���8�u���1+�*��r��Q��{�������*"�5h���~�'�u�MO�U}�m�	��M�Ic���OC��#��R֣�|3RkPb�̹$83X���QB���xdc`zoi+]��l݉�j�1g�d��0�^���AB��?�ԉ[>��L��y-���˜e$,��^���p����ɲֈ0*��a��[�2l��L�.%&Ѕ����Q6��z��a�pWYZ(��&S�6�ۚZ����F��|(:�m]��2) �d��͙���A�C���M'G���-M.6�(&�:�d2Pv�>�F($�-�ww��K��cE�*�59����6%���\�� �}�4�w[�{U�k�`��[���Q�!�))	��B;Um���������yŁA����o �|�f}#�_���}~ǩ����o������E 'J�$��t�V�C�8E�a�x�A���%,m�_϶̑�$��eU
��<���B��&��6Ȏ0n�N �r�[2��{���W��Qa5��k���� ��r�V/��YG<�Dq�B���񬠣�������嫮���4��S6E�]��a�3><[n��
���>�Z9Lk%�Uٺ"�1��,wk� S�Xn�������Ʉ����6w��Z�R�2�`$�T5Y�1�$Rɑ�:����(�R��qO��0��g�,�K}M�#���,������&3§�#ӝd�~�)o)���}+�n��dw6	�p'�巧�L�$-)Mt��Y�Kq���9`�M����2P �D<3���D��M�0��PF;����S]g +�aQ,]Bby�t�ޖ��	ݔK��rs�$X6�����5:�C�n�da�N�,'�*���S�oexJ��|�Y~�����׿&�(�*|4r�Q�C>X�R�w,߼vܟ�Ձ�28�MO棍��%��� �m��v���Ƕu�g�N�OcB�zsgU��~��ӹ�F^��������!Xa����bV~���Z��c�f*0��!$�'6L�|��:o2�X×ྯ����|���mT���!h��Rә��s�Kf)�N��=�ߌ��U(�TΚ��Ϙf�cҏ\7�оh���ۣ�YJ�j�'��e�_"�2�??Z���^�~���a��:E�.	Ui��6��t�ԘeyȈTlM��+����dڿ(�����r��R�z@�.��6&W]F"x��y�s�Abos�
��!�i��A�x �����+�O�8۫`��kٶS��c�ڞMgG�vb
�&J<M��[�d,�88�Kw�D�����B ZΨjE�լb�nw/���E>�qmS�o��j�T����rHw8L�������԰ ��ɦc�
�ce�=�����V- �͎P#���`}m���Q5�4`�^���t�H�x�6@]�	u�*�5�o��k����)E���=�-����27��螕w<�5¤eut�6�����
���N��5&��	.�c\���m�&��:���9
	��}��m�I^r���<p)L�'�yR����$�X���I�����i$<�0}>A��tYK��b�8�\��o�4�3�2exR�~��=��I`���6-2��oo9>�N�l�E]f� �EPx'��ݘu4BK�@�\��W���>V��V�h��#�։ǋ�W��8��Y�`�T�-�ϞfLȫ�� ��F@C�PK��@�g&�:̩ɾ�/�����f�*'�@gs�Uhx��l�w,3(phv)���{v��̑ה�@f�j���"�Mw���n��U:|9_����4p|eշ8�}�0���mҎP��Wϕj7ѷ�R�]e�U�#�x��y�� �����j!# ��2�j�5sF)&�F�UiC82��2Ik<&�EnU�z�A�����4(�/��U����F�@��_��n�;)7W�J�ڒ�bB%��bm,j��˫���� �uܫ��s�CD�7qf@�1�3�.H�ɸP䟙~�>�*�H��Kg	�ܴ������F2u�w祲�N��0��06���a�y�0r��"�h_f�}�s^"����Us(ɿ���wq'*��5`�	;Gi�
x�ɳӉ݊�7S�`ǌ�����E9t~|n	_QX�~c�N�p�'q��0�y|W-��R�k���bp�ү<N�=�J��G�R�K=���ޗ)3���.�R��ğ�����=���B����z�Aڝ��A��T[����0����u�Uk#K!�p-D3,*�]�
��@�IQ�=�Cv�&�u_�n»#@̐��@�qR�\�Y(���-f�G�%\��( ���P8�; \<��*0=��mپ+�<љ2�Q���_�J�S�x`)�� ^�Ɣ��CU-F$��O�;�{�l�y���%$$�#��Q_��"���<����/�.46;��[-�'@��WB���%l-T�#���0v�^��l�|�7D��"�����Z�/�	�J����	�B���z�z ��$��p�t�m�P�*D����@��!�B�FU��uW��7�Y��BC񐚃k¿���eB��ށel(���:37�
\��{+}�J�盜����b���5q�l��Ѷ'���3GU*2�+j������P�����H{���"4��p)��0!c�%�������~�97���M��С�;�A��3���~��怈H�u�O\i��>}�Í�EJgXؚP�J�6���9��t9<'�t��\���JK��e�w��9��_��� R��p(Q�p�$L��R������>�sm9��W�9Q�P,3�2W�C����g��K�b"<0$H��/e��O$h��5�x.��1тB�����ָ�_}���΂35s�i���2De9;��X�	oR&�L�<�M͘�p{{�C�c��x�S��ޥi�?3cж�i�Yp�[��L4#�O���l�ܰf�<z����e;T��M%��k���㟷�Ā��z+1��z�)L�%KY*�����-Ȣ`�(I>��9?Rn�I� Ǩ���Y⏍�g�Ѥ3�Ú6
��IVi7|�Q��N���?�٣e!�}�"�����ɻ���T9G�&�u�l�V�K&8��m	�y�Cه�e0E�b�P���L����I��N�c<�!�ݢVov�B�iE'R����6�M���g-�Wm�itg�Wֶ��p��+�6N+��e��A$�����J�������so��z���'T{� ���_.o,GX��>F��U�uS�[�t��#I�-<����0��QZw�-�,�{X�j��YN�u�d�p��z:�o�� ׷�7��ٷ�kV	��᯦Y�?�}!ݕ���v�ߟ�hw	���R��x��\5gd��&��|��r2L/a���2w�����[��7��Q���Rl?/�g��+^�z+�Á�~w�md��nX��z��4^ݝ��t�	T oB�G�x����74掓��G�{U��iG��|wn��ĭf�[��^5А��-�Y��qBǗ`�n�+DO�Rѧ�g�v`9���aF�Z9��y�G�8x<�S�������rɁ����q3���TĠ#d	.��:_��	?�<8{K�~IE��I���������� �ԟ*���O0R	A@��iPX��!�余��e��͕����WK^�E���*�Yi>�@���;|��\Œ*���Ӭ˲[�!���L��T�I��05�^��d�P]�� ~m�N�ܷ�g&�(��_�N�:{OUi>�u�p#}����Y�2�!��<��k�/�w�`lȦT�΃�}�+\MO����Aw��qn-�5����ipq�X�\o�_���f"OK��뾧�\�$������#���ڬ{�!�Hoىl��3��]ܛ��7�*J"��]�6l�k��GX�}ް�h�r��]�b�l�;Zo���{p�L�I�����*����	���`�C��<�Sc��(��`F����x�+�OE	Ƽ�o��}h
*�}���p;�X�����[)����57� �\`+?���&����֐m�O�)'�k2f˂�o��D��qp��1�() @"��#�\⽩Ƥ/���R }F���	q�Mr������"6?ğ�ɫ�l�S���[e�2�m���0^Le�ID�����x\���&���� �ߨ���#�=�R��j��.,Ǽ��{�>�7��(��5�����@�Z�<�^e���ӿ��ıb����&O]'����'��T��K��"����2*n6A�O([���O�W��tـ��I�q|�B`��|@�,�w��3�b�m(��#򓌠�.���$��kM
��K0��?��61b�`�rة�L-�"����V7̑�0���Kl>�����߲�>q�`�Z݌�RK�}ʓ�Tj嶾���:���t	+NM���G�w׃�A z~x��^/�gU?�e��TG�� �%!ez�m"d��"�ь�J,ߕ���g����S3yP�W�X?�zt�P��#�1{"a��/̀8��� �{+�&Of
8HqY��t�ZrA��g���Q�=�X�gj���%)y�;�LlM��� �4���q�����3g���J��)]+��W����|>Py-c��>�5iQ¹�2����wI���(pj�S�G�<���tc*�xU�X����nTv\�gX[��G9Y���|4�RSz7�Y�����;�L�ȁ'c=�V%>6hP�u�R�mS���+���2�l��1,N�V�P(��0�9�+|���kVᤑ/q���msp��S�"E��.�{����8PGN��r�{�cLP?�P�Y��Zd�6SI6H���|5 ��vb�YsQ居�+7�?y,L��U�E:�Oaܨ4.a��5��Z�:�k��K�|F.���dm�<�.�J��B oxSn��@��BCli�S:dN�9uƱC e�����{4��h�:�e!K>��ѿ��!���O�,���\k�s�*֬rVB�F%�.Og&>�no�0Z�૧A�Lq0A~��`Uz8����RJ��d)l�]�������gF��R��\{��e�X�Fe�6Wj����;Tc�ĜG�#�����٥S�U�����e~ܛL�:�
�@��Z�������@��4F����5%�lrV�J`�Ṛy<��e������t�4g����Z'��%!lue~˵¤��n�XG��Y��L
v$@=�\2%h{%/Q�̹}!=q��9��奻�� �_���sN �%�д ���G��,rI���W|�d����Je����W��z �-=7j� %��ଟէ@x���#!uz����IѬ����8�B��f���A�1n[�E񲀾ڌ��<8pF��fK���2s�)99�ӹ�������L�c�"s��u��!C&?h��ɪ2�<�3+D����y��-pw+�ͷ�-�/~�K8�r}�4j&m��B���ܱ��2.^�ӊ2�䨨d9���搻�R�?C|�,�U�JXŌɺu���n�PPXS�VjƗ�,�=��	63=g���~A���㇥�%�[z��܆�K�n4f��hH����q�[(,@�l�!��?��?�8�%ҩ�j�^�l���Z����M��'ٮ��B^��fg���o���tq�\'&K�X�l7�f�$�����y���L��)J�Jӧ���x<;e=N�",��U��E���u�:Ǧ�z�ѸO��OFD.<��}�? ��$��iй$���"�p+��܏4�]b��&�GH�Zsv�EnL�?#��ޱT��^�� 4t������ik�r���h��P9N�UC���$6�>�U�S
5�o�Qt���ҟ�]yQ��z����K�:�o�[s~�񑧞�H�	Rq���o^�����a�R�F"��rCjyz��R"5���$����V���<n�r0f8l�T�_ E��k��i�Ft�޷�@I��i��ȁ}���q�%�e��@��;Q��T7Ũ�k��\�QS�
۹�2��ȍ���JZe�L7ܶ"��E���M��L`�f����E�Td�EY�f�G����WZ�.�
��g'�=Υ��#pQΆ����u���������T��|��nʉ:R�"bzc<�e�Y���/�w�آ��Bs�̜A����{�7?jJ΅Rr��wN�����������|�2i�;�FgTR�lP.�1�V)�ưNf�[��ç��O��j�*�+	<Ax�\��\]��QUG
Ry�3?4��:B(�~����˷�['�E���`��PS��ر�������ϼ���&
ymt����b����	茔"�{[9J�� �o�DF��NAw�e˚R���;�g6�=m�hk���H<[)*`7����B«��G�Yi1
B��@;�抈gܪ�f�>TI��2TU���>�ST�j7����<���T�� ��`81��(@��3}ϰ�g�=82�Z,�/5w�>,:�0������q]�c�q���e�7�^W�8�W�h��D�vgބ�,���  m�B�:*`t��D�t�w��F��������g���.����!���ã�qr�a����\���YA9�m%���^��7Z�_C���H	h!JE�8|2��R�����`��/Mx�m����i�����<6� ,Ϸв�g8`�g
�"W���<�90�X�x���JUo�="��hX����R�w�?�Af�}D���=f�*Ũ����2������snk)�Ж��S�(:���'c��֟�t�zz,��%���8Ul&�>.�[4���1P��[	OV�e��E��@��oB��`?<���?l��,�;&�@Il;�{^���]�?Ĝ$'���n��:��A����� {!Z2�Uxߚ�O<�i��W�Iv�v|�n�Ղ~�`�fL��[�
�@|�0�m!fī-lz0c{c!�-�.js���Q	�/�ӗ�9]�Θۺ�����{�ȎH���i���-2��k ��7.�6%Y���'�~\E����k|�����(\\�7��R4{���
��C�4�S����d͵�oZr"}rQH{�Hi�JsldI%�Giُ��GR������i��/e@��ن�0������m( ل�l����i��I�"�<.�K_���fh������h^Em4_��r��aH_�(�T�|r��r-��(��]�?P�h�������~cڃ~d�Pp_���[�@)��?|'hS�8���q��X��C?$`�n97����J�yG��3����y͍�"d�kߌ'�n01DrU���nqt%GV��6`dw���s~a��Vd���LQ�*x�j��j� ��j���)G�Xo���rFD��
k��]���-�	쁊V5��x�2��B��%#�⎬�?�?�{���gyD_�h8��A���D]Q���{4�����W;���ba�����ڛ�K����lJy"���]���$��t��ެ�y+�D����'.ֿ^	��;�� -�\�k:&'�s�Q�H�]ܲ��M)l���r�s��'�Y�g�ye�Y�>�!Ū,���9UW	8u�q^��j�.S4�	l#�ˡ�^lF9�%�l\��=��!~w�浼��/�,�y�>JQ��4=�5N��`���/�D�1IXLA��)�Ԗ*(AL�[ni��	�1=��j��I /�e�4eu���}�7�����lԒ���vZ�oY���6���F%�\a�~=e@��u8��,�)v'k�/M|Ol���6/�8-(T9�Κ��D��O��	�$�=�ɲ����Vxy���\��d��ջ�Au 1���K}H���Yħ~�����0:n�! =+��*��N�b���ܖJ�ݵ}�J����a�Dc(_�c�����? ��P6=�V2����F��ߌ^�ŻͲOA�O��;Nt���dt@�P2�c��2H>�̞@>�M����c�D$'q ���ܐ�'x	���,r,�
� ��r3�/tRx9TY�qs��gM7oP�xy��ç�F�!�<ge��:��3K�_��q��Y`�K����mo��P�W��ʉ��E�s|�+z�1T��I0x� �7��Qt.�pڣ��w���\�+���wR}��g�T���H|ID��6�!�Ng!z����T�c��hM�bآ\a���']\������<�<.��l��I����C~h���r*ϛ������8�h��ĩ�&t�A�0����F���2��S�~ȟ��"ρ�G~���a�xQ�e�8��,q�{I�s�E�98�Xڠ�)]V'qNg�K�"�VkCVo�+��KoĶ(��&Zo�,�?Ha�4�q>�����w �;^�+SW�D�v':�,�9>R/H��ʿ#�6Eq�^K���t� w*��,L �IQ�K_��bdp��O�����}5�;���˺lG�0�h!#*��fwJ�Y)"��h��
m��✿�^P�=��C(ɵ��%G�������X5����v�����eS7S�����[��4�E~�Y�l���uZ��ձ �n3�m(
���M�XhP�Q?iI�,�.nW���U�7�O��6��0�>6B�M�
ɮt��!�C%�ˁn��b��%{rSp� ���d�p����R̲_DPݍ0�txr-��j��1���_���A����2�?pѓZl�ɿ.%��1�w��P��#��Q}���0Ĝ�~-е��N�+�$K�i�C��7A��8{�`�������t?E�B�M�j�>�$�PB�$+�-5ɏ�F�!�l��<Z$���uE�|">*���th%�Mf�������ٸ�15p�����"M�u�Pςk�V�J������+�SK�׉3�`�ZA��&���#�J�r���$$b�fk҈�FA���[�ŵ�'p�o��$�Y�����c1$ГpB�Nu��0�_�^���A
Ձ��	&��`�9����ɲ���^��#�ǽ[�i*�G]�y��!�@�?���;�����ɉA�0���p7��pn�ي�6Z˻jᝥ��h<J䤸Vhg��!B���|���Wu��X�s(���6B���l�
|mM`�&������f*.pKu�������	�c���wj���G�u� 5���Ĕ=� ���C�s��Zu�Je�O*^K,Z*�!:��#��)�\'���zc�W�ڬ�Sߧ-�Ԯ�n}����2-��<���5�U��CCN�)���ڤBH~�9�b2բ����OėA�0&�$�d����@$��`?~�i�l�;f���l�{�?��U�[��j�D��7A��������xI���
����<Q�"p�#��/Ը�AyIy|�%�z9����ceG��:5|��XC�Z"�e�^�Qǩ�.Dpv�R̢٫��L��(�~���ޚ��a��Pe�4��^���{������>�L�o�I��+�q���ߴBM&H�õ���pϸJ9䔢_��h�\S�]ss�ok��W5CX���'(5Đ�F5�ߖM�zT��CNNu�8{7V�~�E�$g�P6�t�t�	G� �.�;B��J����e63�ە��n���f!����Q��B���h�Kt��; =��Ѧ֡���Sc<;�w��I&2W�=	l^3��@.Q�[r}��Lr-ǐu��S;��"Om�1��!�
Q�m��9$�:j��J����l��`%ְ������W�2s��
�������V��6+� A�G�H1��u����m}�f9�	>a��O�X)/)4ֽ߇��]�.�q��2��b�3(����y�ԣtr�f�
�U��D=K�zY�}r+���`D��H'��:������9N~�y���K�0u��%m�@O�v�n�Q3A�]v&=��*�$���;��1��m�N�X�<�0v9�sߙ!�v��hw�����(�̨����3�?7f��͞4�S�j}�
�����nTĐG�n?՘<@���ƴ��l�v���m�je������$�(���Ԣj+81�ŋ(�l`�n����8�
��r��hC�^�vo�2���" ɣ�����O]��ܾ4��w�mǷ�~b�|Q�*��]��A��Y�D�뺟0[-�t|'���$r�ќ��j����g.��ض���^�-�� S���8J2k��k���Ѓ*��i8KI�� ;�:�af�0�%c�M�� L��Y&��S*�������1&�uG_�9n��U�.>5���d����&����F�)��ؘ�_�[躰uh]�D��1�9�O+�<��N&f��3OE{�yk��8)����\Xu���yh�~ۤM+F���\���V��Z3�P��@N�����!WbF7�� Nvö,Y�3|d��;�$%���M�	g0��D�7��/���ۈA����zf(�!R8�~�Mx�w�w��UmN➻X�,��0#z?/�̶����j�*A7V栲�G��O�R"NV.��+f_�M���3����݂�?��u'��:�L�T��ѱ�'_71��i�z�)��7���-��.sW�o�L��f��lЦ�b��4���0w�.վhm���%�f�5a0v_�W��^��΄ ��ӵ���Y=��T�ɧAo`����ʻ
:k�A��P�B��!�y�K��X�8��r��*��}V�iRk*���ҿ��3nji�(䀸�����\�9��GY��fZۇ�s�dPE�q�@.��x#�~n�����=m�_�S}.��?��}z���#@��0Un��.c����yiέ����Ҷ�k41c=J�3�(rY>^؄_[������B��M0)��SO>�»��HΞ�pY�,Q��M�2fx-OLd>J��ѦoUK #R� �Tg*�m��.��Y��Q���O��'���
L�CM�ׄ�W�KK�NP}�����q�|��אJ�mvp�����^��EED7j���R�����deW:,�y.�"�_ej�F���'�"^ׅ��=[v9	��Ô#.+���fܸ�Tч��S�à���d&	����{X�$%�.k��qPu��q��>�&ȼ��r3YB�`٫�W	=uړ�d�1H���L?��6v�su�M�WB��u�t������>���o2��bёQP��Wa��2���lRS��֘�4��nI�Rx�� ����������Z�JҦlFs�*��rF}� Y��(�F�V_t�p�5�0�~�4~������������D鷶a�|�Ն� ��ڤ���y٢ޕ�\q�3Z#� '�"�Ӛ^-k&dF�]��%�x'ڊ]Ɔ�蟜�{@Ӆ�wG:5Q��N�ɨG�ھ����\C�_����Rܰ{�G@��$�/���\�Bbz�Xd)�0�1��M��1#�"U��mǯ��M�X�n�/'$�\L�6�m t����aӐ����)���]�ze]�s`R��hYB��.'`u�*~_\3[�$_���%����9���B��U��lS�Q+�b���J��2�{I�BwrK��
0Lrj�z�`�����'�[i��U����M~g��0 M���H{b�����7�u3�r0Ptq��^���S���` �p0!2��@ 4�3���I3�g_�D˵G�H?�P�3�nZ���r�{��	73c?��՛&7&��ߵ��>\��.XkʺG�g)���uTPHp)�_��j�Q��s,t�Q��NR���7[G\!�~�����cE(���M�}ݘ���8v<�zV9}��@pB�l�,�~��6�]�a�`����x�>G0(2��|��4��"G���RMi�>K�ρ�c�ל���Y��� ��;���)��� ��fL�!U2v3R*���s�)Z���ڬ���2"}�^�[�Ԑ��_?�	3{�y.vq��va�� BPo��m@�=d_��/�\yP6=�_A�l��gݛG,��1@Oã�I�9�1��9�?T��>>����ځ���?VØ�L(��{�~����I�4Ƈ�lmڡ?�̗U�Nr�U�#�hC��n��Y��r<R��"9� {q���%a}(��l@�1Z_�Y��>B)����\
�a½����1��S�[	,f�"m�[��N������AK������%H�S��|�T����^�2g(��?��u��#!�>_"����$�Vu���Ym���N�9�2�3x�k�?a��I�ot�$�c#	{��5JF�W6������,�_��w_I<[�n�-,(��f\�����*��^Ӱ+7�����f�im_�M�q������e���j2 �N}��n܉C��nۜz��̓�6��/��ME=R	�I�Zx�"bD_�i��R��kiك��	v�d�Ϲb�]�H:ω�0z�\�)Ȼ��R&��~�Z���ݾ@,zS_*�Kz�;]���e��uuT
�R;��	�!A&��±(�p�&q��B�2���9,	�Wu���<�"�lB� �����������'"o���/G��70x�a���)W�OX"���=ar�9��\����V�]a���������+g���}bD�,���];O�� M�A�2O'p\����-g*&��Rt��S�+Mc���Xe��p1f����:�%������Q�p#��ht2B�
��ǣsI��S�o���e�ä)
�Û���L>��IJ�:�x2^�H�г��q�n�aZ{�Lo�s�,���A=͂gC�Άj{��v�z\�Չ�����}�5?����&I)���iQ�y�8��ⓤD��������,����},��&@T(�P��4����pǨ4��'�	���kA(�@�b������yݨ��q�0d[k527S�|�+�E{=����8�K§E���fV >��gg�`�z��կ��%6�3!l���~/�ho�\��X�l��2��/����s<��ɸ�J߱���[bp5{�����<��"gl=n#��2�t��B�<��-j�&n��FR�0�V��2E�@{4��9+�I��!�e�C�
��8~�����J���P���ag5�2��൬n��)r=vd�[a"��,�q��P�a�q���P��?�����Ul�~��[��z��慑��>/F ���4�/�V-;bD���u��2�[_����߽vU�P;��Sɔ������8�=֤뙙5����8[�fUJ#f]��p�ɺ���h��0&\:^ە�$����G��XP����lF�,{��t�L�t��L�Mؒ8;آq �K!U��<�� 0��B��� {����F!�z�X�/M
،N������<G>��D�B����k��"M��ؚ��a|� Y,��f���ІIk���%\����`q�{��+UW���\�Ԑ�T��Š!m�:Ni�f��Z�+��`*�Ү_�S��i �Sqo����4+S!��}'�筲i�7*�Jp58�)�3��E�רD(L,g��Ճp�.t��+�큪�a��<���ȱ¬3y��S
>�+��27e�/NH��u�[:������q�u�;M����T�&i�4=rx�!R�]Qݞ���zWf�R=.g
w�_F� M'tLk
=����*tӜ�~N"Z���D��Sx�i�\�]z7FY�m<��5�J����QD�p�����_����dK��۱�o��8鎢������6�f��Qj�e�Fg�BGU~��S�����k>���5��y�4�!,x�|�R��g��h���@�F�x���>��m���Pr6D�t�����_��l`�v�4�r�2E�DخM���p0��C�����GP�j�\e�D����vU�p��a~i��etZJv=�d�~��р;ZE�����p�:��������T��偕9�2'�Y�ۧ�����ΰ��뛙��+����V�H��٬����okK4om�Y6����?o�Uq��6U�/��4#W�T��f;&�&.a)��Ob���@7�/�X#���D�7�L�ьǄYKW��K�v)������e�R�5�N���Bwd^�]��ͼK���\�E`��kgO�~�8������=�:9W�BH�t�ξڞpв�1�tf����$��*��R�W��]A)��T_.#����$�0��5�������0;��� ��gL�[?x���S�	�S�R��U���?k7��F.��ǲ	�"֐���z��[E
[y�
z�d�!��(�j��R:���ھHT	�61���/7�&2�[ �0�7
i*��|��	���I3���� c�\�^yL�����Ő�S���/U~!b�b������&wC�B�-m�o�K�w{Q������w����(�G\x.�s��q>b*�A�t��#Kqa�֯{����M��#.o��Jm�KBz����'ʲ5��Rm�hm(�CP�z�h�k�$���UyY?s5��~y��Vf�j�^[�'1�Z�$�������҅��9^5R[�;FZWt$��4�)P��f��[��ҋ�b����O{����A#ۋD�������n����Ƨ+��i<��mf	v��'?U�ǥ���8r�]���اD�k���^�C�`?#ob���������	�
��/���D��?�|&>��{�xQ�O%���JMEM�0���IE~5�Jÿd�؇��������Q$K��I�EU+u%�~^�^xG˫��D@��̳��$d#������^�&).�UZw&���.`��=�"��E��Ě9_sWҰ���.�+o�낡<5���B|`u ����ĕÊ {����<88r&��t[���4�@)x�=g���ĝ�YF�Qô��\���[���nzf�Ť&j��EPD�G���o�V�����2�Ù*���16ǻ0���}�2��R�ڒ�*�mp��'��p�����.��JIN;�(~-=56ȔAI@7:�u㎖�\�,Yc�����"�ɶ�%��C QRDts������oKe��ݬ~��Y|��k�J���X�|�F�%�G:!SZ��4b^�����2��6��=���BޖQ}��:#����u�qj�IqE)���b��I��?�z�M�圑�z�7As	%��l�ρŠ�>E��΄���������͝h"}�JT��ŵ��(13+��Ǘ@��	���k�����<{�a-��;Z��g�]w�z����t.I)�����B�)������_��L�B��ځ��/�L�#��D,T�Ƚ���a�
{w
{iN��!hG�{���!F��oa��y�u ]E�*3$Y�I������U�ζ�ި��MC̛�����"���OmD;+`�d	�=�ڐPWo��}=gZ>���ǟތ9ɧ��1@O�!9�Zo�,48�l%)y&ݎVu6\곀6qK��7�~T��m*/���9찯�J����� �ӥH�̱g��#�_�8�^LjV6/����6�K�+vs�p�rY���b�����3�3xo�9A9�Q�7�����M����,��Vm�B�\�#�#�xBKP</����}���D[t�Ŕ�3��N:(t���� �υ+k����N���E����˞�A7�h�X� ��>�j��w.���U���R�~�7�J,$�]�B'˥?|�r@��kP�~B���|<.+ /U�X�XѤJ(�jH��ҠI�=T�3=��y\�8q���Y�K�tn��1Ԣ��b�o��k�T��B�?`�ޏڃ�1BS^��SaXy�s
tb�!�CߤH��xrW�<l�^�����i���̨���~��G�Zw�. ������L����y
��d\+~�9uD� �������6u���Cs�첲M�G��3E��c��{!*�*�Qs�Ĕ��s���H�fy%K9��u8OeR6z?�kv��\@<���Ӝ)׭Y+���xE�9�I�9�`��^c��$ק�G\���%��p�O���3/�1�.���O��G��0����xT0r�E[���+n�e����[��C2�><�̉�{l�C�w���}N�|� �[����G�_�?���F��c�r
�ir�±Osc�m[@oR���g����@8Ӄ�m6g�S���6�YpDAߋ�O�U��1���٦)W1��_�{��XFDW�'�����'ia�lTO7/�"������F�;�j�Y^I�j#zD����ʪ$H<Έ��X�c�e�=�6i�t�J��,b�^�t�L�T�����I^� :+�������
���y�3(M��l�	�{h�Nz���U=0#_c}`��֗"������#��y�P��@����_���5y�/2���ə�hsH�M��۾tw��|��ȱ��+�4�Ԝ	�,B�:����,��8�sA��IU�O�:����k/R�-�+I��]��vC1���_�l0`�%^"'���p\(P*Gױ���~�?����o�D\[*&��% �\ܴv�YO�2�Xuؠ^\=D�����H�Kj�ꬆ�o�Ge�B�&����CA�h�S-��&��UMj:�F+6�Q5��۱�6d���u�5\h�d���#��C���}�"���Iѹ�&�)�Eҳ"�q?1����{���0�|��1�����C����:;�}�6���:^[󵣿bbߤJ���3~8�;���/����>�Kˁ��0���V�c�h���3 s&����˧�w��P�v\��X(#���~:�޿ې�4�&��F���c�񷒞�d~I��.��F�<�b3���u����'��$�Ғ�T��\dꞆ\��b?��k[�W�S%�gm̍�M��@��$�cQ^�PJ�r����E�1v�i��,Ei3��ɡS̞m�h�gkj�|Nq��H]��r?y�P
g�zG&��YiI��2w���ʯ(��8	��5W��	�����Ц�+�)�^���&������^�܅���5�a�+Z0ɀ�0w'�U�p^��:��rlb��[Ap9�!�@��^;X��R�i㍒��������Lc��n�^-��7�H�׮A������5�و3(�}�N.?7�e� �W�F����zHa�"Tp[R-й��B3��tpR���-�%Tڊ��� V��W)�S�q>�e�9���	����/�Ʌ� �D�
��1���K��<ǈ6k�e�wdD��kD�%?Lʔ��H?���oe�I���seN�7��Y��Y��*P�G�kOMKK����ݗ�'w^���+�IA��f�cᰁ
,������9l�c�1�X+�˅��m?��W�|mn��$��g�5ae��`3>��I1�n���U�.~��s4�S�Dn��f 笳����LY�@��1p ���kʏ4?��#��V�n�nF����*��_Cxr�5���9:H4J��5��V��"2�-h�<ڈ��o�L7���o;�z�/2=��+Ç�l,ͧ�� \8@j�#60e�d���fc��tN�Q�V�Hd |���Y�3��(vG�xvZ��.jm�s:�L;b�i���"�-T0� -�Pg#��_�O�\.t�:)u���0��e���Op��pv��)}�9�g9�-Ǵ��&�EU �Uh74����X�$xnvS���;���v�Ь�R.0h_U˲b@�{�����JlCH�"Z؎~��?��?�D�ZA� ����( �:~���(1���ICW�р��#�"�=���n�o��v��d�'c%O�����vڵ�>e ��B֕�b�t}�Yg����)yQ��+��5��+�aU*�Wo~޲��ϊz(�l��o��-����}:U���h9#4Bw~�<�ժ��G��	�z Զ�Ɍ1!�*���2����5��DF������#�~0Vmu�:��Q������V���,_�MZ�gW��~�൨��׽Ddup�P)VS���R���T�72�v������sz��P���	k��>⠮z�#�F2���qO��q3��D���ѐp���[wP����/y���*kS��L�R��aY��bFt�m\��!�nWϹ�֦�ϖ�ĕ:H��E���c�9u*�����(����ڜ�k��w�{N�!��=�����uw�����ɵ�	�ؖ�G֪�46x7b�*���JФ���)N�ZNF�{:��� V��O�/ܴr�Zم8
,��׿ƑH�r	9o�'[��͚�[{�W��V�O�蝲G�75�/��V���{���[�KDje��j��V���fX[~T��Gg���"Yyb�R|�d?�_|���:j��`V#1�zVdj��]~��a����yq"s;��	X4%��j����e�.8��||����m�Y+���Be$E��5-�y%�Cׯ��`�X��p��s��:���O���랩��\_{��gR�5�ܒ���>؈u�*����D�sR_�ц)s��	@�g�F7��v�aj�Fז�;2V렣��������?{�gF�4g�����`���+I��%�I*��&���ҸO_���u�8�ޗ��q��Q�B�ұ��/N)! $��K'
foCn;jV���?~������|.��g/)зO=�fX����Z-���yl�"k�7|�������[os�M�Y���	~��HЊ��㲢xJ>��
�hP�A�sZ#�[h�/f�1&�������}��l��O�+L���D:�ݙ0aw����]}��t�]���J0 ��������㌬j=� �d��_�U�l>#W��ʺ��U�O�Ox0"!gy��V�T���܁y+��k�5�{¦��*�9�����]dDF`���j�l�>m���k�qq��6G��,N�Gge����f��v�{kQO~r"თ��ױ�0�(#Y�aY���,�g�M����}��h�ݨ#��wM�}����L)3'�D��(0d����'��yK�p*jLL}�	ӝ����V�&}�U���zU}`�K	
v���-��XS�Ky�!�JWLqv�&z��j�{�����n�8��D[�J�{s,VZ'�8t����:���.����V�Y!�zz���J_޴WX`�@*R�~T�=��Ш,���s�-ڄ\��Q�9E���X� N���
t��^��/IH�pH/"o��(��ۨ��Ү�%8�H�X+h�SQ��ts����0;t�K �ܯ�,�m��a��Ĳf�l^�3�="��`�6�sk�l�� ��-bh���x��d@6F��6=�]�;n$7=�$?}�� �̢ډblf�O��6� �zl'���a�����f�U}���k���dO�1�DrRV6�݀��jY���* k��ڄ���S�\�Ʊ4)'o��󈪫��`���O�e9@��-�3�=�d�6�N�k[������bT�b�}p�}_NU��&+�*��C��( ЁxA���o`CB�,K���}%��*�L���*�K���2B؉b�p�����75���'a��)x2����2'\� �4h8�bB�Do`�	�҆>-^���da���\+��Л2�~���sZ��xRZm~TJufpg�r��Z�L�M,
H�57��Ḁ/>��͞R��L��*��|�>/��t\b�)�>�풷���{�+�K=�[��w�:����|��,�r])߅�Y�IF���`�V����ߎo�~�~�깳�6�mkr��1�j��N/���,[�U�_80��SL3�m/��X|��t��a����W�b�o�t�����
M,�l��$�)I�+c[�%k��`�.x��〉��[��YWǇ� ?*<����%
�!x��K��l�~G�ȏ�Jֹ\+�x�@f9;O��fm@aj&�N����D.�ހ��dM�Z��HG%��3-��0y0z:$��DV�� �"�h��i+%�L���{E�ʣ?�0�]���|��c��u�bB�7#�ϊ�Q2�f$�9���k���{�m:�*���Q֌5�c�ɠtv��1A_���U~�����
�`5�w�w����9XC�a}��>.ܒz�'����2ihC�q�P�����+�;��� <���ǬX��eߝs�}�;�u�Ȼ�	P!6Y��>��@['\`�&�!�6�|o��p?N�E�䁧������#ü �լ�"�=��a�Ȣ�M.3�
�%��8���k�3��2##Пψ�d1L�뎑`F�p6f`B���(����7����܎��^�NM߱s�B���1�������N�z�6nR>K�1L��1,�m��5t�a�M��1H�P j0���h�=4?X_c<.��U�3��#y�.�g�[�xU[}��]&��ߩ�P�p�b����f�U�On�|� ���jv'\�;!��%��Y�S�� 0�1�� ���szE�.9�$
Y0�$�b���O�!DMZ����X�H{�D���k�;<?������{��r�G��1Ih�Bs5G3&յ�K�%�2=�W�����c
d���h�����G���ҷ�uCu�r~ 4�̴����#��F`�4��g�f�G]r�e��=������"��mM"���`���'<=2��o����.��Qd���G�����C��H�^��*R�ܹ��^[���YHi����(�0���ۨk��[u�Er�ȋ�6|j�uQ���d.���*�/ .���M,�X�M�
���M��2{e��.�j3JDb�sp�n�?��=B���KZ�$?��h��EԻ ��9�q���?>���\`+r=��Q�$<#��k=N�e��/<�8�E�u;7m��c����C�/<�8/Ұ�r:Y�X�s)¦�b���Bg��T�l��:������:���mI�S��)�:���Ȏ�`t�ϴ�˂��DJ���<�L���L�,��+i� 5R��yҥ�d@zPR��j|1����_�N�z�`-�W�E�C=$��չr�J����6��AT��mM1A�6�P��	|���Z��J�>b����Z`�x1�.��8�^e:�����Rh:u���n4�P�2���鳔sq�����9�k��p�.[���Ĝj���t�h_�S��Mz��}qUH�G;�o�Åp��%퇄�绳���v��D�����:��1���6�� ���[�y�y��/��hv������S<:/qH�˥�����1��ۀ�: U�vj�|,�Bp�?ئ�?�B~�}%cIWL�]h���]9.�;t�#[͟Y�G�j[H�ք�T�$?�pn�y���3� ��I# =F$bu:\!a�J.�>��Ldk~��i3S�ߵ��cy�l�+N�P�$ʝQpy�EK;7IA���`�[��ٛ���Z�$"��q���v�R���۠�u�#���O��_���Z�n�c�~Y�_����Mt;�J�*�N����?�w��N���Q]g,&O��pt����h3���,�k��2<�3x �(⊁0q���;��z'��� �Pt�a�X�F��G݁�����9a�pbZ��/Jtv�F����b�H��(Mˬ��B.���.�H(�d�y]�.ɾ.��)j��'��/���\���C�4� %�c�Rԙ�8��'0ܷ�h��B>NK��i�g����B۵�:��ށ�^�]��CU]t��M�(G,e����=����A:� �񾊒����f�]匔N߳$'ȴ~��4:b_(��R�_Vë)���!>��� R [�Γ�W��#�9l�6����bH�%�r��L`�="���t4�,vA`~ ��|��:�L@e�yH�fM�oԛ�m�U��Q�,�q��'g=�7��/(gϻ��(����V>y.��	5hU�����C�E���:^����F?o�{tB���3��/е;�zK:�k��o�_qa��gl)O��#"���g�Xm k��D� �Z��߉�o;~T��w���~D�ɢ}� �E�:� /C;��S�2���9��Ys��M��U�g��D�yE�a>A;�}Bw�&�:]ޖ�e�2F��ܵMF����9���ft�jr\��?��	��I��lۈ�𢡊�r�Ħq�5�jC��%���/�_�c����0��9M���b\.�+��(���N�C��L�36��j�t���]��3%`Z��s�L�B�7蕙��	����q�uh<��L(�o���[�hd�9#�R��M<�U�.$Ӑ�k�j�g$�x��c���K�x�)XX���c��X�Q�������� 5}���]����c��L�d}�R@�� @�a�Cf��C��'�	���t���.���d�˸s�TF�v'@>�Dlez*�}�1�?s��>I�TJ��	�M��D��`6PD���'[�m܃S���a�1�����D����0�F���Y}�s�\\�ǖ"�x����J���ke��XKK�vˢ9�k�+�s���������.#�����~�ĀՖ���@Q�<�ߦ0����L�~����A%U�J㄀�e��"�s��}���.�%�e��GO��Wh���ƃp��ݮ]�>�%T�6�j=���U"��>�� �h	ݢ����"e4�xM����8e�;S\Nm����:
	�_��d�'� ���䛒<�e��|�ǎ"N�O㑰}�����S&˂,IW��T�-8�7����݈�Da��&U�^AO�<�� �U�=%�jĬԢ	l���_�i��nk�����!'�{<��+�l�H�#�Jj�L-��-։�>������3���i�=�Y�Gof�2w�؁�`ךAɩ#A�p*I�F,I�;m�nD���P�&���b��V
��3�,0hpS�\q|l�Q�$:^�*׉|�q��Q[p����D4����+4<���c�Z[���#8���\5k�-�2��%���Je���#x�B�6VrdC��V=�OB��3�q�f�#�S��d(�*������O��OB���bY;������-�%�Q�)m��?=d��UBz��0�c��6,퉗�f�r�� ��g�ˣSԨ��F�V�ug<aV�a�!�@9�Z�l�z+U
I	:#r���I?�B�	����0������tI����k��jN=p�W�s��/`��m�i{>�-����u�e��������x�c3��:l��%�Iݰ�=�[����^f���3+eh'�)�cjo�𩤉�p�Rĸ0����
�x�v0)��"�t\�?&	��o!���ϰl�+���L�	�|ЪR%8����&s�Z]հ�h�?{rB�hu��,�kg�]�9YQgss�$�� �q�̙fz�y��n~��L�ڭc���$�^)h7��tKj���_�uR�3 ��5��̝GW�`��@���7������u�e�	HZ�"�ur@R���k���Yv�S�0���P�y,���&h��/�s���	p��[�,%�#�ޯ����ɥ^Y!h'Y�R�i���K�`\������k�pV̲��L�D��n�ӋR 
�L�WX!�d��ٗx&W�-.F��f�WM�y�����XH0��%5y�vOm�y݋�b�i1���#�%(����^C��]��
o0���	�u���-&�>#���hx	t�h����[�;�`��*��pb�r4�\7y�ۉ���ˌ��g�D�H/M���&�r+:��D���]]�Ԝ����H���'�6#��7>Gi�\�FkZ�*H�ssy\����2�T����=W���w��Ӂښ�h�"���H��P�3��n��O���P�Fl�1{:���3�j�R$�����\���f�7���閃J79F�J�5@�ʝ�}2�tq<m�h�� N@���K~����`b9�J5�0"���ߕ,�_�Nײ7�_ܞ�O��Q�X�ϛu�|������Ͷ��{T�;����``�4��D�{�ND_�UvN����D���F;A�,�U���.����zn!~X>�V�Z� �
���HwR���_�KB��Դ��N�Y�oƂl�Y�.����W�?�֠��7��i�� �&������#��P�ȯ����6{QuY�s6N�����#���A�E� �����%��2u�!�l
��Pw^���pq�,��V�����Up���z�j[��u�|�A��g��I޳̢}���6�߳�q"�Z�E���}�([O�<m����ꢚ?K�K�U��~������@
�t�wbg�I� F�];��9��qiZAh�+�.L��� 7�j�M?8Y�d���&ٔ����2Q��K�Q�<�Ν[���Wv1��M�
��s����o�.��K��X�D���x�}�O��:?]��5����u:������Ƶ�
å�l�h1��OY����[v	x=YZWJ�CU��}�b��J���cQ�ױ:�9&�.��,��#�B�N�鏄���E� mS>�MD�yK�w�9�*r�Hͳv�t�|���`V\�v����]@׎��L7،s�{�\�;���꼉-'^_ �.u�!� ���B�~S��F�+�l�Nt�Fz�š_}Sc�p�&���@�(Sѵ�1
�u�3����@c���p*[2z�Hc�1:�^f6�7b�(8hV0������TM``�3���a��V�>z���ܸJ�'���$�4�89i��D�u��B��Jy\�R��x�����;��wZKa!ǜpF)��MމWu�L�8��M2�Ov"�L'����)*�hCק��v�w��E|XX��$]6�Tߘ�X!G�|�F��'1�:3�@�Kˑ�}?�]���dby��BsTX%���ɿ&͛,�sb�]b��AEL��ع:����i�0T���pmdk��4#�uf)���7<����\�<��};����q_�<x��\H��r��Y��haK�3R&J
���JO�^�7|���v�l���Sd�	M��љ`O�����d�?q��N<6pK2�@��]`�Yp�拻�r~�P���L)BQQv�ޑTS��T*�E������DM�q{��R������vrA_=��f�K4�:i+a��W��-<_�ԑ�=�--i-���6;����1D[�4�Bp��P�e�l)s7�S"n/����6v�6w�����QY}��1��ńo$���j�>��_��L,ݏ{��Δ#�<�P�p��WnK���}D����[/�B���Ŝy�k{�����^Z���L
��FH�F�W���	��p������FL	��o�~��5o�ԽA�hΣ��g���h�������=� �3vD�1Cd���Fp��;zC f����lR<H3�������h�RyQ�n������ɭ�~*����?�v��:���<kI)����c���I�{�b��v(�����MY�C���nS'�:�ͬ���� ����� 
p��f{�>��p� -=�o,OՇ�bĄ�e��=q�(��W�C���A����ҵ�0��@���ɡ"QCi�0�wLyY��A�5H���G��anX�d��i���t1v�o�:��p�cǋ�IV<�e�X�3��"�Z)Џ�*��i�=X��}�Qfh�Y��%gC ��l ��a?Z���)��U�V�,�.����o9�\��$5R*X#�7S�0�ᜊ0�Tk��7��s|�5N�6��לD]|Sk��������ܰ��I���#�:����՚}�zᩦ-���Oy�V�u'bDӍ!���`���CZZVzW�O��R?@��3ǐL�C��f ��B�_1*�%�5���g�����tVCh���!��Vr��CAŴs���{���ێZ+�x��_PJ��ӵP��o�����"��4�����_�U5�	�������.������n(��C�AkO�
U}N4�^�\��1l7����W�_yB��U���l/�y�)�&я'T���)T؞� �2����k˽���ZB��]	�o(2w��
E�0�X�KZ�ԃPU��6Leb���ڻ��x��4��'VX�t6�4�Io�����;�)K��0���ہ���q,ˣ�����|x��8OP���c�t����<ؗ5�h#�\�
�?&�ƞ�1Q�d\h@�@G�3wg8�Ң��n4�
��Ɉ)"�0?*�.rfC�Z���J`)�8��se/�m�4z�ﳉ<���[\ŝ�r<���~f��*z�pV ]XG+?�X�08s�jhm�#����4�v���B˃*e�-.Lk���3�T:��*D+n���)}v�IC��mM�1�l���^M�AAt((����sxQ/[���D������U�Qƭ"��B�I��Q�w�hU�Ld��u�q��0��CwD�!v��=
6�-�>f}��-�\���}��>�m�k���q�m���1�H���v����#�+&-2�� ��L%�]w��t⿠yߌ���$��پ�^�8����n'��v�4�jb�`���kɾ�nҌz��� ����L���{f蘰�����G�Rߑ���5��gL����h[~#���<xY�s�t�0���M7�{�^�ǰ��"�ȸ��!��[G\�"��)��P}�E�h7VD5mFY�i��nٶ��]xql�>L@Ə9z��پ
�80i0R� ���zu�
[[Мל�X_�"�R+��@���l�]_���]c�Ӽ^�p�2b %��zۍ�=�3���F���Ġ@�0n����f���7��i�K��рڗMc�%6[阀,���t�C�0��-ݹ+��dkI���{��Q�P��&3jɱ~��+Iw��$u �[���<g�����[���C+�R�]��Aٓ�.���q�#5[�?z-��^�|1_��E���F�7�1s�J9P�i@��b�Ȣ��
F%a5����`���q�*���=�g��"HsC~Y���%�k*�ͱ���<�}���K��JE��D����תuO�[6�o�ĝ`:���$�X��H�E,۲��d���-٤�MKѶ��J�f�Mp��/��7�q���G,&k�������9<��*&*�1�d 9S�߰��Rg2����#_|i~�e^��C��^�뾁O���1H`�A��x ���3uګKI��݊zN��{�E(�z����X.�����-#Tsf���]K���.[����:X�5	b���1�C*r�`V6�u�\�Ք��^(ԧ~���

:�w^�:��S� cp�.��2j��GQAƆ�rV��v�ҝV��ђ �gBg��Ȑ�uQ��⁙=���C}����a���u�ü|����6�%��[�=2���rݫ5��O�����S�jQ#qw������I��	��g�QWJ�SeA��1pxhoa���o@��� >K���5u�;�8��"��!�ƅ`�JKY��(�<��� c([����4�� ��|��}w��[Q��tbj�
ǖ|�[޺>7}�"�j�H�@a�_��Ѕ�D��X^r�7�%M�k�����.�?���J��X�CG����s���4�`���e�qIe���/'��ԁ�����n 2�p.��B#p��=p4i�V��fv��I�"`�/?!,�?׆щ�t�,v�
�Kٲ�̐N't?���ߦ�ӏ���L3��E�Y��K�v�������7�U�~��r5�gT��
Ӏ@����d��`ԦIv��b1� is��p�IRM�z\�6��y&�Cv��R�{ɹa�d�$�Em7Խ�uj�B<,���x�޼���*�q|a�{��Sb�@h�՟��4+��(Ŕ��H�Q�e���ԁy̶vn��\�) ���L�h',)��aȓבI�{����޼kw�N!HE��E�#�X�l�y�Z���n�����E��b�k�݁N�������7֤�PU�0��g�3?=s8��6���|rx���RTh�^])��y%٩{T����¶3e���Ⱦ�:�w
�Vk�Czk/6ۍH������w�G�Uv���d��S����OJ+,��t�֟��mم����h�2K��b��=��l�t�xK���8-|[*��f L��j��7����I�-m ��@�aј�Q{����jş���s6Q�R3=��ΟKC�7��%��h����՜0��@�� W��牤���=X�\ju�oO�{�=�gޫ��h��*"�64b�o�q����Ƥ�w�ʋ3���X�w�"_V{7�&�/c[���G�@�G�bCH-ZG��^@���F�"�؞4�~:�]�T�@����̑e��������.X��w��t�V������j*N�1��8>���#�P���CvU�;p��4����T5[���O[��ہIteR:+.�>��5�%�����	/?,1+��^~Ҡ�r�,U��{�b,���(1�5��dqUl>�xm�m$I
-0!) ��q%r�\��I��Ě�f��[ͮ�r>��6���]%=������j�(��L����bj�d�w��:n4R�o�?���~r����B�!=D�7��"p�
dmi�{��N&V��D���>��!�{��Uk�x_Ok�_�c��������F <�#l!l��A
�t��8K��u���卽Q���5WC��¾N��]�[����(��nSk�'�c
�Qje��(��j�*�ݿ����~o�amW]���RF7�|��cN�d��M��vS],L��3<0��7�� #?t�Ρ���B� A_V���0��[�wxg��B^����LpBM�3��$�乌h��"�ڐ]Hd��Zr[���Y���g)N�e?����\˵�n����\���7U�7v;i8Y��H2�áe�#6���.���pT3����6��	|�&N��m^���q��ƣ����P����sb��,���ώ"�[8jU﴿F�i���kF>o�x��X�3�\ߛ&�/\ �UO!½�O���s�3�R�ERᅬ)��C\e�s1�<�J�e�c�0Tx$�ݧ���+���Z�7��
F�� ����-j�	�h��t�I�.MS�^�����(69Y�%��P��oz}�Fi��	f (��[�@L݋���4@QZ��� �߰/�g�
�K �c׼�e��R�j� ��r�-�՝��Y��Iyd"^ҡ7O�Dd?	���,��vk�΢͉��X�aLCRd�����8<�S��,��7���w�ƽ}C@tc�?�0���5�y����@ �6��ū.�X��������0׊D��oDv{�����y�[��?���_8"�/���R�o�?,U[���?|���#E�M�c�co�;�mR��N����U�Y0e&��<Jv��iI. f����p9ԃ�=���<~�$3�:��Y[�)zT{&���v��o؟��Cݙ�$�����[k80F�Xl�*�����Wt�~r��근�Qzk��\jN<j�!{���I�j���;�C��!�a�\^C�_��0�x�D�(ӗ�zYu1 ���(�(u�F�'DH��_܋m����>�'A+��Ɠ�+V+�a+��^vo��J�H+.�����k\�ֱՉf2w�yNz*CZ���7���er�VOrٯ�wq�J;��f�*y�����0���G�������r!�	n�U3�ra�}�^� �{ۖaܑ"o@r���/�#D`��ʣ?U�)^��$hA��PQDw��n�*�;c��i���(ʌE��j^V�jV6��9J#�1���!X3��A�����F��=�
sD!�^��J9�HvA�9���};�f�(@�"�oQ6�4����E8����P�_�~h)�a�K4s��նi�e��58��k�s,e��β�E�I�0s��y&�4���]���n�w�F/���q]W0}�0,�3E���5�]2�~vp`k�����g&v%�����p�cP	+�&w$�h
E�7Ԁ�$1}�V�&�qN¹I�]]�p����-��em>�Fz��^�P�-/\,���+�M$]<|���!F���5��Ґ��4*�P���Nv��1���B�����/������	c��oZd��<����KX��0Xsg=����7�;��B�|�gdmK�8�:O��N8J�>���t�����W�@�3�!)zDE$ޱ�V� 5��cH��m��l�fm�w,�Q�y+b�1 U���R���p��>6����,F��2�3N��Y�Ēu�n#b�!��������������s[i.�*�ϛ�:_Ϝ{��%
�{G�?_�!�]%��;��b`�:����6C=�	�p"T�<K�#\�% ���� ſWx��mi�M	{*�߽�-��#� ���R��T�d+�8�5��k�R:K#�;��ͱDƩ��R�?���9�ƭ�&M�A�@q$5��< �'bEL4�Y������9�tt��Q�Q��U>1KGC<��b�)�Jǎ�:�X���ݧpT�:.���0��w5���`7�'V-+����ّ~	}q��Bp�)V�����-,�Z�\�u�T)׃<�,�n)��r}��i���*
��d]]5Ý�Z�,[���v>Z:e5X�֩+�R}���!��",��k)cmM@��ѵ��JG���gdޔ�����{u"�v
��bG)&f�&�䴔6��� �x����q��/`G.�h5o�l�v$u �l���I�dc��]p8����\�{��~z#o�����H�}�@����[�ߪ]�΀�����`��,i�׹(��׸�e�#R���TS�`E�E݂�e����ۦi��DbF��PtY������Q�	N$V�������dm�0j�(3������0`zg��P�d$=��	Ï�y�6WfiT隱¥.+�y+9��&����L+��as~8oR�W�<����6|�;/*����%�4��'��G�4;U��/P\�`�TL���]�L��;��
��b ��
�zx�������;boKc��:Wg�C@:�:"���;�^0�lJ=ĜgP�4f�ؼ�.��D��]@B
-CA|�\�_Ԕ"��z�r�`Ů�k,����cc�J��V_E(_���c佮���[��FZ�q
���I��	���-��a�˘>w���'�`��x=�i@��N�p��@w�?G��dX`�*�kv��]c@履����R�{J@��� 4�fύ���O�o�b3gp�\=�IX���p-R������?�I<X�,#4] ��3<�z�S�}���<�٥(9^t��_��4�f�y��DSx˯
k%3�����쉯�ۋ$2��䁭���b�07=ef,������7wD�����Y:�D0�U�����oN�G��{��qB1� �q�['o�����|�0�V��=�H��a���O�=��g�3�*/av���U.!��&�SA�~���7L=�\�7���,�)�l�O[��o�de���,��e0rW���9�=5[p��L�G����>��������2�����Rp|��e�n"�
�����+��qM�ס_�DK��&�
滞�RԪ.��g��%Cl��79��V3ц+�ͥ4��������l�D�_�-�[���f|@�rX$�O^Dc�G��KV �u���"���(H�Z<@O9��Wz�?T�.Ϟ������Ow���jc+pI�Q���F�}i��崏gl�h�FY�F����^1}����x��7��8�ş���p,�c�"Lt���6�;	��L�&76y��ѹyy�ĸ.���V�6'�	�"�U�(����N~M��͒�b�I�h%Pã���	�`�i��N��>E
g��������������J�����0�Ѥ��bX���4#P�t��ఌI�C�S|ͮ���r�ꢯ�LR���ţe�wʖ�^�3_�?B9��h�Q�}����D�
Έ-<$����P�~j���Cݰ�rM��1�W� ���ӣ:��LwPI��ǒ�@My�{�i!=�e�񻒸O~��7��������d��.��3��U��m��ZQ���w��B��u�*Tū�����'C��Q��nS����H�_ꏶI�����!�A�1���o+�g��i[5��!�J��-ףN��NNT�!R���֜���!���ג����V@a����~��)�2���1�嘴��LW�R�G�e�V�O�D�V�m�b0gf�z�J`$�I��$��?2���FH��yJ���)�'r��%(�lΙ�ȇe�Bk�J�CK�Czgc�ռ��i����1������U]NN`	G��^8��6�V�'4D�	o��1���S#�zU�A��ϊ��7�*WO��C�0XVM(mђlR��Vlt��/�p��Yc=��eA�WZ�J�rɚJ�����3����io��t/AD���B^��� ��Ɣ��L2or(�4����5J�{[�əyq�(N �%�^ ��_��R>�aʿ�m`E��(E@D;�Ɲ��o���D��v��q�( ���i!�7�͋�1=���m��:L�0���fm#��BKg�v�$�%-6:����MH���+��aْrA$DPN,��!Kt��%�ڔ�v�D+0��#�
��ǲ�P���!Fq��Yd(���� h[�{�~Jr�X�
�g�������$.r��}w=o��0LRW�_@Mu�r�����E��'�eϫ���AV�|j��I�sz"W��7,l(���a{�~���%u�����;g�P&C�\�eV�j�����97�����$�< �[̫���^�v����M�"�A�I���*$��|4�}�؊)�?a/(o]�v�s��h�{(�`�|.IF�eE�1=!I���sxC'����q�����S�Ѐm����,~T����/�'l��U�j��Nd�D��INGi-ά����-�0��H�>��&�ib��ˡ�@%��j���\	@�޴�����V`��Q��s6���9� 9R�k'sKi�l��+����PQ���������w�_�' �ɏ%C ��� �[���[),�KSMm�n�-B?��Vb	���|�-=Z �L1�^�����I�5�eLo�_�Fg���P
O&���@��K*l�{��K�&G�e
k-Aʼ]9\V����/,\�7�׌���M͇���&��H�pHX�H5W�u��!��PMNwR	MՕ&��!q4{!�8�S���h^�l�<T��Ԫ��Taѵ�C6H"�(o��f}7�� �$�X��?�/ކc������P���7��jB���N����e.2�[
uA/k�m�>W��"��3����so $k�����#��X}�8���~�>[f���M�0��շ,�ٶ�D�j*�q�a��k�a8��"��~���Ps�������5㧙�2?�gO����������W��e�#%W�W9GF�]C�?��Φ0�Ī%��|��xk�sޱ�2t����ǨGZ�K�>��a�x��cG��N�;����z�M���)Y����t}�W9��5{qU8�ԅlLQ�7����>Z{�}t��mlL�zLH ��
�"�*�S�b3*~/JK�Z�!�7�U+���FI{�Y��n[i�\��ѝY5��t��܄�0D`���6�L:a���M/�����n�Z��^�S�!����na�<�BQI7�y�)QqD�)��~��ɽVh�U�u ev���.w��K��UL<�t�6c���nf-+Z�n\ջ 3����=�5�_ODK_��������]iE�zo~ÔN{y�k�������X8X���U�KWv��zC����w<Y���)j`���s��sN��i�����r��ߧ.���q���Ƶ0���Q�%j.dV1�<~b�r�%���p�$~-�x�j@;����s�s<
d#1�蜙�Ce��oU�P� R��$���+����nm1�d�A����p�*Ν��n���5�өs�r���������)n��Эs�$�^����s`���t��e�ʖ[����>v�k�M< X�zeMOZ��R�.)y-�W1P����e΃��T�]O�T�|{9�.C7�kMt$�/P��:'�8����7a���?G�Z��c�0�H�URJ�LK��;��/	��*�XcK�]�B�C��TH�|@>��}ou���b��R55����������6W��P�D�a�	{�g�>4`r��wq<����ԋn¢�ٝc�H�A�0�Æ�wl��Ru<q�me=/�N�b���`���a�)!�^�mF��N���c�dY�R���G���,�Z��М6^� �@#��G,�{�����B!�f��m��c�I
�`Π��#��N׍�N��B�H,�&�&:+�x�T��K�G��o�o?N���������Qk{��`�Юi�q��q��B����dJLQ?4��R�]��VY����]	dY���%&�D���6����R�N]�����Lf|���o̯]I���E" 	(e���F,f�����j-r¢��A�s�
~<����+�����3����8u{%�Lx�,����0\�:1�J�qwg��7ADA��Q�#�[�K����a�$>w�$�L��`=���]`�IR ��I�C�����y�ך;�s�Yb;z�aW[��
��?�ќ���b��W���m�-Q�R�i0��Q�j��]f-9ES���0���Y���R^6údy�Q�ta\jy��M�(����%�:6y�Z�,���n�t}$I�6-�����5�Qyp�B��j5!�R;QBN������Q��2r&o��yt�M��y��T�6�3K�������Ƅ|Be4o#�K�f@�Շ�	�J���|D����������E�m
�T�Ly&���p=v�ٴ���uț��,O�c�q�m.',L�Yr�P;��7�ջ�iכB셣��F��Zl�Y2�5�B��nh	�����^��_Ϩz�H��I^�P���Sd�K�)��%	������˂3�-�6m�l8T�S3/�=���׀xQ}�' �g��c�˳���g�a�5Qz#jYস���pH���aD���@=2,=�+(g�?8Y�* O���Z`�p�:��^�i/ num�ϨH{�'����lA�Y�:�).J;�!��}�	4HE�1�.��dVǩ4�I�����˫��  ���y��(.tW�R�Y����͋�'(�QUu{�>#ÍlaM�C;�oG�<`�����w��`6<�2J�y���6ʳ��=5���g��V�渼f��;�1Ƃ[�-�\��э]�m.��Jw �g�%��蒡�+���
��r����L#v�Ff�Ky��A��ʿ*4����١�dt�e�ć��C�.e��10	����v����%	qB��=��+bP%72d&m����,�c��5�.�Hz�#:[�#��lI���H��Pw�mr{7ڥ)US�%Pq�x��N?;�+a�A'��mG����h��T�KO&$�2��&&��}�?�,7��f���L���0o�sJ?}n�`f�Ø�0�"U���&7��s.s�haMק�]SZ��s�p�]k����3)��r��{Pr�'��,�7\��dʝ8�y^*�	��e=ջ���ͥ�LE�2����Ƚg�mT9q�m���Ϋ&12�����a1Ģ}<���۩(��|u��ÍYVP'H����"�!��3o� �Ԛ������Pg�!��!���̊!�V�����(�t��W:�Dhg7Y��Ί�Z���7��m�sT�n>�'����68��z� [z�r��@�06�]�C�(��s�3��.�;"��c�Ͷl�jFo�F1#�49غ��%V��O�P��� �t�j�%��m��#l���t�H�/7���v�u�� ���+��i�O1o�@/�
�:��np� F��\Ñ&�8�?��*x��UQI����j[���ө��_.����/�M@�)tu���R.m�U�I�u��AC�}�d�Z���Y��N;6
g�u0� �e(�.��tA&P��;b�q��u3�B$��u�i��<��C��+.Vuv�H�w�!��vחF}!A���ۨ{&�,h��Vv���'��z5���2.��%�na�I�'��K�P���H&����Z�EiV��QL�P���?��C �^���a&ͽA��ż&�������������p���a�ț���'�T������6�G<L�k.�TO�2�R[���*�^S�N�����!�l����r��T���]NӰQ; ���	(%W�Y����E��q}�l������+cEx4VE���hE��l����_5]^Gɝ��e�����SS��R�=�*�+��ӎ��,<�L8$P'�<��	A�-n	@%R�`1�e�U:!��ȗ��0��;]Ho����mDY�Q4'��V61�7:}�a^:��-e8mB��"���mK��.P�s�{: T I���u����;�&�Y���R �$Tp�A#6&	�b�?�Q�8j��"&0Ҁ���B �W��c�	W��ׄ!�<�����nU[��z�2j, @��t@@���M*�!��AҊ��vy�N�&�$�uQ�e�F��}�Ȩ��C\K�|��r�)~�_�U���(�3�����:F��p#��L<d�^}҂�z���aI*��x�q񏼷7��@CI��q�c����;@u
�j�Y.+���_8
�H=���ǊR{/���Qr��/�/V<���:`iB.��!������%
��I�gE$%m2��+r�u�;�HFF�Xf+f[��K`�hAȶ�B�и$F�,t��ҩ���vj6�p6��BY�B���Yh�U�F�� �	����hl��k��	ȗ����@恵7:b5.�1���P�z:ܭ�ޞ��S�YY�Ĥ)>$��B[��ו��e�Lk�_`���v�矁����	�u�|��e��_�f��i@Dw�(��?V�N�*s=�`�9�]��<[���:paڑa����CD�~s��ouE�U���m�UFH'r�Y��KK�*7�l�{CA���!�_i��,��9�+�5`UvK"�2c��7,�)���:�}�4�5���C8�~�<D�+6v�ڲ¢hMR���-@�̦R&;�s�V࿆P�R=�vV�3r��؛R~�d�~�3u.�)7��/W,��|�#�FY�Lp���^�����0�]�E�{�0��+�ت��>s���>e�vBW��y��'şrG��r�6���k��c"�ˬ���j�wl:Յi`�����+N�a��}6M�X�g��{������s܂
����q����$�]�3|R&G�_�|ZV�~�LD�7N�%�1���ky*��d;z�
;���.	�o:��zq�@)a�7�$���I�194�2��i8�GI�m &! �ӣ���j�����)��g~\51zr]���Xަ���?mD�n^(Ct��e,�uQ�+��Ř�9���\l&���ؚ^�Dy�\�� ���˾�hr-�vT�i�m؅��DG �Di�������;`��n�3��8���0+.��Ҩ#A!�������]�ր �(�K����ҨP1�\�#��e٭�<!0�U�ذM�g���-�9����2f�f�9A��,����._��y��P������H������ǯ#ơ�᫔��
����~9B7�
���L�����!_@6`]V��eZ�֤�&��E�b����An�|d0x� A��Ue�vD6����h9��vWU�[�ɢ�)R�ښ65�v�[� ���U�wm��a{�Ei��l/g�Qažɶ
g��ׁ�ь`�wT����0��P>k�c���t��16��-.;�͐p ˡ�#3��مǉ��
�#~�f�>��mV<��(I�ʇ����?=X��?NK�2��#Hi�L	۔R��!A�l��Q��0vKʣo%�����4�.2�î��ǷzD��Z���sgk�dz��ң�Y��z��Tt�٣�rt1�o��� �ϒ$$,c�q�r�"���2��&m���X,��ԩJ��v:Y�=9��D¿D�FP&�i��S��(�O�~�R_�P�P顂m?.26*��ˤdO�'�191c��??񛄓�9Z�z˞|Ž�84�Z����{0��e��[���d"Q��/G�,�{�X������5�yf7(�E��}f �#�k�ȷ��ev��'�J70`�|/�j�1��5f��i\�ot������Ƹ��ݗH"�z��fl2|Ѷ/�^�l0�%̔k݊���6M"�b91P]}��HXJ1ȡ��`�h��݄Cm���M�Ͽ*��D�uD��i��0����݆lv��u�����@fn�z�qϐ�����9����S8����mw��5~��@j�a��,b'Jμ�K����F�d(��h�:�oD`h�\V�Ǜ�L�h]�<+� �g�>;��A�7�\A1%S����|>�H(Av�H�_aj�z��5�֟F��qw�ffqi#ߝ�Ҽ�TzJ#-�F�\�P�c�"&r���%N%�!�r����&�5������O;4�s�Mj�i"G8�m$U��tIH{��G��nnK~]�t�q�"RԺ��e�m���K���؂iE8%�(f3����R���^�e���8�0��ō텆4������r�nVf*Q(�e�QP`�����B���^�@m���98 ���3�A���Q
�`�>�(���9�����ң������>������Wd����f�5�w�F�Ȍ��/$4*cV��K�]>Q��W��V�
ʏ}%=�߾Z�!"az��v�^	���]��9x���������<e�f�k���r��E�t<���/ KC�������S)8���	-��J��-���G�BRHo����t��EʺPe���[N>�[����[ͺ��D\��i4�;p�R��]5���ꉧ1�Dq�1i��
��[�+�����%k��>%�T0N��f����y�cs�N�F�;�@
l`���C��8�A�E�	��J�������^�)-]m	��"9mEύ�^E�3#e���.�������~�t�8�.���
��*�C�!�_��M�?�PS�Qd�t�j���ѱQ��'|E��Y���c��Ti�F&����F��W#��0��܇�S<?����m+Siz'?n����h�0���=Q�lx%��O��@���n��6v�a�+�ro.k�Q<�͂;�^|�����E���"&f�pnW�(�.� �r���dM�<-����&��=���i������3��+����u*�6|[���p�h0;���1�YH%������H�e ;�#x�'Pv
.r��1H���%�� �a�����r���������Ô�U���\�r��*>#�&,o6�ўIԜ� N:�Q�s镘� ��{��f�"���ޑ��&J�X�)&q�[·"�� A���3������V��cǍ���p�-����V�S'gdiIR���Zw��WW�$G�	o��X��d�-�������i���{�X)�H48�X(;$�o����&��8U-i���.	u�w+rEO�a�(�<G�A}�J���0���Ƚ��I��Z�>Z脀�N�1���]�%�`��x�;��`��.r��:�櫏ƾY6i���9:`����+3P\���n:k�������1����T�`g\Qa]�B9��M����\�3�.4&JF8�S����~�+=���&�T����:�� ���oU���L���#]����?xGy;���2*�y�VI&gS��s��ԛj\�2���l��IZN��r^�^�C���h?�~��z�o��`�!c)1�/D����lb��(T�FN9�֋���!K�h{u� gjk�M�ʡT;���Ή>�q֓ �d�����8��K8�V�3h��𼄕�On� } KI��)�����1\�c��lI���U���EᮾV^���NC>��BN��<m�N���ߺ�MV��"Q��ֱ�~�!��[~I�]���rAJ<xdU�|�#��X����_2+��1ڦ1ő������E���jA�!��r��Q�yG�{��S3�i�zQ]��u/ܞ�0������J1�N�[.����B��0�{X�o$���zT��Gۦ�Y�ͤ4p�5��q<����>"4�<�1���7����[Mf��㍋���ޱ
�٤��,ᓯJ{*H�,�y?5����_p��ທ��������'�dS4&�K|�q��E4	�b_��jRj������Oc����ފ~ne0�����[͐��6���m�9{� ~�W���+�.I��qq������N�
F,ݥ!;�}yب�m;���n�Ӝ^]�[���|c������@<�"���e(��)��u~���n����SMBH���1�u�1;�Ύ�S�p�@�EՄ*��IoƝ���2��jm�V2H� �������/��I�B����@!����@'���O���Y͖n��z*E��H��TFF�:�x}��Z��E�<.tp��A����]�lZ�i��9�7��􏨔���ԲG�ŮD�a~��ri!��_�<����V�/e�@���{K�u��CM�����dp�
��?��b&$�2��V��YX5�.6���uM.b��,�u�2��b�(�`��� �>�b*}F�%(�/K>�+ S������,3�<�b܀ղKC
�g2Լ�����T"*C�e'��bo���n���c蓦)*�I�����c��u��w���d-�O�,-���wNZ�����S��.�o-�G6������	$ Ebv�(�A{c�8��`���cÂ�6W�~�A�.�K�a�sR% 4tJ ,@������T������"�Ξ �*�5	���v_����t�'�e�<�L��� �P8h�����/gߦJ��߻�4m��s�}aԈ���Yl]���?�����# �I��ĂIM��iW���F�s?�.`� �ѐ�Cn���'��$�%r�!������Q�'��ZN2s�܋S�An.�-�s��y5��}t��D�{|EM�X�A��0�sH�=����]��lл��" ��y�A��O�ul�*`(h}���/��K3yc�:͟�ؿ��j��g.�c����PE��]�������Ɔ�H+PO�i'Ve�����@��������;�d����k�c=]�����w�bU	(�&Z-ע�d�9�
���m8X���EW�BB�ƔF��ג�&p�|-HnM�][��s��l�4�i�#sJ�A�H0�-��u�a�O�9vc���E�R^��K>�:S�>	�Ԣb~h���'��fx3�+)�g �r���Ë^O��������o^��X���A番��^;�]��k`)��Y (�4�:�M��ǈ��ǕY�H��-�n�p>e_&��@aҘչ��Z,CȆ�bo%��Z3�j�_��2P�ZJV)�ßj���%e�.y���+�NV5F%� Y�y'6�[�?�ք�iD�
sr�='�p[�*����Y�5�g��Z��"�ï+��`��t�|�a���L��y֍#vz�3-QD��}d\�$��
�O�� l�(�D& ��ژf~����am���3���	�����V[b�^�Y�f.$cI_�XY]��iӐ���C�b
$
O/*�m#9y�ύ~lGg���R&�qaC��V���A3�3�ﶵ�$0�ɉ�|���E���,zJ�Gd�8���Z�c�ߞ�.PvEӝ��� ��.���S��I=���O���Cm����/�xB@��M<�S�3��s{��딥�k���ۣB�Gts�qj�Zx���2vq)����TҼ@"_z6?�����&�xF��Pc����cv!�6�D�w�GQ�cN�Z-h���ʌNu�DғdމCY�TsT��HTŔ'�7`F.�����(g�.�8hbz���f<2�9胠*K���bn�ܕ�R,�cH�(���!�k��V&Jd���0\�=��1ҳ�� ]iw��%=�ki��u8�
�����-�khe�1�_����;JRP$��׷��i�q�ܷvp��$~Z���Y�E}��b�C��}�C��uo}D����侄��:.���HU!��ffɔ�q��m��|� ���"���7Lhh'yi	����cg|�x��� &�E�����f�'\@J��R(�0G,)�h(q�SF�Q�G�M�v��(l��_	fP��)Z�|������nx&�CL���#z ��N�D/�d�R������ W�\%W��+t�{��G�a���t2�A�T�4ZF�*E[D��Ѝ���5f0ޔ~�<t4
z;�����,��9�Im���&�w����(��tPtᩚ�7��QTLp��gs-�i�i�_-(�E���a�:����h��P�*�Ha��}j���]]��
{p+��E�=5���}����64Q+/�!�U
�xpP�����}_�K4N�}4��"d9��3�X����L# ���8%t�7�w ]��74&���1�Sc�
��Y���C�\�^(��ZZ�F~�8!��h����{0{�`~:�ѠH~*�-��~�
v$�!��/��mߘ�?�|��ڢ��3��ϛW��}>��L�rV�9���h����|a�'�1F[dS�K/���쫦J@�0�ҋ��M���P������ҡ�vs���(Ȕ��x]'[�j�Ѱv�D��Ʈww&��ge�����1��x�!���WbRxr�I�?.&� �@,@e��� W)_	k2�` ����Q�,`��_������T���aT�]aI��k2��N*d�"R��d��u�Cf��\��e���J��_&���]�q�Uy��rz���6X8���g�E�#�G)�{���u��[����q�nU�5���yF��'����ֿQ��ނ��۞8�w6FV�z-��(6���\ʃ��Tj3�eȝ38� �M!=g	����NJ;H�Iմ����4�#�~�_���-Me�̾� k��l�Y`$��v���d?Ϙ��:�R���n�{�G�\��j��*.�w��dz>����v���������q�Y�f�;1���
��~@9u��;��O9]o&���E�]�~�!`�ѻ��-��Gb8\Ί �3�ڡg!�:�z
@CΡ�0K;�N2R
�Un�.���QDL�`�b�l�V���Ƹ�����E�*�9�C{�vy��~4n�C� /F������
�A�=����$n������O" ��h5�O����ա���\�:9j�V�[�J�p�^;�W��-
s2�C$.��O&�i{~%ma|Д��g�5���kK��V^�P��J� 6�SŻy<,�?��V�j\�������V���	e��DBdo:�[Fh:��Z��2���H��ۊ1c��Bֹ{Q�����.z�;��vf�c�R��*��q���|�3�/�~0�Qx7<��z��>��M�������ճ��dY���}}#�6P����3DЍ�-�ҙ�ft+(���ĉ��j9��ØA4хv���lip�U��w���IH4�0��Q��/N/���,&=�O�$��k��h��cW\^��*�A7�^��k���'-�<�� c������8|Z#�k2�l4o�Rlj+x�J���$�$��֩�Z�l�P���Np��ٵQ�x+^	i8�c�z,��Ov=��eIu�P�٬1ŵBW�vd���M8��1�A��x�W�fU��5vr�2yN���?;(Jx�Ɨ�1]���M��]�����>]h"=�7��Ǫ!v`�yu1ƿ����1�y�����;wІ�����?�g�Uh��P1�+C+�%@z�C|1̑�p�Ӕ��|)R�3�m������X�as?�D\>�B����;�%�����2<#�P+�-U����y(V��p`����=�x�U)U@Bc�ƭ���L���s��P�� ������8'T�U;�>m�5�CAk?N���%��T��:�����Y�gM����a�~�s
�P�����uAOϱ�hc&1��	�0;S����XF���)!��v�ǻ:n�J�\�E���ɿ����4�X��֛%ؚ+di~Fu���i��i���g,B_��6���Z�by��uY�*O:���'�3e�m�ߋx��RA��]�P;R��BX�ҙ�1��\,1g���=�xe\�bt�a\���'4S�J�d�|�J�����њ�dф��7Ώ�C抒X��(�z��t��\Ya5��?F�xfP�$��bS����zn�������W���>���o�1�74C�_G=��V��NZ�U��ʰ�@�.�[e�:dV+x�O���,� 9�O����$Q�~Z�]���Uv�:$�����B��-�.+&���������l��u0Cq�v���Rm�ݩā�Ыܛ� :`[^jW��+���T�C�c��Ǖ�7T׳�56��$N�0����3�}bfVf�Ti܍���C pJ9�Ӧ��Z�{a��>(|������В.�8�d�5��8���FGQ���-}6~:;�pV�-�S�r�1^�,�\FG#*�v4m���t}H��Վ�^\�)��ŭ�Q�[K��i�h݊?ER��B<�֝I:�q�L�D�0��NYi��R�0	IoZ��z�)��5��L����|�w�(8]	d��mK F蚹�/4L��:���O�|��u�!��۴F���(�%p#��|�?|����)
�؟2Xa�1��`c��}=�|���k>�@&3�'��w�j��l�[�N�s�\�b�2��y^M6��C�0����yI��`��� Ͽ���
�vU���7l�z���}���Z_%�jCq�ڥ�<K=b%*�^ ��:3�4��WS�y� �1*��J�Vӵ��q�fէɶ��B��J6 -<:�_C��pyޟ<�Z��U�u�1v�ͧ�����W�"s�͹I6�M�Fl-Ƽ#��wˇ�|���mbvG+%R�$��&�X��
�T��X�ad_�j/�������V�ߵ<EХ���'P�zi@�:���Y-92A?c�7ʓ	3k*\�%��6�����>������"�]�'R�Pc�6��6����i����&�1�F�BM��7:�4+��b�Ƿ��	Z��2�Γ73`��_wwȂМ k��D)�`�q��f���%u6}Q܎��UAo�!RW*Tq=%C�ר3���?J�E7�����~��&R*,�qF�BZu6��	���ݒp�
z�KBJ�����uQ�����O��͜���j��:;=w��)y����9�N��
5��'~�oR�!�V~���YU
��z��K*�'�Tj��4��Zm��Q�*�-'���p����8��/�L��5c����ڙ��� ��'zO��U�`k�������=�=�6�y��� ��[M��˄4����H����X�:�mLs��r�P���iN��^�u\UM�&�L�x�s��٠�Z��ڻ���4!Px*��ؗsމ���Sd���	=�-Y(����C��(DLE����>�˷�C�$�ɸX�C�G�Sl�&�:9�^D�	�!����"1us�E���.:,�E��eU�œL�����<.�X:' |O�EX!��/D�pe�՞wx��F�~:��@(�f�1n�3��T��f��V�%�=�V5��o*"{�,��Z�ѳ�F��\��R:������{�}
=9�G�~=�1��N����"��./��@iXly|qA^WS�3�j�[%�V�z}�G�����1
��U)�Y�q�iRę�3|8Ì�+ Q���b'-�,ƪw�I���ISY�tkG��5P;�ʑ�%��Eko�e�:D�m"P������Y�`�{��J_WO�j}V��f<�tf�����"ם��a3��!���P�6��"�Kݓ䯀,�%�9�ֲ������郺��J~�`��tǄ�%���xc�sQ ��]vt���,���I ���A.x���:���b�&�R}�al ��UxΈ���.͍G.����0�5����"��
����A��Q�/���f;V�܆����Ai;������=u`{����[z�KGѮWL�3��c?�E����&C�����z��o8,屺������ C�	����%���ۣ��W����$Q~z�-ŗf�%O�n��V�/��hjK���r?~��pҟTXa���ZV�V�rВ����m?�x��#�U 3�Ζd 0�?h�Y}��=�L��i0���?l���]�_сL4�DSD^4z�Ì➏��ԴN�w	e��w���2�����X�B yW�C��-#F���J��/t�dR뼙$��D��K�0qZ�|��-�%��ӱ�d����#=�gA-����b�-��8#��2@әY+�Z�����!loو4��i�+���_H;��o%����>�(�z�o-q�(0��`�H�mjw�����X���p6�1�j��ewe�(b�=h�Bs�D�dG֝P��_q
�-zPM�IA�(����LS��E�1�_3Q�������JAb��,ُ��+(q�-ra��!1�d��ل���)/�ؗ���'�I�_�w1k,e�e�`��&���:�ᔓ��}WV*_�yce�\C+��*��qE4���دL��h��^���̂�=���B���i?O�`�\Ä`tz��Q��H<V��ŷ�Ӕc��л��*Q0qUߺ���XV�����$$_۸|_��Nʭ�\?��-���7_5���7=>�����:��\.��a��C䱆�ӧ�V���I�S���:��rPITk�Uai@���A���͒�y��G�$�jKc�5��K\-\��(��.z��`�����~��SȊ�I��g��/���fQT�.|�A,7��^`{jQy��5���
�#)����{*����
�ӿ��_�T׈t�,���T�xR���V)��Iq����#?X���Ȅ�]2K�d��2>rjh!�7�t��،��������$}��!����a��R�G+U4���g�*�}jx��W�$��d��
,4��HIvěż���ª���E����W�G�����r�r�F�m4@N�0��&�*��LD���K�����lD.g����h^�&���D�d����x�eh�%>�'K�t\�ᕯ��({�pu��~��䈻���<��N!�ڶj�/�kb���"�A�7���Y�q�N@ثU����6$gzۗ��������Zծ�+;���m\��,~e#+
���bܶq`�����Vı��͢-יg:%sŲ �N|n���^�Bu���=_~z/%���w� ~�����j)�;�L7�&I���. �Q�ׯ;�?W@h��xکvf>�t I~�,Wmq�����s��ʡ�kzM (�]�`8D���"�̑�|�������z�;[2�d�-����v|�;8	���/i\ZM��+譬�)r�^��XЙ��@�l��Ȏܶ��*�����phn'}�W���h���@�1�0�UY�Fb�|S��y	��;5��l@��@g��@>��"���MD�	�)J��L����gZ�w�ƪ<��.�o��T_�j�а&<�u��iٌ}��C������B����is�

6�_kmV0s�>}S�uX��q�p$M��7_Ĳ���,�~���`^ly5�U�x�{cʹ���~�m�`m
�.�>�I����x�z��)EzINf���n`�p����_'�+zpp;�Ĳ[䦀K���5* G=7ۓ3�Ưu��T��e���]�Q�f���
���)I���M6߼�� @�W}��A��.�v"'�8�ϭl��^�l�_8���ְt0q�LK o`�]���k�7V}�OJ��
���3�o��q��Y����T)��W9���RG��˟gz$%r�N�P��su�y?��'#�~T�H>�����W�0���WC:�Ҽd``V?���?��9��F����,+R�-��wk�s�-T���k����*��sŏ�����V��ѫ��0ztf����K����Y��Coy�x*a�YIҠ��ߊjj�|;t��{�(����/l��[.s�iʢR���e"/�H������Cq ʝ�睙 "�$w_���JW��m+�c������*5WR�ٮ�y(�P�A �>~4n�6��)�����ȭ"��K��\J.]|���F!u!��\�wI3N��"�Fş�+���P�j�%��L_�]���]����E��b
[2o-�^��(�0X�ԅ��Ш��+1L�{g'�|(�H��]|c�y�GR�݈�l�k��b�"$��&��+��LFb:��c�$h�1^� k���V	8���.{Si�Ef`!�!���ͅ.�͠���Mk���T3��o�nه�x�Σ �^ka)L�,�/s�$�_!�.T��F!�ؕ��"�Z����(�C7vR�b�}� �:Η̎Y��S�q������$Bf�R����c���v@���Y�+�;�ax�����XP[�$6,�' *�z�5��[&7a3�A��:}S�e���U7	c��Fe2�w���m�����[~���3o�dGѠ	0�!7��䤦�W��0���ф�bR����7��$>�wq���X���nW3� Z���
��M(��ﾭ�3����5q���� ����g�g���F�?w��@B^VI��g�ei���v1@��I�Ԉ/��Wؙ�h�#�TV>c��f:�1��|)$�&c0�u������o���
���"�t/�Χ;�i�K��=���Z�c���E���&���W�#���^mA�g!�}F��i�1��cIZ뻹{�^j�n�+�W�!~&�l����_�^��m H�t����f�e�g��8wb��sBN(�@� �V��*��=��B�����S�Ԋ�˕���x����e߲���q�U�n�6~����,�W ��UC_��äQ���Kʊ@zy�0���ȥii�Wcbn����Yؽ������.���jP�2#վ�'I	�eD����|i�"c�[�*�bay�TqT��5uc	~o�FI[b������cL>$��<y�Q��Cӥ�yeL�Lu�ᵿ��^×|��!��m�[c�}�L<��đ���r��x���d�I�bb�\Ģxݑֹw��I���JsRu歏Ugh���y!�=`Al���ҥD"�4a�\�'��4�\�҆�<�y�Čh��w�	)��T�u]���k�c��y�����<y��xB��e�6��T⚬k�PM���qV�+��w+�th�	�ڸ��+���]$� ������k%��ڕ�g0V�w;���4:=�+��=	t�.=o؂���:��ZΜ���v��B�cǞ��rM�t�S7�@�{���u��	��SD(I��7��~�Ny�W�:A����U��_<f� �J�{ɉ�"���O�K��2���D6%�����
�?O�,�Zj��3��ve�	�z�&�B4�u�9~2��+Э�8-�h�iI�9n�9w��\��
���PODY�~x�����3ز?��:��~�0��h���5��m�[�}q����{<0 �,2�B��v�	�b������Kj��)�j�ٴ9XE�id�v@֜%�s�C��e���Sz�0],iW#?��(�j�t����J|k˹2�ɾ�T��̛
�m�}�H,!A=��p�áz�U���?�<6�>��~3fX�$13�*�q��4+du�#���Z����nwT+���@�9�y��Ua�����zC燣E�:��{v�Wt������>'���������Po�aD�Lǹ��b���|���KA�%S~��i��0ؓSnː�h=�7��\]��R�=K)
�<9����,�	�_]0�0��}��'v���酾Q���?��2���;%��O+����I��DK�9���af���H������SZ��z�$$u]�L.�5a�`���A9M{��g�٪�k j�{�^����T��m�^xn��")��9q�8���R�L��0c��d��\�m��&ủ~] ��l��ⷠ ���� a�[4c��ι��h�,t@H2��ވj:���+g��v!�x���*�
�l��p{jHw�Cb�@���@_-_�ԋc��_l����8�����#���s��*�bK��U��p�Ҫ*\]�����j�T�����F�*��]���vE�%�uO�O��~���b��Ad?�r�4N���o��x\���<���L��ʤ[`i�:Wqn���{�c�N���.�����"��Q���[�K��U����ATBu�+��^xI..�PiskFj��;�zJ��r�1L�Ѹ�
�^��c��K}�7H=�R�"xhO�r�FU���,/ֱ~�B��)"�X�J(�Y����,���/���ak�ťq`Owfo�K�)��z�`F|��=����r��j��g����ćl�^SqA8	�QxD��i~�2BDv�ֶ�`M^�R,;L�M�t�U��dP-�K��L�؎�2D��pvű�^�c1�y�I�� ��ҹ�4��Ѹ�`�DIA:���'`/�����l��̊�*���`дnY-J��ZG�;v�+�:\��wz��G(V��k�<��5a�nj�c���Al�` ��~�#��(���05	uP��tTZ��8$�Pn�X�b������p<���7������[��6}]�M������2�,�Q:�����Ϙ#2�KN
����k_�\7k��Mlԓ�󨧏��M=n��|V:����ֆCx��oS5\���i��&Z<����ُ�C�.��۫�x�_�:R1���X���c+	�6���'FrP]��9.
 ��o��~K����E��(l�����X�N��
�s��WC�����P�S��/�ߒ؉b�۝$�cs�Џ�s|�G�(I1����q�;��aQ�2��@�H�4�]5�����k����#�\��K��^o��Z��-�N��	�>����xBp�����ͣ��|�2
�`=)9�3�H�aҘ�@L>E��6�&�A���rW�_rS�y r@�m��t��j^;����§B�\�*/Ri��̃�ʂtR����T�����>
�&�f��
l%{q��Vd�11w{S�8p@a�(pg�[O�\�K݌���JM�/�00$��I1c;\�p��汥h<	2� ���3��D�@���>�C4$�(��٪��4F�m��FY�1pJq���O�R�������o9��9�&4[V;�Z8�d5?�=���l���3A���/��$b�"�݃T{S�I���gX1L>S�B�\�?ю&^O�Y���m���Q0Е
�Q����G��0ޱ�e����8��<|�W�:�9p]��Z7�<�ԀV�K2��
�n|`���Y:_pVk�?����6�DɭSX�~�p�yy�;��jU�YM��1����E[��U��JL��
�7�O�2�-b������[3p��\a�>�7�c��2�1��MW
�Z7�]�N�M��zqX�	C� }\�[�Otܩ�7��c5��W�z�[�vq���lp�&��%޻�B�+��[
������7�V�%�#����Tʚ�?wBx֚�C�#4���K���x0)�4pYQNn=&�gʁ=�N�Hkf|�N�����sU�f�꬛�ݧ�2��3]V�q�Y��l�`��������**U��2��f��v���Z��J9��]	�3
>@]>/񶗛��$� �z^S ��Շ?TX�G�1�� w]�eYG/B�)t��F�Gb�42ڏ��h�Z�v������~�w�0���)Et�ީ�92�����6���0�p�ʍ�L�{V[�Ll6t�'a[���
N��H�7K �qoц��7)��#gQX?@��/����X*����Brz8��,Q�;�#�;S�0�2ek(̼{E69i�Q�#Jb>��O���� ��ٸ�p�&���;����Sk����2R����6��z��p���3���S���tu��d]��w����i}��2~�La��������dҧ�a�����DA�k�S6��X�[Agd��G(y�� �*+T�t=~�G��K�*6��EB��(%�=���$_��gK��:�S:��	/�vr��C;%~*C�,VLE��F��X0e[:�EP)ձ�+{��=,� A�٨Z�u�i�!�;�Y�#Ɠ�nǇ��$�9#�Q�[��z���U6^�����֘�*
��C[���x V���v4�>�^�6V�rK��{/�j|��Cr�s�Q�������X�2s
i�$�����%l�])(cy��Je=o��o
jFO�.���Q��m�mm/��hlf���Pҁ�%{T�3�om�/?�o�+����Q����S.�4����C�$@��"��y]HOƨ�{��r�|[����XML��4��!&�l����k�u�`a(M��^=͞����������ֈ���o�Tȋ؛��Y	ZeirEG4�(ݡ�~E����Șj��(�lu�k&L	��!���l��pƨ=�x���Y���U���M���ԚSRxR)?�$��"_>����Y�=]���]:�"����.m��@^�'�v;��`S�oS��ɩ�9A�F�~���V��,����ב)��+�?� �-�bt�I�Ⱦ�]���涵�X�l2n/�.I���DR~��v��P���d[[�1�պ��}X߰� �VX������
x�=Sp U
s���:5L�1={�����sC �2>�������Uk�tWo�$���{���Z�����2�taB �&[d��G?@��5��dʨ4=��h-@����i��m��_U���	���B�0�#R�כ|.Z1{�(�[��Ee�ۂRW ���	K�=�����TW�NN�&��&��V�e����_��:�ׇ�U���_0���S���h�Y���:	�G�Qy�~A�A��9��o�%\�b� cKqͳdp�s혯x�M����)N�T���f��)�q�El!�z�O݅_�*��<l�l�{�����C� i�~|N����q;���V�v[��r"��t�Ί����o�2N�U�F��T@0���R���),H����ݞ��#To��
�;�h����AZa��.�D8[�j��0,O������vv�Ғ�#޴k�̦�m���~m
�u��V��|�<bH��ՉT��$�+wٿ�+�Q�Gr'���a�x�W��իM�y��M�5Pe�P�������\È��W(3~��)����1���Ս��ˈU���H�����	FT�_�A#df.���s�E\���)3����$ ��BҺd�&u�x넵��J��.��L�{�\�Г� z�������^�������i�ҡ��M4_��j�� h���N;m�2a�y}㉫IX�x���O�\g{d��9�Xa	)����X�Kը/���jնh!wx����+��)a��D>��7�*aۿ9�'Ʒr�g�����.�_ȱ
M;!x1���ڷ4]��ѓ�ه���.B�AЪv~� q9.e��R�0����l�ڥT�C�X�hH���Ë��U����!�n�Wz��|����&�*D���;|	�^wE��~�ז�M,�}�I1TER�H��|��{��I�(�4�p��ޢ@V[&r�T�i�D7;���p�H$xiq`�%-G%t�38��2�>SۑG{��]� w��%VPƑC�d:������N�<�0 �q��:g�rd/�P�[�F�9���9�-b g��E���4���Q�F.��Q��(pD(ʐ�S#P��Cs�y�)1t/��Z�Ѧ[���g�&]K�yڪ����+�;�Ɔ��kR
���J�'�K5��nu(�{����7"���D-���|�t­x-��8����:��(u���]�u� ���u�e���K7�̳�6��j��[K>�񚍼�w��"�KD��#�ekX+,~j煇�J?A�������cP��-B󵼈p����w#�.��^;π�m��k�Y0s�Z�K��\-�ᯰ�#�g� $�+����o��A�rPT��f��e0����v�)A����t�����)����VZO��/��N��C�Sϒ�$c*�̓�N��2�?,�O埬�my�k:�`�r�6��@�B��(z8���@�}��U�����r �8�x�6��I��g(Av�����6 �K��R��e8�	&:���,����u��tA�����@��(�H�E;�D�De�>_��üo�&_���g�-N�Q Dh"���@sT�$+\Y��cU��YTD5�2��\�[8W��vq6��M�Ya���D���0zw>wa��9sǂX��	?K��g��G�Kh��B��>��ǣ�����}�mZy�JyZոU���^�������̼�ZrZ@`ؗ��HC�hT/B�,[�.֢�F��WdӼ��]�Q�=<w����h�2�O�c/��D��c��idk�_m�E�sc[��;]z(�������l#d���Ѵ�M��݄���} HR����/q����Z�P�0�F�?��:w���<b��x�K�qh/kZ#���c�B�p��gg,ş����:��y覤o���|����h :		ث�j�]�|���5�5x\G��ËS�.�cᷨ\4U�0�k���(�壿�}��̍��P�w;%��x�~-��+�H�8����,��c�Eo����WGط��4z�K��qJ�ח�����<򌡸�r�=��3���S��	L�	�<���ᰵ�IG�;�;�"Y�Q����*'��yo�z�����B��8ƥ�*(�|�*REl�Ý���)	�Q�Ξ������#6Z �büt��R��Q6�C'm"B��@��QfL��g��,<���n�XS�*V�� �3 �N������ �Қ�9�8ЊrRe������V2��b1����NL�l��
���u�(!e3��_�G*B�A�����37�0�����gc�f.�x��q��щx�>�Fr	XZ�.JṼ�`���$�ԕqR��Z��k����X��N0�M8J�z{���\��3	�� R��=�o���M<A�$1u�K����*��_�KsY����`�Z~��(�7�cO;y�;@�AY��Kݴ� �u�����+@Ɯl���WE8Xt����ڡ%6��l�T��z��.�ZL�Q1�Gf�������6V�+�#& $�K�I�������}�n}�@Z]�!��<%0�5��r�3�W�q����P#�����%���8s3^���u0�w��8@���H�o<�y�R v�hY���<J�i���Dނ��{TH�cғ?�؛"�k>�_�jv�B�K=� ~�G�������њ��T��%t�MQ�i�e����0��:�v&�,%���z���*0��5/�z�j��Vլ�K�/I7�:�d��kV1���b��w�"GKU}u�"mY�m:%I e,�i!L�S�g5zy,V"4<9_h�(\����ۤ1���[qPWLx��ZyϿ��j�"�5�����0�� O#��
ئ׷�P)tTA��p�~���������*��#`�w� /`\@�ס�:�C������Z]N:7���Hh$ �LV�{y�UV@�6���Cm�^E�6x��Ri��҄���;k���q�Mԣc��8t��	c�R�Z��Ti^A`����p٦�F�g��j�`�]��|�l�|�_t4.I_u�ӍS�C�_�4���5�k�B��fB=���Y��3t���'��+�?-�0&"]�(���z7����s�߭o�uPp��^5g!מ��YE��z��#�cS7ϔ���ۗ�2A�Ѽ�,m ��r�j�7!�hePCP��e�n��,��J�hn�tX�ک�-o����\1��)�����ZMLDS��3����J��cd��j^D.q�A�h��������S�3�� $̦��d+8d'Li �pc�b�o�q.�+q��Pᡍ:D#5���r����A�"^��U�P &Q� G����h�>���W�����@�|f�p�/H{�_U2n\�1Yt5Y���ʖ�Z��n6�x��8�zld3�d��T��!��m�tA�7��8��5�DI�G!c}��~��EX���YQ�
'�#.�<�T�t��ML�@eLyү'������o_!�>�����]T���+l�.�p���ܳ�X����Z���=(�N�\
:��}J�-�e��Ab,�g��l:��ư5���"Z�e.�7�����23�8����/�6Du'6���ۢ��(�1�Д
�9�'ϓ�G�ޥ�|���k�\�S4��'�p���1{pa���6�	b� Jv�����5�.�����u���=���#�R~���I~���2�!7)hr�����5CVuP����V�]ȏ�F|r��]H>�.�.��=;�3�%�5@��Y;�k̬�_���T�u�g1��χM$AF]Gw��"�
r�9�ct�p�/��C&�qɾ�M���I�+rC`�%�܍8U6�>�W(��t-��2��	�i-c`���LI7y� a	<r�����3e5�S�
`#^2���W.��l���E��:����`�j�vGxվg�B�ݝ���b{�l}=JtpPV�됰	*n��6qmI�?�a��k�V�8c���a���ցE��q~�u�T���HT4`�B��.y�9���~ܴ��:���.s���CД	����&�v"D�\���}���'���dP�b�J��w���<��QX���+L�V���+b?�=Ў���0��	�f�ɏ��ߑ?��a��2'B�-�靪��0G�(��	�3h��)d�Vdp�1�*$ʆ�u����A�H|p �S9N���hyO\4Y[[�6",�0p��qlІ���&_e$9Ӽ��8(g�{���]3�E,S#=�~l����?�������J�x�vyJ�x٤׌�Ĝy�+J'\��[\�K�VSa�Vۣ���oX��o~}���"b̈́0�@͞��]��"Ft)�(��z>>��t���q&7��S��c��F�B3��X�9�[^��<׉ �:�u������|����뭜yPON��q4^�9�L3��נ�[[d
?�ٗ����394ޛY��<IMdA+�w���[���%�p��4M��b�{�����D���3�<T}-���[1۟��?6�+X�X�*E�h�A�$Ӧf��	�%�D�[Ia��0S���q$
�[H`[�p�͢j\���KE���	fDU����d.��ňN0��d.�cVAUp�_�aq��!T���=����z7:�>1l���C�IϚVo��}���Һ��:K"X�ԀM��*JSe�_;���, ƎV+WA���Ӟ�xjk@M�t�g��{޲~�_�J���5��3���MgQ�� [s�B{���hhj����#h|�f͊���/++n�&�ʋ�!['f�
��bQ�x�������H � ����)��{Fb��h��$��bOɑ��,me�9~s�ˏ2�V��g�M�h���|��׫C�)���h�;� �,�	v��^�֭�E��8�l�z�V˓�֤g�����z� �2��|>oBe�H+%�� EM�NH0,U��Fe�i�'�U�׽��v�
�9m˹�v�݅_���

�o�h,'謯�FB��L��=��y	���%�Z�<lߒ��/'@Ȏh����n��(�9em���"P(������?ww�0���n&���e{k,m�n?�w ��7՝�g;��|Z#MI��Z�R
[`-�V�VT}�Cv~VJ"v}	��-�P�
�ws|s���]~v#B^NG�R�t��l�}�aj\쌤x>�Z�Չ+�_���w�|{+n�-�.q��o��\+���(\,y?�x��M���Iu�O�덶��i�܎�\o��7��ʂ�}b~W�n(f|�0�㥺G֒}G_���'���&h�Ӆ��l��1� y;Y&�N����YDw�I jN�����������65�UlU���6H��F�.=h��w"/Z���SmU�Z&_�zo%���{z�76�=�:i� x=��}C�P��X�>�p��`�� ,�K�&��.b�+���`F�+�M��(鏜D~�/%�<q6^���l]y������:n
�����eu�?����^1٬lũ�V>
~�&��^�s�9����Ox[U@7r��Ծ�7.��
Y�u�dTb�A|��Ӗ�~����{�|�#c�)*�2D�e��eD���.�P���ėaRʑ���N�[$=�<��cM[(JAN�`��6ūRA��k�{�IT����}C���p&����9�	��k��ځ�VRmN���q���L.�@G����fs�Ռ���bA����`e�������VǗ�h�b��Gl9(iw,�icMA���&����dX��[��o��'�;Ck�	��)�H��0 �=��z��� ���=Ȗ�`��W��Ì�Ƶŉ����w!�[@H��W�uq�	V}*F�J�#h������Y�8�nB�iHK됊j������&ƀ�VDL��J��")[�Z
�dp��(�,u��%�znq�1���)!�O� N��v	+�g�f2�*�T=}|�Z��[��9��4���T�������'�J*t����@����'�`JxJS$H�*-����ib�o�Վ3�����] �����'����묟Ǫ��2�Ҥ}�S�BN�T���I|�x�5��-�Y6a\T�!NMp
á�I�6���|f��5���=*��;��p%*�9����n,AW�'�����ֵ�4��r ��'$X/B�|����D�!��4^mj(A��
/��n�(C�(�#kQƋ���K3���ޯ\t�﷡z�}��yV?<�Ψ�&yȹqI�K��}9���7�T������p���"mKa�F!��`��+"7&��QwI��*GM��Y(��7�a*�<��k��0�����<���j�W�|��7,\��z���֟�zo������N����F���YP@:ón=d%H��_�>�p�2�h8�$�Г�7�.��}:P��R�2n�~���M�\0.��H�ů�.Px8O;W��y���ocu�z���iݿt��N�KcKՇ�
��@Sv��IC���.�O��0�;�L��I���q���?�h|��i\3�\�zH�|�x��Q++�Y��=�73����w715���X��SY�~l�P���J���J�H�*'�����3��Z��L%֣�R'�${�/��ak!���;I Р-i~���g�"Xb�o �������F�)�R��loWK!R�M��ݎ�E|z�,m~�yF���K���]���~��BM������^��9����J��ik�V�3�D�m>e��J8U�ʠ��i�5'I+�c�غ���w��
EV�x�e:�B!�+�X@cW�d�U��/��o��T����S��+���wt��N<�jx����N�?�k�R<~�B�M�@�0�-�~W�4Iqcf��ٰPz����!�p��F�W��d�k�P��x̗�m�fͦ	� �qۋ�.�4S�v��r�n�w���R��,3_D-_�+�����]]��-���&ͧ����!�k&�Y����!/G�D2��:���_�-d
��/5vOL�Mx���0\�5�4�ԫ�ɓ���ʃα���<��蘃��6�ۓG���b,�}np�vʰ��	�G4������������<�x��Ы�B7E�P�ƥ.��r�r���m��G�
%CBg3<�̝�_����,�
�~�Z����e^��h&)5��k�*(��(Q�I���5�eF�����$>nٸ5�:Ű��Ty��Jd�B�E/���PpX�����FT�Ӄl�k�[D{"���m������	,��XL**u)K:���$��	�?&��C	��g%X�Rr6��c�b�K�hI�r������~c��J��̣JOi������H���,�!=���Y�^7T��q}�"�.�(����Q�X��y/�|1A��v��̼ee?�ģ�)��iå�K�y�������kO�_w �%`�Ii L/0bNy���<����\$?j17�(��%qJD������N��h�x�RA�U-?Y�l'|�JS�+8��<��ߋ�����|��t�3R����%Wg�K��2�i�ݳ7�R���t�>�m��x��{vjw�����l� ���!f�^��Ə�$� ?��q�q2Ao�����<�-NO,���b:�|V�G̩T���j���Y��-���KUߞ���zw�L�o�!NI״Sy{��82�Xf�������ު��n��*���Û����)��pں�{$`K1�y� �����%���s��6IN�Cv+M�Y9����8�n��P�mK�RH�h���-��p#f���)Q���8�H�������m��p���e�u\> �$f=�.DĶc�!G<�)����H^Zs9NQ�Eu�u7�CM�c���.}Ƭq�L�:}�=ȴdϭ�h����y�GT@�	��A����/t���H��*���Ѫ� [{�����^��N�B�j��H�JYG����_����Пt��q�eyp
����B@�#��3h���Y�Ƹ���3�'�jg�k�8�����֑c6��2r�$��9�]��-�x�m��N�x�N��:�8�B�o � Ƭ�EK��QЂ`H^�.��jI �)� ��w��ޮ�ᮙ�^�'�0�M�����TDmbu���q,͂L�`��`�t~{���Cr��Y	?���R�;�`�]:\I9���"QT�v�C]�� 8�YA��
?�ӛF$�@~-|�Z�bp<�d+��7*�X���9{�Xơ�P��l���
�JU�j����G������6��FX�*�§(���{y+0��ԔRr���P���"�l.�����Ђ�QE����*���iܕ�"2_M��t 	�Q\����Zs�%q�I-m��S�VD�zS`�@ʢ�2��Nug�����Am\��q���}p��v��~��q�-��^ȃM���0�#��|�y���S|l#`0Gѩgdk���OBőo�*V��"��Y�F+����� AH�7;������}n%�����mT��-p��$5�P)Y�Ҷ>\aU'�bH�;_P?���� �����_hUS�L[ ��)V�p�l�����q�_1�!Xp���YA�G1U����_Aצ���mߒB��QI׬�nRD����#�7l@�M|Q�@K�8l�9����1��({�kwM��G�jiBv:��h<�v���Kx#��F�����S��v<*�D����Q��JٯA�^��ѕ33�y��Ε����o9\+�n1w�É�[i����'�/��G�25Mu�y�_��{Qw��<�n����ύ��<o�3}��U`���B����8�^Uf]��s�?���g0��mlT+���F���ui��Q�;�1h�3yhm�qt�Qp�O�h�P[T��ޱ��-�PRE���K�s
\DK��v�O`��U"t�T���lN�81�	�����t@�i�Q�tN`�s��ΕS+ny��g�^^��k��(���\l��������ê�.����/�[սS��b;��e�fnZ���,tx"S
c"��z��_�;�ܙ����{��U��2)sh��9)��da���`��G�e #s6��gt��a�}�*AP��_�h�e��3n/�h��:+�H�k	�j>�QB
z�����.Qy�Ǚ�4�Ď%Љ�&��,�����O�ci��!� ��h7�w�:(r��E�:��Cu)���