��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��A��T����,=?�����G�F)4cf��4�-�#�	¸���b�ntV,��q�~�-���M�c�Yq�+�Q{7�O��a�{,�|���.��J�� T�=n��OLj(���l�|��u�^����^���?�����r���HQd����Eg4�h�z��ݿ#4
�ŇPuO�|���FhU��SU,�S���p�kVb��*KgL渔p�A�P�g�ܡ�:-c"�t��j��./��$_�4֭�.�?앂�o�LE%M�G�~���4������YUp!6:�՗��]D��}�O��Y��K��m�cеz.ٲ�KU������I�+gS��0u�D�%�w��.9ҹ�R���^/đ�uzq�kt��d,�*ފ	��ޠ�2��5�O���\q0f��ss�s��.�>�{�DUQ]oٖd�S�O�1��;�#Ā�AA��" ��Uj`�^r������_!�y�όs�-�J���0P`9�gCh�q���%������?� "@9��)y�\rY���
��[Y���7#e�#��4�"�pZzt*�h������B�ӕو}�#�}��Ⱥ��Czz۽U�ʽir*�N�3Gz+��/G>!z������h0���=���I�"8�Nn�� О��-�ŠK6!����#�C0!|��,�jn��#�d�>v#!���A�	�jD	{��6V�%%�r�B �i��d��z:1�D�h$��^r��'H��`6�\�$z#'JNa�%Yiu�o��Q!�6c�<�m�\կkBO�>��!�E�(L�x����Wզ�L��"�!Sb�=ȫ~�Xr�M��<b�aTN���#��A���J��K���|��;�dQļp� � ˂K���N��%Y-l!�#YM7�պ����5�5KA��0u7/I�].#u���Mͦ�O��\��g1ܒ+CY$/y����9��Y|��`�fQ���P^C����`D�l*X�P*��Ɉ.��_����2 o��?�_:�:W�c����Nu����w��2<Ϗ&���W��M����+.Z�1�Mɺ��x,����� }6�i��L�a]���ZŲ�%�>�aI�����+�-vS
6�����Ȍ�M�lY��ɕ6<�.-��V�cG��hľ�&��Ys@"�
/r�+uM��1 ��Kp�trz�w�rM�'�ϑ'�NIO˫��"ՖSJ��>ءG�n' �6�hX�!o�i�WK.Ò��ך-|��]&#۸�n`[�.�@^��*t��x̟fY�p�5���<re ��؋R�������ܖV����˚6Ĺ�~%���R���p�л�5H��q.��d|}�(bz��5��q�4��l��ii!d�[iBtjw)��RcJ����
��u /�?n�@��lT"Q��p:����\�b��}��nl}J��������m2ӣD�-���x  �r�w�����!�K)?���� �q�ȆI�ݟ�4��֏��V�6���f��j�oh���gP�(�����I�V򞛲M�]R��8���]�����$�z�4GsЋn΄Q�gt,Thz�MZF���ew��q�F�Vic|�v�g�DH��u���t�_w�7����dR]ȑ�isjB��~R��qU i��8F���
,�q��=z�K��B�"j;;Vq�p��ۼ��=��#�9ٙEo�~Τ߯�(�������%ɺ�"�N����s�ß��^-�8��֜`�D�0Ʊ�*��,�������3u�"�������
IǊ}1�Z�W��r�i��~LX��T޺��@��W^�����t����"f���ud����N�3����"/v���p~���qg�'�B㰏�ˆ��<�y��i�1����+�N;�V3��Y!�aSCʔ�9�
�~�U��C!��N��x��^/�Lo����K*'ee+� #����S2O^^w��'��I�쌁Ӥ����m�oDgŤDs�F/�X����1��<���@�f�\�+�:.����y��.w2� ���H��,�V�ܺ=�>��՝��H��?��r��69�W�d��axD�cB� �!�	\�a+8Ț��1�"���և�9V�H�s��ͺ@�3�̒&�%2
&o�'d��.�1ұ��-�F �!�޽�6�� ���&b|�c�J$�BEAr�m�)�i�ъl�@�%Z1gy�0�$F`ō�$�R��ut��Q
�Fԙ8S��E֖z�l*n�����I�%G�=d'H�=�HnD�1��@2*�"Mv ����� o[s�,C����Fb�<f�c�%(������n,�5e���I_�m�H���1)b8�����F15�����3=���ƿ�v�Ԛ2kU�r=A��ḏ�B��0����"Z��$`� 3��xa�i������@�Q�q�[yP�6�U������ $�/�6`��I�h�OCt�Kc�j���$����hbp�!�|N�~�OEE�6+eY�82+t�"�{��A�I��;�Q��o����2�rIK3>mzP�UrZ��6@l!�m���IU�7�<D<챐�42�����@�c ����MV��V���f�k%��qO_�W3���Z���1ƿjrK��A6:T�.���)N*_�5Q���wd���B$��>�N^&2�����(�t�G��Wn��2��$��Z����;���f�������^@Z9�?
��8���Pׁ5��1���uq�.yq�2����yɨB�˜��!s�0�qA��[�?M �0�����Ӳ�ŉ����R�*<xR���dӍyj0�iS>;Ns�UB��wF� �G{��U���~s�NH�b\�Bb4� |�B�& @�
l�~v{�d/2���ˊ]�m�N��H���*�A�r.qL㣟�����5Q`%��(�K9?~Sa�<�Q�0-�׈O1b�Z��a��	�g� �\���d��Y�� ���{���zS;��쪻��^9S���c���D��_ӌ���t$�E��*15^�/b��5�z���v�)�����Կ���e�k6"��K#��:f��X��iB�+�O�h��#	5�Q������"�+6Y�2g��?�	EC=gĆ�U�WXG�!r�^RM��ǾT.5h�O����=O�0'��6�X =�Ct?�1_���)�'�!.>Ƕ���m��[�K��4(�ʜO&ܯ��'�#��q�)����O�z��wa�l�JK��b
*3��J�R|+�pz��s[8�e�TF�!� Q�1?��mps%�L�;r��1���S_Tl�=n*
J_�>p74;��uY�h@�#hD�����dO��']�($��i���bXjk�H��٥�w3}�`����Q�׆��F�����,^�o���Ԃ�0O�\��av��8�AB��td��
��E�Զ�$o5���ęhs�g��#�j�+�<�V݄ZJ5E���:?�*�$������'�=	��\BQ�ls疒���Z��ƅ�{����4��T�������y�v����Jg1o�-(�#:�FѢ?�m�����;Aߏ����ޠ�I��V�w}���*�yb��I)n�$�oL��K��l׭p<��E�]��+]
�~!���?��X���>k_a���(� Y��т_c.�"��Wɖ�BY�$;P&7��0{Z�{:�xeVl!C�;���眏3y�p\q'P�p�mhf���h(�|�d�D��e�"3q�i��]���{�Q9���R����]�k�#��:���0����,�7�ȟ&��D���L�TГ (�T���!�S�;�R����T�Ɯ!�&p��Cj�	��q��9����x�7��TV�w0�Z�c(���ώXX��/�O�a���FD�QA�ަԾ��\T@��ajX�"(���4Y&��۬��c(���y]���t�qaV��ye Ϫa��7���%pmw��0��3;y����N�U�U;�UqH�W\�;�����=��L��XCV��Y׌�����h��K0���9ѤlG�|ZL�J&�7���e�M\{��=(�=��jr����G��~�!J6��Q�_i12�Ąsv��;��nܵw�F��w���iL��0�cM�	B�!�~�b�&s`��*
O]��γ:p�Od|�/��n���S��v>��fI7�l�/!�4�%Ug:"N�^F��B�H%�|���W�2����j1|:�0������+��C��R�{�å����&f���CM�M���w�x�ʜDn)a��wP<������m�,'%Ӥ�,��7���Xv����7l�y�/��?Ɔ�t�<��^8)(ڢ[T�1�#�D�Y~�w�2^�P7�.㌂�Ϻq�͉��- ����h��W�b�9eFY I�	;6Q�6�L��n�l�`+��)D�G��> �SOY��$����_X�<~���ћQjQ�R�❺��u��Pȩ̑���i���o��l�xY~��|���jn�j�5��Ycq�u�$�󮮦a��)��c���(�����U���[������<od��#į�X�)//��xi�U��-�my=a�Ң��f�Xm��44\�6�����P�(��F�Fw��]��W5��@�#�I����#j6��"h�O=�k�f|�[��F-z��C���sD�������R�����B��^��8��{��A�gNz�?{{-~<f�"c�Y�{�ׅ���X�
?�<���*��������8a��F�%%�)�#�/Hνv�tD��IU�3�bE��)x3������_lV1��˶#�����)�'ƞ(�ʈ�GGl�/�fjB�ڸC^�x�$>r�-�ߑ�ۙr�rEƔ�Y&�V\��Y5F3��F���myN�Jɬ�if'�G0��(ቜڰ��s9������8t�a��9�G��t(��PdY�p�Fi<�K�p*�z�A���0 ��w��Xą�(��x�0t�����Q�2kq#�9[�����v$�6����Yt�,��Bz%�8m#+�L�chwf[��r�A���J_A3{p����*$��Jn����\5� �2Ȩ�����Lθ�����lufs�uZB+�G�د�H��?^�3+z�Eŷ�"D&�ڑ�pAcv�/��M���Ԫ��w%CH 0fW�>�ς�j߈�g���z]��R��I������=1�E߮=~��e�Q�(IU��e�C�(���eG9���x�GJ�������������0��H�s���%�� �����=$h��*�U�+���ks~���e�#g� a��HI�6�Q��?��܉�����K���'r]o*�$���({������`��1#�h��T��ϤV3����\(��p��_�y�--���u���&�,��q��~H�I��&���=�n�v>x�)���-i�2�7!���:ƴg7�e�÷���4	�;0�w�F7
E����c^ÛYm��,Dք�;ae���c4��Y�Hz%J���тg�	$��-)B͙�A��P�>�cx���{ܪF~{ᾯƣp0 �e� �Dnyݲ�� �����Ar^� �xW`ۭ͔�Y	-R,"�.��y�e���̫C�)uHXXv�	�i�-׫�&wڜ�@�U�}��FE(�e�� �yM�T���'�CM)M�Ьz� �>k�#S0S�vGҿ�E�΄���G���cA]^"�^Ί1�N(+�ԟ�BwV�svi��V�Eg�_Y`Ā���gi^|4�NE9<c�(|ύřM�}�5�yG�7�����Z�ǟ���������3QtY�'嫟�b[H���'< } �Bh���n�^�j�������I�`��f?��r��ym�K#��O*ף^>>�ѸR�Վ�b���(~l������磑jG'ZL'���"�C��v&����1Fl&h,w�Io��-�ae��p2q�����#���>���ݥ����?�u��(/:���5[}���� '�Jզ�d�Et�\H|~�$M�~ 9��W8� ��L�A#�j)����X�v�>�VY�����!���>��:]W�bJ\��K�-?�	a�3Bd�F��6� �a�'D���δ��"'r�o7�͇�>bcz�\�P�x����hK�Gs��㼀;���C~,��X����5�ɋ�0��)��v�~��X ��M��@V��f#FUE��ǎ�~�m��ʃw0�N����l�DGPԠ��h�"�
,���$�����0�&���Pa������p�]A4a�w���4���JoRUe��&�V\?A��&�a%���I�}9G��og���)B� ?�.K�d(�T�ˊE�<�ǫ����u+�����rW�����a�3����t���7�=��z��ʂ[��;Ph恴	>	�fnI��[��8[���5�'E�p�e���xqT7�rkUGԯ;�f�c�'���s��b�w�1iA�Sp�H
5��wm1�B�(�M� �c��D�����[��̷��F)�Hv�\��آ*���0Q�	 ��S�@�8�d\���3W��.B.+�F�K?I���j��'��>��`)�Y�-�^���YV4�&)�$�u�>`�A>�M�!}Lj��Tټ�v�j�C^�L1�_�C�thB^�e؞��яP铹!�{��i�(�ƿh|�.x?����F�t$a5��6l]�jFTO(���BC!�g�YEq,據P�ƾ*���*��9�J�Xb*�;���%=�S6���1n:!)��9;��S�H��S�sl!�eX�k��Sf�֥-n�~a���U.TI��W�}�dyq�jWv�W��+��]9�0�8Y�^He���G}��������+]�		 �6J��b'��U��w?v���F�Zh
�pL��r�י�T{�ʙFZ ͔�������knˀ�O��4z���}v�}˽O���W�	����=٦�󱒌E�㤷y4����t����2����]��e�.�~%iY�6e5۞�o�7�to�3��U.&L�d��2s,#��:����O���iY@���k]�%ՙ&��y1��v�*rR&��d	]����2�Ղ:񾠇*��a�MoqqCu��Hsz�)oB�-���<��<������cь�{=Qh�V@M��ɤ��
a�x��U�+?^��3slv]����}�C\���3 a������Z+�,m��-�X7��찿luP�$��Z�"E�6�|GR������A�7��
f��g�ԘJ����UXo��:�BAl�I���F�����[�_(��ј�o's�3�ih�e�Y�I��<Y�l��D	�i��-r����#�C��J��L���!d��(L;�d�r_C������w���J�:+�-��g;c�`�ԃ⑾�/�0���C��6a$z�.��fU�g��\Q�3Ә�j<����� t4��}$2�/�W�c+ͨ:�x�*���H>Q�t�g6����7�����������J�L������H���+��F�V��@�����e�
>�.Ӗ/T����9o��v�>$J�Hx�K(�TP��(��Fv���)����I����L��uv�5��b�x>�ⱀ%]x����fi��7�*{�:��)�	{S�
���7>,��G�2�~�n�H~���-
�_~X�8��sh��[|���{2̰"ƪB����a�>z$�����#�8HED)"7�{���Β��t�EC�J��U��/������֓���d	 ����`R�Y?ώ��Rj�,�l�9�ũĝ��	�$�V��$��Q��x#D����܀o����#]X�9���`��$lȵ�-p�ۭ��E��뚆D���8H��2b�� ��9p��3+��X��hƾ����[9�&L�� $���r,?��J~���RW��E�V̥%Y_1��E��-B��*���B.x!��-\���#x\�p��v�_&�hl�����'���f%��^�rI�e��' MB%O]�d��մ���l�W�~�����̏�nwB��l�S���15[����F���g5���y�	����T[�P���p�X��ޓ�7����@�0k�`������E�6;{��A�M&r�\r��&�'��ྱ�P��r%PP,��C�*ѳ�zzi9c�E}�Kٻ]I�B��Y ���U�������|�d{��w Z�Em��Ľj��qy�E�1�S�#�e�ΘLeD�U������<s�/R7�X�ɣ�1]˷-Ie�|��Q�g��T�T�!h�G� O*��ח#YK,=����e�l-��������Ai��	�*���1v�}䌠��E�ݚ�bz��Eq ����1b%��0�0�7I:/���]���W�OA� Ov(O}?�=�� m	����M�����6{�����mi��$q�ʵ��3^��Y�.��stn!��<[�z�!�7I����Y�
F��A���K��z�D�S���B�%���[���wJyK���z�"�P�
ף�_��'	���iO���0�g�BLr�ڬ�n�6 -	�r	,v�G�y��<x&s��wp>��5��~�,x�c�q���VcFQ���\�&lʔ��=QK�'_�� �/�s^xPϧ����Y�|�=2p�@oRaU/�M)]����{��l�ZzXL_�<V
a��O������F݆`�_��(�{n�皛pG2"T���	
&��	D�. �h��Q�O�|��4�b����A�bӵ���^݈�7�PS~W�,rvƎ��_W?y�^�؝Wn�/F�^��%��_�f�Q1���=��p�^O:�c�a"�b���������b~E��R��j#G U��T��svq��z&�O���6J���K�E>����3��Vno�ڳd��lԷ�mr�;O��KN:~��/.�s�����lQqj6�?��{ji��9��1�N[K��tB
	�$+�̃
]@��~���u�����\��/���0���u�����(�0W��/��礯� S;l~��z�����]�~M,�%<@�0��T�ҟлqs_�p�ę^�/dB]�������sb�Z��U��d�(O�>G��콺�k�F�}�s<LZ9��e�-�%q�O��|f�z�q
ͪ��c�<(x���M����X�-�;qX�X呒;����q��i��gf!���L�9:r���5GE�ׅ�}���)�"�2ɩ8¨�$;�㥤�Kg�e�4]�yz�Op��$5�����n�`��6��V�H��x��0��}r>�X!�d6h��[��.���L�d�꩎b�ŎP�m�QӪ���2�c�;C�D��f����a����C��K�5Cx�o���×`Ĥ�0�DΓ
�/��A\n��^ ��Mv��4Z��%�n�� �d�Kظ�� R}�O���ɽ�FW~�m�'`R0�� |�Zޭ-�A����� nE8Nٱ!]�3ֶ�xχ�������W;*�ur]���ܫ��N�@�'�,1���rL�&�|�a�srP�
��1@M���X&q&0NҚK��h\af~mVm�A�������%���4�������,�����U�����k�<%to��������Z�g31]�W���U�,ytq�7��XU9����!/�tG���L͗Y�f�Q)�"��p+�ځ�֦g��<��s��U�O`�4B+�`�t�Rv�_���+���ѭ�S0"�%���T@s�H�o�BǐN��P��k�6�'=T��~#|"N��c��)X!R�7.��q]��t�鑗��u�w,�i��$?$?b0H�e�ޯ{���>��X-�\��, �'�"|x�Յ=wӔ[k(�+�tCȒ��e� �i^�/�NAb�}ū��:G�X���+;�0A�6�s�]T���)3�F�2�8&��8������/y�Y�U5-�5w��Q⮥q�a�egn����"��x�@��_��"#��ޛA�q��ۙV�j�٣嵘y�����_�x�����0�f�\_�h2x�׸�Y�����G�,�r�9�Z}�'��s%�?���d��]�f�prX_��"�8^3|g,2Ll���xb��V��w�ę�uP����1�Nڒ�:��`lv��,N�X�w�f{g�q�^P����I
��A�IX�8jb�L�9a�G!�BE�m�&@ֈ+�Q���
dz�����QD���x���/Tہ�̟L��y7HW��#>([�+T(�����l�����c&f��/�3giý����W��V����jLƧW�f(ʯD�]��pM�=JqzXr]RDu/)��`w��)�L�DaF�s�7��\�#�I����\d������I"qOVx��uC� r����T���C��ʩ�a��f�j�y>L	32�s�5� ���0N�.��i����ţ�+q�۱&���%NԚ�NS2#�ɨ�i ~>!�����fY�7\�[���}��1Ymda���Q���d��ʌVB�<�Bݐ�n![F��Qq����_S["w�4N�n	Ȑ���L�g�o$��h3l1���R�)$��X5e��cV��d���i��@2�ئ=��SR��Ci��I:)�)�)��Miz�/�_g�/�{�0�4=4�U���cOX�%W#���/�C\wr�M0��.�1Nm�����r��oz�V�t*�ä�@mI��	оM�C=�ǎ���wE��W;"�k��2�[u��0!�iA�����?��d^���A<�\hcr�E�����0nu�Kb��5���.C�6��N��(?��x���L�$F<GY�Ά�����M�q���"/�j��K�\�������kV��TT��QP>�y��o��1�v��_z�7�I��p,teܲ�d杧�G\�4�4h�u��L�B�� 3�_���ɹ�+rx$C�o�=���Ӵ�.p=_�a�)L$î�٨�NP�{K�� �?~�Cl?pC�i�߶�d�3�9���Ӏ`�t2��]�ʘ�T5lΰ���~�ÎO<�3�o�rݖ(-����N�J<y�f�[���m,�m���$�ຎ�[nzl����!�K
0gy�@3AA(����O=����r���������C�"�E/�UF*����7Ɨ$z|��B�B�U������l8=T������2�������F�*"�I�N^!!ˉ#�S<I�]_p�d�����<�#n�@����Ee�3x�~	E���OA���]D�0���
W��9dǷ䶞�<��O��P;��a+*���\7���4*J�c*������xWRA���˘W{ݷ��j��?����xg���3�J��\Ai-:I~�xQL	�d�����D;H����tɓ��*�$�y��7��A������K@T�'���7�a�d��E���Vu$E��7o}�"~�Q�-;�%�}\�Q������O[Y�!Ur�p��;��0<k%!wf��*�>��V[r��	��g^���!��+�I�.�a�=ɧVF��ܽH���D�(��`ci1+~$�s�Q��QSL�ji~�b�5�|Y��n]a�F>��\WÑp���&�ަ��
BRq����j�ߑ���55dg r�W��d�<S�%���e�z���E�H��K�O�oj8�w�����4�(1���N�jh����6���K/���Rl���F.#���k�'n�������e����CE��xWTx"��\K~�9�rۋ
����|9P`����B�BqQbބղ4��w�cP	޼
I�cB՜O�E�/�҈+Fa\Ǭ�X(�B�vf�\[��wYd��H�+����U�Λ>oQR,)\�9(��F���sa��#N��\#~�K��22�d��o/�{�w=���0_�E�v	^�Jd!L�B��[ڰ���f�LNo	,���Ҽ?_k΍������FI��ck��S7.��v�,�������3?>�j������1pAn��~�4�v����=�ʝ�Wy�=��QOv5e��0kq��p�!�-�{	jgv��mI䛈��!�����sT�8n[V�,�}�f9t�D�=V.mq�#��
��*�'�����pHG�z����{a&�5�=�S��~Np,�N�o	��B��h�� ��]!��T���Zg��X�py�L;��6+�&R���C��jE�[^lū�X,Ax	��MX�m��pSͱM�����r� Kv���:@��ȩ6� *8��=j�zR�|W��6�`��2��C/р�y%5����4�Wh@�%L��r�7�[���r�2n*X������#�GĿ��������)��+�Y5�`�4N�!.��y�I���N����d9��3��mv�4,M���x������K̞�ϳ!�YM3�׵�|mBn�|�6�b�?åDv"BZ��bRF�����ləVh�&?�Wۉ��Z���X*H�]��K�p������$B�\+�r� ;���K$-`��փ��~��_!{�p ��;ʛ�gv�q7�?�
4�r��N.��Y��)HZ�3�T��A<��6 �wؙ��-
�ף��I�\YguQ�����B�Q��Z����X5�M�ԭ�3&U{��nW�A2;@�WB��CI��M���ĮZ��+�3�N��+�ЙQ��E�H`� :����Ҳ������p�:��T������Ύ^<��G��T�e11}Hx%9ϱ��/�������^�D㍙���e����z�$(Bku-_@@���V3�;���-{�o�_D����)��^?�0���C�@{�h�6��
${]���\s�پO����f6� ]?�U�}L1�^�E�.cX�Z��':��qt���m�xD���V��4�`�R;���*A�|@�n
�{2��|꿜E��A�m���(8\��{C���K$���d��_D8� ��q�-�W�V�I����>���y�m���[�pu��lˬH����$1T��>������ ,�e`,{��f�xH�R��.��v;������}���{�B�qh�fQvӼ:�����RMxT5]�3�l�M^<߶�����_:$8D�B��z�I�T	���Χ
��G��iD{]�?SW���i�?�w��T��唋 pV�k������(�������;{2i��<�Q��r�_������<��.��%U������l�~�Kew���N�3v��lT�9�����]�>�au�����H©I̵x">�r��i�za��0�mf�װ�� g�![�R��l��}���:e-2�a啐�.C}+����cCk�ڢ,M�J�o��:�Ҹ��Ҍ��ۥ�[�]@&��-���ld
�<?ªX^2�,����Iᔹ�Z���͗m-�d�PO�8PoA�1i�\��u"C��ug[.f��BX5 $ms{��zz/,�*j(���^&�Ų�n��C }|���2J��?e�ֱ�t��z3SPI�d0V�ǌP2��_��w�q.o�F%��h�Υ�/2<f?t�T_����܌^��$mwH�s�rc��v��B�����BlGkI����h� n��Ibv��.� `�Ó���8��%�6����1��Fn����HG��/y�s���B�qiR�|X���-t����K ��֞�N)[5w�	���gEWj>@��K+��$�)]��@� �#�3���S�[�]�j�`�����~)�F<�#�����ɴ�-�4�O]��k�4[S0�#�W��=������v�"�f��$>
a��X�<��\�i��l
gȮ����6�h�l���D�cd߰�aXv�eK�ZiD}Re�z���ұܿ��I��q	�����h�����0�Z?��b~C�1�)d�g�B^roI�O~L���1֑ �$���.y��A�WHK��"h(�/��S�8���\�E�{��|�3��54q8Ls~h�QJ�a��u"�g)��0B�v��[��)񜢷�੎VD5=�<����|�:l��)���p��h t��.ڶ�m�:a�lb?�>v���f���-$��@��렖,�`�xYu>�w�]A���E����q��GHA�̆�G��(�M��1�x�0��{\A�|��d)uԷT�MF' ��_o ��˶.��ߍlB�	��f`H�'�s���4ږ���8h��F�X�Yi��C+�j�+��fK�ٺC�� ���0�&��C����(x�f]m�MP�mz|����� SY�	Ԗ�f�+�_�/�7�I�1�~�{�
 ���H�V���x��R3�����mg�����W�"'WO�����+p�l�ڀxO�*�r|��)P�AA��R1�/����/om���P2��n�\BՏb9�:�.j/����X���x��G<6W��#2�6sR7�R��v��M������u�z~&�㆓� &�1�,~%f I�s�����˦�eU]$=�{�nb�/�Ϧ> {�bj���^�����P��i��6��iK��{z?c��r��w���Y�R확S�P��A���r��a������&Ig���̋���#z"I�r�d?�����=�%M�������V6�%� ��+S�
 ;3�����xkW3���y4�@�� ^��>��R�F�X׍2"S����K�=��N�OZt�MN��b�h>Әdc����u��ݧ�\�Pm��.�ffV��Y���p�	2/A�Іi��0�� ��D��P4X��@�wO��ۻ���'��4z�!�B�"����W�p	��0�sX���]��M#�l(鎃@���_[`ގ��d�c;��gwA�P��jܲ	l<L5/\���� ��iǲ�/�7����ϟ��N5��P��by��CH%�!�a�'�s}�8�C�e�J�8�~������*�����Uʘ쇖����� �"�������mn��U��]\I?��>����zZ�TcZδ�Fǁk�G9�˚��IsT%.�ő��cY/�P'����������vP������@�K�ښ�HlJ{h"0����`ڐә�DX�y��v\��O�J�6��}������4��#�Tظ~��8A��F�O%���� խ���y��D-���:eK,̴����yl��k]�9�t.����ZW,�J���.��C*��<�1�_fQqA5>YG�G�ŀW~3u�^į;�e]	#��'����V"QLwL=�γ���f��]������P��	�D���� $�q������0���UˠF�~N����6V�Eg�ɻ�O�l���g���[��d)��I�!�I��pۦQ3(��y�++%܄�5lyB��n4�T���ŻHq�3;�z�f��Jd�S���G�*$1C�n�Ë�B�{Ϋz�en�Z# �
���ҩ�%"�E�N�E�0̱��
5N�^����&�����
�<�Ă4���TqE{�l�F�&�~`�!
�!8P��63�C�5E����'Pܟߋ�\e<���e��+�S�dc[( �I��M-+��~�u�
����rq0�rp���	�<�U�����d7�#���ҹިy瘪�F1��I��I��qQɗ�Dʠ�b�b1�F���s>S��\��Z: ����K&_�n�7G��ֿ�p�����Gy�,24�\��D�X/f�a.I��
Z+��<\����@٘���A�r�z8nڝ�]A��d�W�P���0��]T����ʱ(�jc-SOjg�ƪ��I���r?lYA+����]�����}���MD���(p&��3��s"䍴�\��_a�އ�pk�~�Qs�Mz��&���6�J%s��鲡C7�^@Xә�i/�.��L�q�4��n�ؑN�v���;��@+9Ѱ��D������Z>�w��W��Y�~$�c����ZM���v�׭�]�Y=j���;��/�S!Y��_�u��RG�b?��u[gXZ2`к����)��H�Z���'�G�0�-����*���,ΐ�3J:�������něGA�>�+��yM�Eb��S��#��C�̹_n��7�ĤYĬ�`�R�\B�Ӊ�A�:�T�:EY�du�o��L��t�жtN���&y���M��b��	ϓIX�slM�������.�7���'��ʾw_�p��q_�%�֫�İ#Z�a�x���!q�B#1Hv�"U�"�w'b��O�	�!<$�F�d=;�0�s��F�O�y_����6�Ô==]�ښ��a7G8q/��~3��hl�H�ϙz�l7c���Z�1b�BH5(�Mμ$�#�.�aݜ/�Jg*<X���6��MPM���!��k7�m���{)}<�ʲZ&Ѯ'Xl���ۿj��������Y�_nI�B����.�e�I���1Bh9�+g��ki[������o�D%�Zv]�KO��L��]�ezB���E�Ң�,�����+�?�3�����(�2#d��2{�6卸�|}��\d�!�X�9��Ϥp��0ѐ��vR\<�\����p���B�<�e�}>|�e�+[έ���O�}���^�hL�8]�;�m�X�=e)���B���!��DfZ��C��^ڟ�����1��K28���LUL�4T�|,%��M��R�C�"����/;���{��pv�ڂ��#p�
o����b>�*�>��{V��ԃɒ�`�b�Cئ���.�t�0^�o���&ր5Q2�\���!CF҄�1�K�\�L�r�I%��w9�����+���C�6�x�A�-�����>�R���9n#�q%�Y}1�H�E�kѓ߾���ܦ��ۑ^��>'����O~��l���n慍���н8��4L�o���Q��z�����w/@,�A�XPD����F��6m��-�0^q�V�J�H��k��[�Y\��5�3�K�I��"�[����(r,�c���}bm�(��lP%#�~��J�Z*D���kF���1M�Ǎ�H=�fh��9���C����CJ1�ǿ��82MiGl�5�`���+k���|���a���I3��zGoG�[V:��SCʌ"	���8�2D���.��K#���<v��"y.R���&�0�ti>��>�t��߸ )���`�G��9+?�,���� &��������"�F�'Zz��==�/on�6hS0o�	7;�b3^du8c�d���{M���O�Q�-�`X~�~�4d�,RCI����R)������mV+����k����7�ǇGb�ǡ�v1lc��E���ki����*���L��e#���P�o�En�^�4�j玧݄�y;�N�C@�>^s���\�]	N�ߺ����x\���$B����=ۀ��m�����&I�{yf��БZ�X'0jr]�$�]ͪ��B��ҡ��?�����g�0V[��7�%_���ۺnJyیH��y-S�k�֭��� �-Q"@�l;�I'{y�������p�&5�����;.�hp9D6���}g4��n�[�=d��hA�*��ó�G	���� �@�Y�A�A������� ��\ʚ����n�ٲ�q{�r�6$&��+/�O\(y$HD�ehY}������"~��ݪ�Gz�'�oq�U�Y�"�S�ã׭:�h"V����[G�k5lF*�0�5YC��f��f�ϗ֟28��9��{���pPՄbu��`�֧�[������t(']'�ì�����;8���g��ܰxb�O�O�AV��f>2��u��0�}a�̝�ɂ�;���ۥ��,����dZR!�6w�����,_�ABY�S�4�8C��c7�o�f�(u�&1�]�K:����l���y$�5����Ǭ:<�i�.�gi&�C��W��E20�b�!�#{'�e�ݔ=��T��~��i>3��xh�W�����D����>�e	��k�.�k�v�K�S���t��y�^lO�s��r
��n�<����Ql4H���vB�q�����<`�o�9]��T�z��ԮK�	9f�e���]���ċ�5@L�|f�7'��Գ��$'�W�h��PL�������5�pMrK���ՍѸ]�u�.��#X���eI�PM�Ƴf�Ç� ��#�
L����7b�$sT������7��Y\3�K���S����?&|ɥ�.تo�1�$�t��;o!z�FuӸ��I��D�wƬ��T|wX*��Ԃ=�o�v[˸�x���@>��VĤ�R#��׆��
{�%��>P3�Vp\à�EK�_����e6��\+_=v��D���.Ґh����c�{h�u��Im��R�x��99c��]�v��	&b��Y�dE#8fZ��H<;�Y�=/�n�(�qa�!`�x�H0ڞ�D��/t�L����z�%AÉ ����Aq�4���f]0E�լ�vf�x��^,˞�Z� ��`�98������s�¦�^	P�\k���}a����㔳_��}�N���r8G�߃�:c�&�y�a��~X/�S�H�����^�����a{���{̪0�hC�qE��D2|���[(���>�r�ʏ�PY�=�� �ORE��C��f���s��\*�4�<Tz�S�9�Z[�^��}��lɇZ���!��Z�5O!=�@����l(��TWN�&B��z9�.0�x�g��W�޻� �Ye�Ћ���P��{�
�c��������l���	TT�X��9IYx��扥&<	Nn���b';X�������Q���¦���I��y��&� (���^Q0�7d��s�i�rЃ��D��ie=nh�ki��_��f���K�ɋS<2~�g�4�k-�?;��{2O��
�"�Gr��GQ^�ߐ������u������O+v��-k�廊�#���~�t��5��M�\��M*C���F�ݒstP"gwD�?I�3�98�]���a}=48
��	R��W�L2V���\5�;��E�����yx��G�3���d�߶6ڛGA�Q�A�f�*�	����ĭߗ$�P�L�L~��?��"��!�K�ca�L�[!�iw"P�o��m>�P�nW�E��&�.��2^���5��VG�����tG~������܍��V<`@�ӛ�����c�p0+
��6}#�O���}|I�N={[�G���>Jh�U����(�!^�
/W�����D2�RdjҺvi��91�LS�װ��:�����^����x|܎�ʏ�e��Kv"��w����49	E���Dc k%g�WБ�������G��`8���Y1+��D��8+ppw,iL;�����yS:��+W]$,s��
SJ�*��\
�3�y�R�gV��yn��������n�K�2�7��9`
����vo�痟���45�-�{��o*s!��RrOH�4߄{],��\�S�;��zϺW�'�t����FƤI��Eg�О��q뷏��0ϻ�83YD'Z���5tnvS�^�P��5Nظ���$���&��^��t��U��AV����C��UlvR����x�4؋�%���b�S��ϑ��O@_�u�]vẙ!S�r=6M��^_��a�����{i���W���:�0�v���N�lF���$���"�����a#��0aT���tbL=)���	�֏�DYtYM�?'9����;��k}�7�d�Z�~ΕU���}R��Sҹ@\�Q�g�E"z0�;��T�x1(�DȒmp�t��xH��f2�`w���3��>����"!�1��R/���R[g����K}�]g�y�A��*��Sƛ�ǈ�a���M�؛� ��j�����W�Pugd�]�������ӹy�[��M���
p��ᜫ�''$酙���.�-m�fj¨��B4V¿����_C� y�M_p�C��D�\�@�Q���<Y�En�PL��W1c�ŭ[w��ӽ[00,?�������#x�;��f�e�6�c�~.m��=�"
�mR�����L^�����z@��y����O�Ĝ�GU��t��ʨ!H�:�����C�N��,�=f������nD��8��^�Xn/U��h��U���䣞L#�7�n^�����w��O�ӕ\�z8K!(�w�[�qC����Y\�@������r.�}fQmH��ql^���{��L6v�u���ɨ�%_J���$��4���h⨷�,�@b�u �y5�s�Ě��4D��hY�4�X����xq�֟��r?�2e��KG�Z4�������4�V2�,U!(e�\h����a�����U����$A;�'�pLw���_�-9�t����&T��P�\rD��ʟXME���z+1Mcﳔ(�{�"fZ^�sؾt�p&��c��<��RR�������-�3.x�Gҗ}?����I%+�9N�h��=��ʓ~��n�L#Jx�G.���Yӛ>����&��s�A� $�	��$`�U��Y�M�4�XX�hr\�&F���ᔋ}G��6A��q9]:�F�5N����	����h/?����)�r9��o��o9,;��5I�[5����Q²�r�@��Dxn7z��r�_r�Z٨]��*ٸ���:n �}b���Kq�O7�g4>���W����^��N'w�t�����0ά3f��[�9F7�e�m�̌<��S���;�����^'`�^S�7(�&�)����b�H�9��qP�7Aڐ��q+d^6�"�/)��}�n�bb�i����ߚL	�l�.ߝ|:0S�
������Yt��$�l╳����y5�*F�u|����9��ե�z��s��ɀ��TH��hCc<���u���ؖ�K*�O=�6&~� ����ɩj��2[,�� �[Ggq.\|-(���E�,�8�5����}����\�i�
�<��͢Q�C���؁�G҈A�կ�7ƘּE{��3�hF��`�hA�?:2�A���NkY�{
Y����a��A��V7���k�w@L:����l�K,�6dY�������I�
�[E��;�Ύ�A�2u~�+/ QkY%H�֒��2��h�z{&���{��m��rNm�]#���'|�Z���sR��������a_:�����rh@��U��Q����djB[vg �T�9i���K���R�Y��Uۙ���`��)��<����0��%e�u�/�I���%����EF"�pIྩ��fa(f!e����a�$p�3�\�uq[��{����)C�J@�K;��m8�EZ��Do�/�I8��v��]����/���M� .H<�ϜWf`�^�0���A\�PwM�
D����!g����&To�! ;�S�N֤ㅂ���7�Q{W,��l{&Y@�y5uB��1<��E<;��"���7{W빎<�X���/��7��g�����˲�� �{��� �YMԛS�;n�ITѐd��X��^�s�]��.�(J�l]�r`�>1N]����MN�����h��Iwm��|��w6�h�ʉ����b-;��JEh�N�%�oˌ(A{�G���z�Z.01��<�"x�B� P*f\c�N�1j��������C�/X��5�0Ӵ9�<>�*�M�m�۔`��ҼK���2�T����VA�;�c �ŧ��O�D����srӄ����� �3s���~���a+�M��a�%̥x�g�8�+������p�/��j�@�NV�jٰ��V�/5�EWQ��ōU�&f�5۷7%4��gdӞ�Ҋ� y�m�-äw�Y� �7�}�+����&�
��qOۦQ����
A�xL�F�F�����������a���`� ��w�r����h����1&��.�
B�D�*�� Օ�����r:�����F&� _&B�}�ݖ ��;�#]n�d�5���~	��ƶ0�t�~�����U�VV�ݱ*>N7��l��HD���y�9�L�Ek�mF����mX�g��kj4!q��$�������T��b|	B��L���u�C�i���^��!��)]��3p��jCX^�:�s��a��k�y��H4堡x���5�?����q���x�΂��y��f'$aN�����]�Е`\W��t��j�ٴ@��>��n7�ڪd�ëO��.!M�����-��a�n� �:�2��/�W�g�X�����ű ;�寉J�>�Lb���UU�ߚ{\x�p���7j7J�4��8�^����p�ǝ� q����X$_�)t�;�=i㜙+�	��q�#�A^\DF�{)&�1�O�Fx�w��l��|�N����0Eb�vd��St�"�t���ϓ��1�/-�[�V�'}f�(��OƁ��S��?���4���!���Xwe��_��m�->0P��j�xd@��-;t�������J&��V\M����ٰ�+:���z9C��RVA�'�����B���D[8C!X^�!K��W"���J?e֥$�LF�`Q�X�X�����~Wn�*Il6e�s�ۋ�����t���Vā=�����O36�1�����8�<�����d
����/�\�@�\�">�IT�����1�Ž�]WK��v�I��k�h�U���β�!Xx$x��T�@5�綩�ӕ]MgZ�GxNVy8�Pt�&�������"Ս�