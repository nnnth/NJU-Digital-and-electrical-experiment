��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�q���4]oHe��zL!���V�I3����?3�k�q��>`����G�"�P��-�V���z]<�zצ(�n���tOH�k��q��h�����J��j��a��N#d#^Y����R�Ѧ�Wԙ?i���~*�s�Y�eqr&')!Ȭ:[�6^�Z$���~gS,3օ��jNy#p�;$������(	�(	�<�^7�@��Ľ-ǐ"L��?�>�i�1toBӝ��gEH��g\W�_h�o-��������>6���$J-*��2~[2��ٓsD6�_Br�VN�I� �Z����-��j[H
�t8{hؑ�=�6#���R�jtK�l�8fͯv�
����+��r�^�P6���۽C2��R�Nhj{a�cq�t���;��H�y��\X�m�j��Xw��%�I�#M*���פ}XU /���2L��|a(�zP$A��� ey���ϸ����L��Ş5�X�F����)��R���=�+b1%r��B$�a�ϓ����w3�eJ���R�a�Ь4!=uSX�C�o�m��Y���;Ćc���1�F,�+�WSj}��P_ط�|�@fY%>�vd+����w�>9� �$��LX��F��uvɥ]�$���a�r��j/�q��$�2���R�K��1*�V�L,�z�m��IRr�_���!6����ȕ,o}��%�5��gc W��S��5��iAz���`�F1 Q�K�\k��}�sa�2�|#�K~�ռ�j���p��!`[%�P����u���:��S"k��<�Ц+z"_׶	2�����=ǉD������P`�ȥ�t8��MZ�U��*:,���!���vg��J��ܜ��b^�J[�qf�k���a:g��st�����	���0��>�*-����+��e�Ɯ|TW���	���b �����	nWK�nh@� ���Dܪ��*-`u4sߛ��3f�"(;�9#��f���>��j-!�bvc%ʭ��Mt���,�y�XNH���ita%+Qx0W7i����X��?!����򴻋�Ԯ�@��.?D� A���Ŀl��-��ѧ&�Q%�g}��C&d�u�	2�h&BG~7*g��o��ש �W��,�Hv�0Q`�!���%�?_!~��$@����?.\����]�N[ptE]a�A.�e�*��7r���������꬜�o���<}��͚���[}U���ɯ�)����3�~����Q�u)����Pu�v����L�(�����͑��*B�7>KӴZ�w�C��;��ux���wT���$Qh�d����'��Fw$Q����#�ʚz��6�����h�w(�i1����	�S���´ZZ�m�W|>d��M&A��֛<�"��9��P׾�� �:P|�H/
#���"�����R��W¯�^p��b�]	D�f�k�^/n�4��Xp!��)j��!&�T�7��Z���N&ݤ"ht�q������ ��[4!c��b����mQ�MQ�b��^�M��y���/��/���Z�l����C��u\�2��%nt,�*���&