��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��3�q��Xà�C��tt��R�d��O��I�P4�X��xJE%��y�m��W��+��̼�`����k�@цSSa�,�sw�O���8(�@�H�RV!�V���;��?�"谎������ysP�>����|I�Y%fMc~�A��a�ݪk%ݺ ��' �s]��E��A�e���F�5������pYy���R׈�d��vHv(p�l�YO���H@�$���M����U�ؓ����AM�����~�t^Z񧓮P�43E��]+~��{pC���C��Kg��H���}�t������Θ�F����WD�:����i�);��iKC>����jC5�^��ؔ��n�&���{)�r�P�t�-�Z)M����Ua�sa��ϯ+��� ��O�WmC�G�f�@��aQ�BI�F9�d�ȡ�ܽF���]kQW���hzڞù4k��}�H��ݹ�0���P�[S���?M.6�-q��F>A���E���/GQ;F<Fr��iH���ZB�/�����>$�r~;�㲉���`|{Q�R����n����Z�X7	+,j[�	��?�k��VA��Z���I;�2��s��;X�v�v�Fz���6�~��lڇe1�j~7�;�B����C�d�mC��/$0$�� �/$��23�d�["�#3(�Ր�g�VEz'�|V$��M�g�љ�E-�=��@���e��v�-C�� C�~�$�,A�\��v�0�eb��Z�Be���,�0y��F�Pd��]D�!�}2��4�L�8-��5�O�=ʹ
��ބ>�&���P~ţw��%
i�R=�y�$'=w��C�7v>yj=	�m��pՅCd} 뇈z(�C!qIj�v�q��jg�&s�Ŝ�ٜIt]���E���5�6BfֆH��}��bb�V^hK�B�1����i$Kfu)���Z���Bb���9�U�M�-��4�YE�St���A�n���0E7�PQ�J�¸I�3p_��FU=�:OH��*�[���W��!a���Ɗ7�)�J#��]�0�T�I`�%%���M0#�"*:� c� � �3��Q�@�E�.9^��h�e,u��/4?�? @@�!!�S��P_9vϕ["m*m�I���\��j�/+m�$�Û#���������,���1�>fu��׬Uκ6H���-3���Bk��{�D�n\#>�9��c�jO��{�F<)d����8R�����'��1�C3|���g��3L��~�e�k�Ʊ5�%�̆yylQ�*96�z1Y�/�L4�S{�m�˿�s�O�j]0(�M�1(���X��\�����x��UwO�m�W5N��D=�h�#�4a�ܸg5"�è*�q�N�{����.Ф���P3����"�3�A�d��d�����=�S��2���u�/�<�WA��>q�����%��X媻H[h"+��$h�\�A2ʛSw]:A5S�d��4?�L6~;�D9���B��Gܻ��}Ȯ��`�:�J�4`��u�'�,��BT��ubU�Ɏ>��@Il���N��,���|$Ζ�8��L� *��E�-����֑��R��Ͻv���C�k@O���,sKJ㇮�:�C�-
_��i�&��F �Z��,l���)iO����l�k!L���,�,�hd;M̄�Ah��Q�
���@������� J(�A}�l�1e�vD+=#(-��
��^��LfNe:�0J[.Y���w�g�?����C8�h<��pܵ�K�G]���N�	-$���#ˈ7��\+ß��r� İ�,�@y�ô�������Ҁ��Xa���3r>�,��ű�ܗ	n�*�_�gX �i���t�	��E�� �1}�*�C{�B�
�AzL�,dnu��� ���,����3�=f��Z7�K�_��&6=�T%�W.P�����4��B�|=�N2��Z�4]�[g���	v�����a���Ļ��QǬa
�BQ>?�@�s;'p&��:�*�H/}��r�2g��Sy)�7���@9M'<����6�fT�"��aa�=~�jn۬^�p!5���o~�ӎ���n�[l��
�k�n��a���h����]b���;����U}40i�Iw�����t�Vq�>P�/1p�mOA/�K�P��n��!-n����_׺l�G(�r���ᶣ������%a�A@ZMܿ[)3n�?4	�%�)!�1���	���v�O�
��	$b���@ᰵs6O_p�3���'5,�訵����:���v���ߐ��.�<y0���b�MĊUq��w�&k��p���H0�wzͭk�@���h��zR�2*�BX���^��֓��F;+����	���6	UO=!3�����ݰ�0��B�Ta����J�G��z�c��7�1��*C��7z�c���$~�
�:���L���ҷ�0	��w�˚��t����qY�#���$En��	��8�Nl�!
���)Cn~�8Vڰ�����S�NoE�-�vI�U3��w/f8E�wQ	"]Txr7ί�������k�����m��?��(2��]�f��[<n$p��)�7.��o#@C?��cⓘbD]�^i;��S�H����/7V�fQ#���=�����f�@7-�+��i��U��,]#�
�p`_���5c�@/�8'���ua ˈ1�Gq׊<y9N�7��wc*��wx�P#߾�[��c�V���VL��~�+N �Hb�0?̜y1��$���B���w�a�I`.
�Y����"�L�����`r�:$��@��rSV�u-';j�d�e"����Fݪ\4������0�x���ʿ���ͮm����&�\�F�s��@�A{��������Z�֋ ��{Ս��JO׹<s��B/�3~��N���ǡp�;-%�/vUT��_{x={^ ���"ͣ麚'��y�5�9H�<���T��S�f}*4����7?
%�O
�����.��/5�%�p_��X�g�Y{����I>���'���I��1~�:1��
i��#�y��e�q�q�[�V��O%B3�.P�d=��[l�9�B ��n��u��G=�_z��Z��8�'���OfYR�>�=� ��L�Y����S���x�[�	ˣ5>�UP?�7�6k��c�-�,� ��͝%ĉt?nWi����QWH�Fط'<�Ŗ
.�_L���]��#�ۑ�}y+2�?O�����&R�*@C��1r���)Ь�-�mJaf�∽{�=b�%���
����{�l�w�h���̋;���w<��GE�3���F����
�Ȋ�� ��%�K�i�]?�`>�
o
�7��>W6�M�n� @�1�3S�!bx��6����vd<Ց�d	�@�P
&�g+!HR���cb؅��x�'���G^
�'��y2�x��wx"cۇ���v׋Y����ǀ��_E�$�?͟Ud���2�.)�Q԰���ėA��y�AXhC'/3�M�Fw�\3�?t�Z���ԯ�9"�Dҭ^?Xi��u��"��#��mg� Q�W�(��6{Ef��q�b��x���]�L�]�)�'����IK��u�>z�ޚ�mF삈�����:Էt��,�]�'��Nb8�E
q{ѐlf�!b_���ݹ��Þ#��`t° �w��Y�XQhGY��a�7a�XY��m�4�Ѡ��Ov-����_�������%����-��YDp�T(f9��'�=ؖ����b��N�?kˀ�s6Y�{��a ���]�v۩B~��d��_~�@6D��"uFV~����,�KdJ��� 
��#�<`�E]��zZ�Q�[�w�er@XB�j8S-�}��H#�2���F����h�p��OO>��8it�)�@��	5�%+T���!��C{+,*�1���joz�p>��V�<���K�ZDO1�$��&P�J��-�KʙH��> ���]H�K:.�<�* �4�����BnbJ����G��֮���&��}$�M�M�vIsk���Jb��mVeZgo�_������~2��ҕ�t����%�2oO�%���A�)�'6ף�X��+B췹/�!^)�©vk�'p��, �6c��r�Ü-�&�����^3���8��Ժ[�]+� i�m	���5zk2�QZ ���D�o`Y�é�;��=�}�y� �,f��Ƚ*M��:�'� P+"��yt0��p<�� �K�o���7�eY�2<7��xK8e�#�|�ЛuN��A=T٩,H�Jn�y�}[ɜ^+�u�>w���yO���-��۬�؏n-p^�s` -{d<�^��N31ɻ��z�`om;��4W�w�F�[1�Q�l7;��Zq2v]֥�uz�Cp]�aS�����lj��Ĕ!<Iξ�A�&���i"����ϐ� ٧..'��w3�;�g���Gk8���(B���޵KJ>X�#�3�Ċ��2��)�ɶQQ"���e����u)30��v�/��H�6t(����g ���ǽ�6;�����4&�{�yq`���ސ�X�8W�)�!^��gp�t
���b���7N#��́u�t
��'��C(܇�I:�l�6���ɱ[�WJ��'��H�2�6��a�؄	����$ظ��`&-�x���B��Q�5��ui�4����y�,iZ�xi���9��6f8l�4#�g�i���
���
X ��0���Ω-�$�f����������`�,�^��8�����)���_����J���c�����>���Z]��e�y�E�T�袼 0�V��� v�̌ʅ��_m%BSZ� �wȊ/�3�	ts�j����b� lb�\�2h���On]8�$�͂)���c�&��)$~,�#\��;�:4�q2�y�a�lU��Uκz�c)��R@�^;�����;�r��-E➟�N�D��:�'��?��)���.�'V�ӥA\Ȝ	�	��^U	T�H���|��x�w�ă �XFQ'���-��.�d��\��B��Đ9�y�l[1�}�V�Ǧ/j�����<�C1���p�\�	0�e:���^mH�M��'_NA1%��
a��e�޼2���QbM	�����k.',��c�)�ݿ�8�.�2{�<G��o�SV�F,����`*�pH�A-4x��T� &K޵��ԕ��I��^!��e~?��q'�E-���d�I�����u0��4�{�ۤ�o��؂�>��Ê�3H	����Y����L���7Dh�Bϔo��2����1�<�c�����-�0�jHx`�BDė�	�#kooJ�rٮ0�����s��u�O�DqF1����g�UL�����aCp=���:���a}�/��]#��|Ww�t�Ϧ��URf�u�Ġ��i��<j�}k��� ,�)�|�΃�,�>�F0I����� l!|jtv�y;�s��<��zS�T���)m�m'�#�7;�!��^ C'>x��<���r&�d�ڗ�O�� =������Q�RH>9����ʎ �=o�K�����1���"{�� aŚ���@�a6�{� i
��a��Aڎ�oU�WѢg�A8��Û)��;W�hyB���M &2q$pY�O��r~�lD8g#��nT&Z�����u$.�ØUP��ֲLiiF�p� �5��O�X�Pޞ����)�ĥB�c����	d�o��}Tr:sQ��-�+IM�9%�K��b4�����R>J�2lG�o.�럾;�8���*���� �z�����n��ԩ�Xy�W�Ř�4\u�("s4�{p��G%3��SE���_W+�k3+���˥�|؜u�/�|�i]�$)�v�����ݱ�F�#q���ݮ��p�S:X�c�㣟���T����!čC�z�F��~��%t�8<�jƶ�}���q7Z���\)��Q]��6��� ��ڤT?��F�˩��ڍ��=���rc��=�+D����X\w�Ƀ��w+�;
�x���(Xc>5R��)��\WW���o�������P�1���e��E8�͡�����a��[4�.�;��+�����P���i�h@ʀ���_O�1�X���6����C�r����A��ℹ��-Pr��A��?�@6A?�ͧ������|�T��L�S��#Ϋ:�����p"Uo�q,�69��nb��f���גBMc�.*�ov����r1����^��$�u0fR��Z���*�N(�Sjd�� rx�M�O.dce��T#u�v^V�Dm[�z��s+�<Sb���{]֙�%&�T�vH��eߑ�M���0RGh�|Ŭd�+%l�a�G�B��3�2���?`!��M�{�NA��%7�#���1�j-�m�R���aIZ�,RXb � ��\�hl�SwP�>o�<�wT���:��/ �a�Z�
�N���w8~���
�ԟ+�k���MڴsZ-��#5޹R�L�(�g�1^{��,X�g��<h�΅c9��ڱ�@���
�Z�>I������Sľ�� >&X'	��"�=K`m�R�!^k?�q����`[�����1�.��v��j��~Ҥ���7�]o��:�ǡ:,3a��'w�y�[���P���(%jJhӄ>tSc��$!��ᦣ��0%~�(k��>��+@�s"�A ��?16m� !�>H���O��%!� ��}R��k�"���}���&*�h�g���?�۫܅
�/�7�n��H���w�����S���B�Ƴ J�e{[�E�)o��q�<�\�Zka�+�A4w=�,�PGO�<�����%�'�����d�ڼ�oTe��Zx�d?�&�hN���j%��٫)�@3m����U��ӎ�n �=���諥+�(H�r1�#/fZ�2fa5��=���<VO�y���&PR�P���qrRd�'��a*5N.%�T�:��C���61xb�Aޛ���֕|I��=�>��|�2Q�"�*�po�2��q�CMA��!����Jڴ���:�%?� 	�0�>s���$7�����/�/�>�l0�wG�cP�oxH��s��:��*����K��u�e�w�>�;�FtGD[)�N$Faށ�!�S�j�����WѼwbGGx��|�7��QJ!��Ϡ�����X�Q�$'B��<dy�C�?!K�f�ﴀ��c��ϲ�UT�Y�/h�GIаI_:��zDב��`�bu��;_r�`p"�Ы��ί��C��_47�^�ܺ�&<����	x���uyٙ�+UD�\1Ǘ>���+���k��t�"�BlW�iW�;��t���
�ۄ�q��*&�d�8��1�75�(�����32TA��Pt�r �iFAo71�x����a,�y]��n[xԥ���谥m�X����^S��b�m+�����G]A�)"�B2�\��Hy��r/i���Y�<	�:Q0���u���;&+(AFsU�zWœ)FItX�ޢ�b^�Z(v���pW�	��3bT��8lg�tE��B�U��p�������IR7�+ϖ4��+P:PQ���	�x&+�d���%��UI5�v��ך�cA�)���u��0��Ȣ"e_O0٨��4�e7�J�m��[���X^��%��GUw#��α�M���۩6V�� �ڃ��{���D3	z���:��
T:�Cϰ�8�Bh�si��>6"G���N��^Z2y%mb�<g4��eD�A��A���Ȫ����r� �I�R�L1rQ��A�COe�Hj�簣���"��p���2SNnV��d���t�;H���*vk]w����x�.�!cB��7ޕa3Ɉ.�D���e���E]�`���N��3X��k���膳���h�8,�1�f5{EA�\7�����"#���1�m��wT)�~�<oH��;�T�
������Y~~._�*�tF^#CC��rЬ��}L���TUP�E�r�4M���_>�srub|/g��)���*���߉Tb	�~��z�Mޥҋ��l�d'�Д\QN��O�=GV�{O�@���>Zkܫ
RQ��*�s�!ͽ���#�e�� Y9��}@��E-�e�f,��Ǵz�����[�|�q�v0��1uO������_���y�&N��)W�������F��\�o��Sx��7�]Y�Wҿ�����NU���&�z��̱��U\�\`�7�q���r9;��X��u���'�k{M	���E����OT��gz��u��ux��z����@�+�P�>2L����	/g���w����l��0T�]�fL;�#a�O�����o�"Ÿ:����Ql�ċKc����g���J�s1�a�j��lm�9Wh扲~����
o��
7��r,�3g����lh�=q�����g?C}]T�p>U&�a~�M�/<����4���[#^pa��{���9��h"<�)����J�ʗǮ������u:/��;k�no�h���֞9\�r_GHJB0��bO��iM;���E����7����ݟ��
U����NC�"�������̏Z>���;Ͽm�
�E�?jQ��P�:�K5�[�� �1�,���m]�C����%�(�{��q��y�"�����l�B4s)�S�lЭ:�)iv�qiOpd���gR���F�@�MO������ٛ�-Л��p�֋{�۞t7���P���𲔔��ND�12S���Ȣ]G�K�'̶�r��Ҟ�3�8��UK���'|E���
I�L$jFu����t�YP�W��v/5�#��Po�v�M�	5Q���:3ָ�0X��$w��e*� ���D
G�}������_���]p�s� �i��~����c����.,�I	���}cŻ|-NOT�Җ"@PM��k�n|�R0��0�v�]����;j�etk��/�|G\U�\����L��������HHt� �o�(�j6����'8B���4�2X3�vZ̼HI�ow΋ډ�'�G�t�L�@��?�\$v��i�,5�fr�I�Nt|��Xu,u�Q��X��&>�֏�$�G8��bs�E��w����uA����3�5�[Es������Q
���
\!$�S�Xo^:�]�K�:0�d%#n@�^�F���y�.�9��^*/Ε��p���~�8����4�°�~*�a���+h1Lc�as��B���|�;�b�ޤT**��*�-��W�17I�Ϳ���Ǫ���M�K|j?˱m.\�zE]���x�9�6�9Ykaa��ܲ��n]��]z
3D�D�Z�T���D�&�нQ�JJ�g�����y<]���f���'�����` a��VB�Mf���lu�����7@m|\�|�o�w����D�؄aE��'�k���K+��\	���%�t3�M	nb�������ڸ<��L��#��Ͼ]j�Y�վ�Lj$LV��7�h�iԱ���-�����FF3֛��я"8/�=)W��6{���C�����M���-��V��y�5������$������+�c|S6AҏF��ym���j�Y�d����b��y�;�l`�#,���bYm�U j�;6���s,IfŨ3o5�ϣ9Uv^>Eh��c=+�tAs�)�}���-�<��� .���""A]�%�$��7aDj�����#��%`8(Uײ7X:1��p6��+Y+Ll�eū��I�~����R��x~<~Cը\�q�����&:Ղ|L�`ı�+�1�O��R��9(u4��+u��%���z}熤4��LU���I�`W|���L�w��	�G�<@[G.;ޤV��a0y/]���h-�d)�\����2��8��:�5,܂���9 qjW�/e�7��%��E�����H���0����z��'�b+�EGj�}*�kKGZ9��9�����b0��N*�	�}�=��1���U�6�蹼bd�$ؗ�h�&�PH#�:f�)��)��+�)�<T�ܳ�v�Ll?�u��i�m��kʱj?6?}h)$������nm�\blrrE�+�!K��B��z~g�V�ߨ�}ҩ��~<󔌯�)d���&9�j��|m�dZ+k���E���j?��^�7���L�.U&eYL���h>)�"��Td��]�8���=C{�1a��6q�S\�M6����5�}��2��cf���4�(���2? ��7a$����c|�̰�&$����dg3�cr�}���$�UE+�^��g��S����X0{�C�Y� �Ԩ
~�ZN��{�Z���p@���m|ɐ�҆�㡰����z�X9�*�"z��x�}�4��O�+�i��@*�[}^��Z�ˬWJ����/�8h0���@Y�
�.���ҋ�X�j�g�O0ׂ}b�^U���nT���j�P$%�3�$�s�����dV6��%KX'����K�"���r������0�Q��.E4�d;�yI/�jO^�0L�Z��Z��9�)_ީދá����}n�=����:䙏��=�js�a�2�Ė���r9nvH�Y�T6W�1t����6.$H ���|C��[I�9Sq��d�����*/0^�'�4��"I�X$��?9��#'T�L���S΄?3K�ҵ'
]B�l�e9B.�&��*Й���E�
L�fXi�R�,���9㜕�d�wXYԺL@���,i�#�j�b4�&j3_����p!��J=׼p�<W��\�#ۙ!�
�y�A��|T�&Ն�>8�����Ռ
a7E��4f (�����DV��am�L�(F��Z_���
��BY�ܣb�:cdTYܒ}	�"��#�{ ���nE0i��Hm��~HEڋ�Z����\�BF��?w�W�*S��i��6�>�E)x��v^��F6�!��2w�8�lJc�/]'	�vn}�� ��g�,���tm"�w�����	�FcQ
�`����c Ѻ�iQ�hi�