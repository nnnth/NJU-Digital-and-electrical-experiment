��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��RKj���B�}Φ#�Q�%���L+��*|A`Bow�g)۰a��Ԇ�Tv��k#�fU���yx#2<s�����_I3"�ꕳE�5����jVcE�����"*�k���6�&]�ƺI,���!�s��S*��y�v)���lA�$���/�����V3�'|^1]�t��4��6�y�я�jx����؄:�&�C��2h �C�Š��{�)4��Yz�]�u�eW�թڲ��QM�YSÉK��a�%�.�q�������B�#�u�p��仏�� �I�.�3g�g�$���Έ�?-vx�T89�Bp�������/JCNJ�xf�Op?�9��C��:�]4;�����~��+��9#(���$�>V�oH���60FuM".���)x\�5F��ͷǛ��=�k�S��?���\Wը=7C~�s�X��k��R�b:�/���][35wLmO䧭�Pj�K�Ⱥ��t@U �Ō?['��z�	����BS�4��d�P�+�CW�(T��{]hԖ�����%�3������j!?�8��ى�͑zf܁�E��N�0_J��f�_��4��"��~�jg��:x����LL@���1ȓ,��Y���S����$pԆ�&��9�Op����%k+��JgY�u`��1�2@!��5C0j�$��&�T��l��wm9�R�G#n�����Ol��vݜ�	c�7\g8��Ad�S[J�x�hO[ D�"��h�B���d�sb6
�=�K�~���5Lv,x�T<5��d�no�R�`ϔ/r��g��1`�����)x�uI&,���ؽ�A�ҝ�B/�TF���w�;!���*��z5)a��Q&H"om�]�1gSi���\a���6��b�`�ɉ:�>{��4!1S�ܻ��I�V�Еj��d��E.�`��P�����	��Ͷc=���YY;;�d�]�dw���q�����s�hFk}��q�کJ���&�N��@�&ܿ�ܰ;�R�>.n����2�u�d��	"�Z�������l|zE�{���8>GBrnJ���1PJ�^Ғ'L7m�,�j��G+����^fv��,xNQ��":������0#�M\җG/�lT�'|�e�q�$�cGA��b�Z	��	�Nq88L
ٻ�
�V��T����חB�fQ�3 �
��Cv�[� ]D��3�\LV"Q\����z��:��Q] ĕ�/��M��rf�:q��م��(�8�5ר��κY��BO��O�4ޥl�w)(��_�a`��H��f����p���"u���n��p���6����׳�~�>N%��;���
v�����h��!�C�/��5�P�n�D��5,���0u���^>�u:�q�*=�r�7�/G�e	��y@�f��M��aݞ���X�O9W�	��	GD��$�fD�.H�j�9��HZ٢<[(S\%G�>ꆌ��rnʷ�U�[.�F�Q���|����?5�-E��R�����Z��`+]sB2x	�.�j�s?��������9}�?�M4�'7р��T�oUL�h���t�g�T�l��l��5��O?&��A�Z�X��쥕S��oS$����x߇��Z"r�>���Gc$g&���d6_��g�3��L?�a�����paPP3h������d�٤����*����(�i�
V'�	��t�Q��گB����ؿ���+�gH�G���F��$yv�]���=�[��)���!А���[F�{�csɋRE���&|z�kx�/;Z�%��6=\���6TX<��#f��C�I�ȍ�FMg�,+'z)��E��:R�z��o����J���8/��o'8"h����[�^��Rҿ� �[��`��-�ﭏӝ<_i^{�%HC2��T��&�I� ��aLF�J~��I������C�
R�Bq������2�pd1 �v�;�����/�ߥE��	0Sfx�Q�Ϟ����2�
��Y� u`��x>T�'�PJ�є�&�4�zBgW�0�P��>L���*�G�)��X"��N��]�7��YM��\v��!�MH�':��Y��J�r�y��.�6�E�F�)���C������!���~��Đi}��>�Y�W��M5�.t�
|t�����?g��D����G��p�L)-'�Z��q`�f��UK!�&�ć�f�� ����\��i����DMu� O�L�9���0�R�CT��m�����M�f����[��(wE>�"'� ��m�Hy.%��h6��q����F,{b��	L�J�]L�a�QA}��;�mT�q�h���D��RBb�U)��'"U����Ɇn�Ϡ�B:1��m;Eߢo6�j7[����GX��"��v�_��!ʃ�>�|tc���w�+DC���<,�������XR#����F���ޮ��S+c�Q�my�������t�v���Ϲ��s�$��8�]�|�����v0F��\~J�;�ݾ)��"#꫖�*G�˴�O�*�wP��n���ĴlQ84���LȾ��W���M4L����Wf���Q���_Y�ő�����-v�'^�{$a/��{�N��4]l���w��5~v��@�u��L�Ԅ�ä�!�`�q$ �	��dUH���ʉm�*3r���?D��g:X�epkI���cü V��;��>s�8�v��+ׯ$\۬��&�� ��_�c�,p'H���m��!��y
������;�{2�֜8R0�u�� .���M���CUp����_�\\�$0j���K^����y�fq�f���v%����E���4��Uu��Å �%�ی���H�(�ճL��oT]]�L(�{˯�+�{�
�݋]DL\�P S��s��jY��,bh��@���DzѪ(��.��A��~a�-~q]!�b�,0ɼ�"7�±i�D����YFBLSB�&�5؜�#Ԗ��- L"�M~Ǭex��U��� �CB֞"�<s�(c���A���>�!�[�T0���k�� H�)���������E��Z1i��5=�=K�ӳ���r(��oY\�r����k�,�S��9�����:/H�$�@U���`	.Q:57gO?��"��
�
|�P>�,�w8�F�!�;k�z|E�.����&�ݳ�@��)�~�ˌ��v�5a��t 	��,D@��9���E�xM���x�;}�rC�cL�q�Ovi���b,Ѣx��BWD�P�9�v_�$�<!t�pUSjÔ��ZdB<�y��.2RDP�a�0#B��\�Rq!2Z��NQ�HL�C�Ws����`eP��gي�f ƨ���,n���`�[y�o���?s��T����{������|O�5��|�(9�b6N~4T:��E�u�����QcS:���.:��;��bXSp8B��Ys+5�E!Op��[��¡+ɤ<xup �]G�4��+P?'�h��|�$�j�FB����4
��1P6-o�=��`4��AϏ�r+���@kƺ�[)�$ yLv�ֺ$�����UE5��%��� �ul_�ёB��jpd��Yj)0W�(rO��/y{���[0چ��Ŭƅj���@�=�2�����S=9���Y��H4�3S���LR"���&g��q!�ؙ��E��
�®\9jhD���F�ڭ��dF�5�bLPU�z#���*��w��� �����9��'�1ßJ �3�S�%��:�e/�Nb4ў9���JE���ض��2����R��+ߣͧ�B�ٜ�(st�`pk����⃵�V���	���"�ݰ�C 	��mZld(��P�m0���/m���(U^��wI�F'L�@�$3Z��d��[�����ֈc^T�XRds�	� �W�B7#�OhN��@�Y� ���K~[A�j�,�q�i�9����^Zc�\T��fJ8oL������l"��_�8B@nQ��Ŝup|�X�׺bN��o�!~�w��W����R"�5q��G��%��n]�ft��V6C��*����@�|�$�:C��T�6|<�|���u\{�Q�3 �XQ�����t�U��Php��ܣD�� �gj������HB?�N��AS�J�4>�;)�"�H
�5�����zjvK�c�+�	M���= �+\�0�܇���>,�_i�{]��D�\�Mꯠ�0�n�&H�|gEY�ҹ�[��clT��s&�E�M�����	�Z�P����4�ب 	;�O�-*rK�3U�F���i�%%��\�
���Glq�;ӡ��`8d���N"��u�`�v����Y<�[������g�f�*�����j��X���z�
h�O9�ĬB�;���/L����,�'_�h���?�)�U����d�,)S�+��cp�Z�/��u�4W1{G�<R�6�g�Czv�R|2tc��sɭ����nN�`_��(f$����}��|�`��I��mn�M����P�Z�ek�]-��<�E��O>*+A4�iAu�,'v��`�m\;�i9z)����u��F%L�E|�U[�������u�}�sDѕ�?��"�s��*�3����1��Q�{���%H���.9���!P��C�	�v���a<C��]�q3�SCԑ�T
2�����4�B'�������U&��OyU��n� 8�y�I���@�dv��}����l�-(<Z�z���著���ckٛ^��:D1���J"��$$�`|DsJ��x�-��͝s�]����J�V8A�}�Syx�H���~�g�L�+��B&�H��}4��I�rT\J�Z'���(� Mi�Z<	�Bv�C��1���N�ڌd��3l�����:9�4����=��k:�F��ys�Ԙd5�!��Fp�G�k���O�טq�-ܜc����G�&�����`Oݨ%�ѾتR����RK�,�)`pʽXb��zCc�6��\dN�)��w��fK�W�M �kT��v�|�����ƅ[�/Njà�Kw�O.�V��ݯ��{��!�<�!<��T�5�5
E�گ9G��Pu��C���7� Lm��+3��\1$�1��d���gi�۷HE�P�)���SB��T<���%��%���NY�ƥh7�ͦ�To��g\Q"R\6��5��P���Ɩ`i���-=��2��3\g�\q�Hz�͐⨒]�iN�q`:Jx�`Tm4�-�f/xB�9l�:xR_�Q�9����G>=�w-��C�����ŉ����"���pY�ψl'B�Av�ͩ-j�m�%���0Bv������b ��@gk,�� �(��&#��F��I���9�M����J���Lۍ��gķ�P�ӳ`��)�K���#�5)V�U6?$�!������]7N� ����.g�.�?>t��&H��b�O���K>�lzn������8ҺϬ�{�<p:��az}���ۤ�J�*>Y��*��e$��u������W�;�-���=U{�VN�IK弅�^��P��R�#�C$��		���l�#g� }ϟ�=>qawsO�7��b�'`��(J�
���A���4HPg��B��DZ1����C7��v"�N����+��7�)��c�¦���#��eS�6h�5O#��}��	�#LS� H�BLV���*~1S3�b�⥗j��r�F�,i�Įl�-@��s�/FQ���qq#�j
J7M�Մ�e��o�SZF�j���s~v\�J��XI�%&R��֖1�*�!���p4�N�?���P|¸�F{
���O�W�.n��"�@f�Z�h,+�$��m�j��fy�J�lP�q@���(
7*@o��ť��ǛG�6Z��$y*p%<�*��n�Ӣy���=���B-��^K�C��\�Y��1n���68a��c#�6M7�exn�BR��@�ɒ<!�As�3%� )A�����΍��oƯ�T+|+���Fwi���w=���Q�ż��������{_`�ܫ�1�;�W}���	d� t\��l�C��i\��<���H4o̓�Ѓ�C�8�B�C�T�.e΋qw��6�=��ca˗��r��.hv`���e��Qb����P�Ԍ�h��!�n��|��Q{s��5��Xr �q�jg5M���zI_�MD����}G��q�)���O��̬��B��'zMA��}��h���DUG�v����b���{��ذV�ll_�<�U	)f��%r�W|��8��(��e�]�������Ɓbh�����/Uj8{��P%������VS���鞶S�N1G�;�S|�$��+��M�~f��}��7w �f��I>��!��_pD�Q�1$�J1����_����|���5"��0�HA��a{��_�xS�����e��rҚ �^!�ڔ1oq��}���YH��7�!]/�f /r�Fl<U1���ATȟ����0B~:�so�:���r:���ͳ�:+H��6_m��ԧ~I��H~�&�i�ј��6����Fۤ�� p$��1����o�Ԩ�xx�WYl���=�����Xx��v�q��!�w�-Op~�C�(�ƺSU��g�}m�>:�11+�H��G�}
��d�1⳥q��Wï#|k@�+Su��F^�z�!s%��*R�a�%�5�d0���m�4P�=-�%�j���P��Bkp���L����󥅢�g�_��d��Z?g�PH�_��q���Y��D�B�UF�<9��9+���y��4Y�x�������+˜��x03ff��� =���1nr5l\Yf��8��0�T�R��@f��V������uD +����Ĕ���{���`�A
χ"�e����L���37�wP5=H�CJ��Lt0�
�|�����zm��`�:�X�mx��v��������E%߫Uh�����[v\zP��R�$���9۱(��uD<e=�st�h?���lmS�c*%��3l�r7��	$�6�;�Dvb@�������a�>�)J�{��fi�;�
c匘�o�D�X��Z
�w����p)%}�qm�kT���-�ٻ[4r������I�נ�Z��r<��U�'4���p��U�D.�G���+Y"���'.���͗�P�$�&��N�f��+u֜�3��;�g�:��s�IZV�-2ࣝ�G0���O����o�7�h�Ճg�)J�_#��� �,vM��<,��4��k����k�l��N)-L��q�����N�x��S�������wX&ߑE��W����IfM�����V �8�I�?VNg7�-K��{��)�Z�k0����IM���^\+ �H����s$��Ǽ9cέ����ᶵؙP�K2"��c҆/G�N�h���BJS,��UO
W�z0B9���U����qLmi�b�F�j�����X9�4H��ۖx�[C�w�c5���{�x.��q��l���R^�	�XXs:�K�Qu�[�h�V]���hZz���7)�\bW>��\Hz�i�����鋧n&Ԟ�?�O���.��L�
���^����K����\�@O��
V'(�چ�����
Ja���j1�:������[3�m���S]ձ�`^�&o�V�"E2ˤb򐡴El�>�!��~���@�r���f��6��]a`n�&�e�{�{�+U�z��V�\���=,z�����7`���G��E9����+�C9��`x�e S�l�X�Ja��>��icLS�#9��j�ɝ��u���	{2fgt���q§9��:�h�������ج^��j�/*�#��#@7���P.�߹�'زǸ�qW�,���o����J�dZS�;�7>�7z
�J^����Ѩl�R1{�u�>�|�8�l;�V3\�A��@]xO��q�)������R��� -�UB�wo��*��D���]��8~#�[�5j>��_b�S��ˑd�WT�*I�n�l�_�Gu���ϲG�=���}��ݜ�c�e�a�9|T��=��:(�D?S���Vjl7C�@���NoTC��P4r�]�>-�H=JxJF�ۓ�^�C$d�K���]g˪�U^c���J�3�8\��[d�gƓKR���8���fkog[JH�����|,l�ŏ���S87�"�ҹA���V��Q����w ��@J�$`�OŤ;���oɈhb�ޗ2�ܖy=Ml�� Q<i����D5��ƾ��nt���6��8Ǟ=�jl�� �v�`)KJ�X��
2.�~���.��H�Ui��aL
Zm�4�2����j�� �s�Y�%�g��
�N��:{��la�t������~���&?OM�(]��S3�t�������Y�j����I������cjb-�l�@H�^�����禗�Ks�O��~yS)���Ԑ9�獸�e{ra������(c��H+�2�E�����v�J��+�����xE����V_�H;�+�v�MW]�4r��䛁K�mM�5�h5 ���q�	9NB�sy���Ȗ�6;���ϣxL�
[���B�y�vR'����7�ڭV&̙N�=�x]�#3���r��
�����\� �7a������Q>=�0�f|�1���g""����Ċ�t��r��,(��6�Z=���f������b�g���z��lߙ!a%?�ҵ�������N3�a!��ļ�x�F!�僉���$3�@L�K�,F�Ů&50���x'�H�a�Q�e�a��A��-@/*���Ʃ��w�7�h$�-p�*I�����F܎�l��DS����1�/r,�p��KBp]x���1���)�`OH�M�I��"����t��3����[��E��t+[�}��p�2v��/C���e��w�?��A�/a���͞�y6�{��6MA|.�fT��F�V
�iT�P�-�@����Ñ�^<.X���$|Ҡ}�v�z�R�~o�ݵR�9�UvOG��gh��wG<m�֛�]G&׿jt�ic�7iF
�yr�|�����T��������.����qN�̰Q_��o�&����7�7�U]��4����py��>�6iEND"Mά۽A��ф�v�/OK����;m8V���r� Py��wug�"��.IQZ����0g�����d��������`N�@��z�V�6�_�g����>9h�؀o�eu� �v� ��j�Xo72���V��=�5�>z|�W��'\u�Su�9ţ��&	m�)pSJ��~B�	�1!�Ztђy�
f�9�{�"?�	��Q��n\�5��2��g<���x֞Bm]KwБo�QQ&������;�e�`K���M�&��_�V����΋_�ô��f��̿u��s��4����I�23�3�-Zjo8�:�W#cD��$�����ҢK`bUq%�����څ]�x��l�</4'$P�ƕ�%��Xq�%� �-?���dN\'��PEXD�?	W��0܆x��4z/-J�ߖye�I��@���5�N_ZW��;�Hg��>��� -d�HvK{���:�m�7e��l�^#���H����'r�� ��i�"��D�&��G�56ʵP�c�{;X�ge>UbLF��I}ɛ����{�'�w���<ܫ�o''�m���_��v戾��t4�B�рt~�����3���n�ݪ{�֖$�f�<�d��BA��Ŋ�	�&�^-W#}/e��%�� X���H׭*��
�O��e�=1w��0�UV��o0�����V��S����#����gҽ���M�X��-ds{�5v��菉��h��ceOɂ@����j3��px?C&���~�$��۔dK�c֣�#�E�1>N�F�uc�}�4� �D���g4ǽe����W2�.cθ8�fZ
;?\,��u<{�`�A���w��.�<UprJ�V�̧Ӳ� �`��j�(ժ]�{�E�����.�M���ɁDD/|U����$(]c��P����o<���Hx����e��܁�1?����C��Pd��b���?ޚ[r�Z)}g(Ak��oYz�7��v��Z\� �G����Ug�B����#} z�&w�AS'j_Q��V�S���+�i�#�X�9r0v�8x�]"�H�<i���Y���"+x}�F  �]6Xt��i��s���(H��55��<�-��� �6����^v�?KN7uF�+EŘ"%���Qb�ћм�fwK����8\�G�z�j =wx-f����)�ʢ'��J�^������#�2 �I��
��n�g��CU6=����ƞ!�ly.��q�4���ߩ�4d�ӑ8���� ����R8�� �b�4}��+�7�[��@�e��IM�y�����|]�_0Nkg �r���EyC/��t��q��#k^#7E��L��G�Ň����&k ��e�������#44 N���$"wp�vd.ۇP��sO���g��=�L�h�l�w��JI�7������ 5�"��In~j�	 5ɇ�)��{�L���Ra�펐i7OXAP-�Yg#�0�`��0{����Ǘu5�G����"\bI8n������s�����9!�zg�# �Z��ЃD+LA�i�Kl�����4��N��H_}����@�¬n�� �����P����7��)����cw'+�+���/*㡭�O��?���uQ�G�񈫖6R���<S���~��0.�V1�.(�V	�)Ga�P� �PN�Zh���(8e	+	t�"K�J��r�L�B`�$�v:&n�jˢ�(�0�I�NE����A��D�R\�#��hn8�Y���6M���fQsMʝ�8'�8lv��7W\������h�7w�[�p�$�y
,	��.[~�2���UY���LȊ��j{�gj����S"�E��mȿ_<��`��h��Oh�t���s�����\��|������[&�f������X�7���A�p�	�7l8,�ɜ�!h��-��4XI��X�-e[4�+�A~���JG��xؖ,
�7Om����q�>���M�3��j_�v���Q����LlC��L�c��QS�I�ӻ�$����[�V聑<A�jU߻�OkO����u��O�l�xv��bM�0Ԝ����H!p'�_�^���zP�C���
��*N����M��&A?<	�B㏡�M!�=�R�w�������,�XX塌���k�Z}�~#.�ϣd;�k��m#U^5�_�V=��'C�Є(�ӓW��{e��Z1
'���-�iK����0������Y$��ݿ��1�+�\ ݊�PUuUt�	n�����~�A�|h|i�	�
�#	c-���$��^@1��� �Ԛ�o1���M�;���Rū�-]����Y'3�D�v��� �U�wό�a�Pj�즂��l��D��>į�x�LcֶA�:��˴��9x�u��S3����"Q��D�<��C�NT�+y���v QyF}���.�S;Ę�s���hcL�;7�ׇ�>x�t�;��d��J��7=fr	�Y�S���[��KU�i��'����uu�{�>���+0�f��ͱ����V��=Wʤ
��R
��(]_ikW�V�����o.)=J=e3��	��qI	��7kC�g��Y��_����8c�H1�'p�6k�����w�������_����2z1�"*wEDјH������vc�U�^4�Ok�� �W��HT�z\r�\����h�pЁ$��2�ڜ�^_v9��;(b6.�Ze����N���ҮW�61��c'��V��f 0q�I� �q�Qr�L��P� �K`�p�������?b���$>���7e��١�,&.
m`������_ws�ĥ�� g���7��,lo����Z�����XΗ�oّ���4h^�@@�p���fXf�2>���[��L��/�"�e�L*��V#�V��?�qX,^DT��]]�uO�5�f�!X?��F�i	W�	����m��KZQ�����QxiyG�aFg��lbSBJ��:svVh�/I�û�}��2�+�o7][ހ����5�S�w�6�K��
��h%�5��m΂߄_b�䝥K\C}ySXnP���q>Z*�dy>�ae�T	��eE8�%1w�dȅ�qy����@��8ʌ>���dY�1S8���A����c�)z
��)����^�DT�  P�}V�3���=�fy��ӥ��ld��$��CE����Rmo��-!�D�?naT�vm��9K��4M��	@8V��r��#�=�ߑ<b�+g!E�/'&�pB P���q�F����b��و�<Sas��L�')s�8�� k�Smv"�Ȥ���� �*k�H4�9��$�֗1z��-{P��K��$(��I؄=�ڂ��Q��������%t���H��X�@��2�.}����2�o[���fP6GF%�g�|`��~M՞�-x���@B��m]K����L�A\Q1�'���`f�״?�5����L�8��G?n?2w[{����"��f��L6��갳 �:�+�Z@B����Q��
��Ln8�鰳��i�{�\;���r�Μl���P��͡��#�6:8�{{�q���G�ۃ�7�𔌡�=y�q'����)Ȧ�fr��,�W��j�hD��v:;^HD��un���Q�B�+Ј�ܼ��5[��*�6���/8����>LH��mQ�U.U˒s�4�d~��;�'��m�����~��85�BWU��>��v���D/��k���v<��i�2R�|o���q�Z�Mfd�)Z�=�=4U�����Y b��l�]�_e!�Z�0�"�pcU��:��]p��BAsIao%u�����>�; 蔕K��?��:�c��l����MR�h$z�'�]��t�)߻�1}��ql�"��75Jn��Re���36�r����aWC^�|�U�ƻw�$_������i#
L���X�+"�kW�.�"��N��i�n��VAٗĎJ�.;�R���+.�g�kGs����Q��.6F�c#��j
��Zh0M�4��w�A����n�����������Vf��]5 �p��<GtZG9{<�lϥ^�:��#���%�{�{�f"4��܅��,3�3J��U��G�2Ǳy�=*+���f[7���L��%�i��Q��I�r-��W-LȤ.��헦6������S"��+�U����е�:*��pŨ��y�/�+ⴛ���q����H}&���*��қ��A��%��E����)l�o��珽+xY�f���36��U��!z��N�*��g����T�O�P"�����>�׋*H�� ji"���6"Jͽp�|Yk�g����!V�|&'-����I���QuWycrs�d�K�a�����Mχ�������Z�Fo,��K��9/(`g��>'E~�:X�k`�P���sM˿����jII���sK��T�(?��f����ln�$0����13ϸ��l&�N1x	_
JS�hD�m�ЦZ1���8O!��L.��!䥤�OT�K��U���ϕ�M�Z�SE8���i���)��x�N����;^�I �]8��Y:fp����ޥ��=&l���rLD9h'�@����AM�ϸq�	��QQ����t��f�?FM�p�A��K�ku<�9