��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o����\�����:=��0XɽC��1�o�~��V�44'����x�/�s�ع�ݤN�6mt����M��d����.	��r��C{��0l�d*9�{�!ߑ8�p�q��}nj=%X-�_�?�����q�w�?<J���t�>!6��������q�Y��Ⲵ����~�<��t|�:��	��	N���:lw��tf���#-���X%�w�S������8���-޴���M���sȭ)�otMp2��A%Q�$�yR�)�� *�*�
�L�ޥ�d[ַ����1����iVb+�f��Z/��n�%i�c	V`����T�q6I�Gj5�C�]M+�0�j�!<ZP���2�>��iZML���i����f,���ۉ\��f�L�����S���B�Y�yf� �(���������(K^��{�]J�&��	��X���A�wl��ߗ�dꚆi
i0�9f���~�(5^_�7���T��݃+'��Ym�<�{ݗ�tS��[���)���w����&gH`G5��V��l���SZМ���"����/�T7DF��x�w���MvEI�r�1���q�&İ��1p+��6�Ȓ���E���'t��Y�K�PK��m��uNW��%�aǊ
����g]!�~�
��9�-	I�[�E�OQ�N8}w�-�Fm4�j<7��.δ*.vA]i��(��3��a��[����tTux���������_�S��&�����*~1y4̦t�� <3�y�`3�����;�_c�j�F���͝4Ť�|~��[P��\�$Қ���P"���Tm=�qxW*mL����:�R��C���̟�yʏ[��冷Kh��}�(�9���X�H[�?�篅���k9��1����'Ç�CL$�^�M��
6�bp�<�� ok�A,6��PZ
K8�&7[�q��~�~`e��s݇ �q��:�(O8����/��N$��������������n{r%�����Ð
߻����"Z���^���7u'#��X����?�Ԃ��k�{檘�c=��![��`���!OG���5u�W���-�-�'��F�S�����t����}"�~��͜�`Es�̑���W>6:�wo~bA���9�>E��:�ϳ��jp2�_~��ꯒ������t}`G����]A_])��ޛ�P�SU0Q@���h�4�I(�9t W��K~�@G1�O<{h���T�^�Dl��#AI��R��?ݦ�[r�a=��?B�V��4O� ����%!�m+S9�~����s%����x�ʣ��*Uٯ�V�VF�l8ˎ��^!���By7�\�Kx���<Ų�>2�m�f�=�9��Q��������lEa��A	]����1̿���*4�I�+'�o��/y9n�h�t��k��ΰ���"�V���Q�XE��M�|��*���`Ĺ��/�D���cZM%�T�2�Y���*g�m	j'_�խ� ���>�=�brUu��������2��BcѼx�s�'�IK�g�ޘ�p��C6a&M:T 2����d��;<�L+�X�Y�0f���֧?�-�ϓ�tjj��:�@�bmX��X�=��P�Ѧ��+]:~���C#��������5E��h:���N̮�h�H��o jW����4o��&�TTss��p|^�;׏�z��*]蹉06y �l�_�:��h�X���{��<ɖ���-�~�P��w��؂��ߡ2S���͝D;7��U70�Z��B;�3�<�F�Irݏ�R,ui@���Y���^[�9ٵ��ך7����mLU-bA�����@��NQ��tt���o�5&��4��
�;���i;��|�,`��s� ������G�{Y=I�"b�1�ٞ��;!2�ȗ'��=��x��&T�1`��Q��,���a�|�8D��)ճC�Q7ִ\O�h�/�(�=�-�_jĨ�T�/���7\����2���(������\���
���v�Xh��J����%�6���e\4�ͷ�.S|]~���o��`��<.�<mG�����Ȍ���B5�VXT�t!B��Q@����ѹ��[�$��%O,R�'[|��)���IL�?�v U�� �<�ɛUi���Ĳ�<F����ɦ&���uQ"'�¤	���x�������ub�4t^/�-�ߚ�b{%nx�ى�<����1��2�>�]<Y�d��{�dGv�#�̵�m�|��T�1(|��R��+��}%�Z���֢�&������-�k��ճ����fr^��,TMzfWD�v���}w)�s��_�GNp��Y�_�"������%ɠ%�a/$�Yf��^GFӋ~ʳI�c�Ӊ��ڼF���5�%Z�"�Û�0��<"�Wj:�o���������<�C^rQzNh��-���ʶ��_`�fM�d��J����;$���w� u�M�z�.�%���d0�f��a+N4��G� u�Zl��s�l�|�l��9��%j>YN�������3l��M-�E�^���K�Jzt�� t�9�j� &����N4��+� ٳ�3{��;dP���Y���te��,�]���5)�C��Dm�Z7}O�!Jt�sÂ�H>DZgo�3Z���0����D(Ss >�g�i�U��8N��\�1��Nx�w�4��т�\ A,�I��i��V��� j0�>+;t��{f���T=�%�׻�'�%��b���(k��}x�t}�I)c��NC
͓1N�
�G���X�E���E�T(y�2�L�K�1��~�Z_\hH;��d��Z�]�Y�E��k���0CCH�y�K7D��bØ��e8,�,G��61� �*x��gx�#�T0k*�N3��	Oy"nF�z9,�;˟��}�#K��lCa�D�_C�+�ڗ��.�^㣠J�ks�vZ�;,�u>�G�^�=$k�B,��0��*;�f�T�M1e|�O�I��*�I`.M���)��ғ�R�U>Dyې�IL�G)0�hXƺw#b�a�*k
 �;���p�{I �QK�ǘܸ���(�2����v�X�V=K����y��{o���l8;߅��v���I�ò�����"[(2�G�w��1�yj�:�?���9���#�t�]e�\7��
w"��L��~�@��ME9]pif�h�x��^��y1���5�13�hh&w�>t-|г�bF �9�V"�#�q a�ڎ(��E|���aA^-�L�ʹ�̗�r<\���7�h��ۋ5%�P<��u~:��#%�V|�W,�s\b��1�$�Q4���'��B̴fF�6KÁ�X��C3������������{�=��+%�t��|�p�q���i�`<�D	@fV���������V㽟9-&�9�w�e+�J�l{g��1�^7!���Gv5Qt}�R [G��V�X�m"liS���y�:IF�=��+U��n��%y�{�J�A����p&��lP�+� ���بW��_�d�^�Qn_�R� �%����iT�e�{�6�Zf�4	�co�Ԧԥ�&�\87U�8�/��ޭ;d��ag*j�4��y��P��Y����.��8��9k��[@�F$�wԊ� ,SV\�Sg��Y����o��(ѯ�>�����T� ����Yj?~a%��I��hd���Z�<@\���f;s��t�$C�*&|�/�-~�4F8$�-�g:����9�سL?�Y</�~�������`�XXB�]yF'���Wל9#Py]�t?���͝hzVa^���9�q����97�����y�r����<��$�!�W����]�߿sR�v�<��Y7bQ0(�S�Bj���&�
 ([$�!H�<ރgJ���.�*�z�����vpKĞMF�:d��ۉ�܋#��}@��o���mMgFh@�_􁖹�R��u����maSN�(�T�SEξ��ŞN�y�� .]K�tpo�5�\OU�ke���AA�vS��[����������I'�������Dg|(ǐ��JU�ڿ�x�q%ضBW�x�3%H�m�%N�7[����k+�tJU[D)��M4W>y-Z�c����s�N&��WO�G�@/D����D*+�7X�..���+|�x��03VSxY����>��	Am2\-n�SuLI�Ir�I�4�us�*���j^�N�F'+�8AnyQU�(*�;��{�X60%�A[g~t���<!�Є�s��֍�:/�Q����XKY)w�p���f�Q�cN��}�H_x5�*���N53� 0{�)n>%��o6�jǇ1���W[�p��s3ß,1�V$�<>WNJ�8n��׀�!(iK7?����)�F5�$�{����b�|��ǃ~E�������B/	�9se�-?�ԡ���^�����y�g������u��]�p�5y�w/�ڌnKϡ#p�Q�=@�d6M���]4�ҿ�Z6E��58��&�-�(�ݵ�d1]�QH��>�6�Ȟx狾�*:�Ȏ
��28�7Yʳ�0��;|/%�S�:e���,�*�+���ҿ�6�.������NV�|"�Ŕ6e��ؔk��i�E���j��;]���;�	�ŕ.��e+
�lީ��2׀&��{�+�����+�(m�Q�i��U�%ݛj��b73@�;���P%*��WXX�

�[�︓U�Z0�f؉NB=��{��rL�\�9�XW����P�=������a޿IFv�+�](Uk�4%�����7ב��[]�����f�lSP%��9������P7�6��Ǎ�0�>�ȅٓd�{cX��A��<�OB��F��	B9��K�E����뇿B$k�$Lz95��ܽA�C�EO�U+�Y�2�Ӓ��	C��4#м]�5Ϟ�;g�0"S��X���jF3{ՠ��^s-�j3�}l���N�%y����\�Ne��{|�,�����z#"L4���	`���y��� ��2����v%�	K�pw�3�	�};�17�Јq�Զ�2��jO�������|N.y�Bz~���z�s_���>�#VL��?�����_w���{�J�R��A~��n��������V�0��w��Q����N�%�Z��j�P*���~���x{mF�C]��;P��(��r!I�DS�cSr@e3���q��ߐN�e����^��
\���O��)�%��A���\��=
ڭ�w�X�d�:��aK\B�{���-1�B�CeZ�h�=Q�뼵@�[HY�N~�#�ܑ
�J�LJ�[ݒ�h� :�Ia���o��*����8rd���0���D��O&� �����2t�R�w��0Rs*� ZZ�p�jRYa+�Gܭ�����h�,����l�r0D>e����Qa��J�T�L��G���pny-D���3K�]fQ�:������O�~�%:&_VNk�����W�&ӱ��3��&:� ����{��g����a���J��A@@���5�I�gw�|5�=S��7��®G�h����T��Է�YԀ�h�Z�t(R ��{�Q���W4�W��p���CCΜ<w�W�����
�~@�=:���X�%ʠ�I�B��]�spE!2G��z�`��ܔ�Wl�5�t��.�"����s���)���&�;r,�d��	�t:<^�B�Pi�֦��Nv�B�F���|�K^#��ۀP����~�-`��Ļ��e��/��Vc�(	�����>�{����1B����H��s���&_��V�F<|��y�����������I�?`�,�O��BI\j<�b�Mj<�3�'h�:+��+x-(1}�Dh�H'�@�Ѷ�07h	JyR��s�C���k	X�χ9h���p �^��&'`�������\��lM�?���[�$�5�F�RHO&�-`Oq՚֛Hs`�4U�Ϥm�_�e��|ٹ�v7ɜ^�� ��h�B]}Y`A9~7"��@	�m4�N�q��PE5�a�gU�w4�"�V�3R�v\Ia���3b�+y�U��E�����Q�(�,���z�i���q��ꉂeǻ��=UEKx5�����!	S�Y@��ˆ��I�xd�/4�����>�8���%SL��=��K�}�ʛH������б+%̸E<"�Li��~����c0:�6$*FoB��t��?�N�$3�Xn11$-����8���@v%�7VX:`�G�qJ��]����B���n�&(�W$�E�V�71�f~��ɤX��?�_��P�&��i�%���p�}#�Ӂ��r ԦҙP�6����QU>��	.�It8������-���T�[�Z�Cm��2%�V��M�FH���Q"��j���WZ���}�S�)�����)F�oCX�d<R�@�D�����(��,*�=$�Ҝ�~����n�uβ5]��/��N9���2L�����'QL��� 6�`���+bW�I���r1��V�~�e�}�dK;]2�P��4E���btG-)]�P���gG�6(\�'-)����\��D#��p��Fv������=�Ӆ���ڡ�XӪ%�kj��z�.~-�k!U��IS0���#�G+�ӎ����'��v��O�]��G��8˵`���bꪑ�p,4Ζ�weՂ1��=�*XjN=��_�3[B{5p��f��`����̲��n���8�i�����&����g��&�?f,6"���5]X��Q�]�}���)�-�N�8�0D9�@� ��Fm�0E�{�Y0��|=2�uNb
=�S��-�
���ҖV D\�T�ɀBݪ�^��V�ޓ�� B�P&���>�rj�}���6�	�Ex�K�؄�[�	���V+��fL����}�p�\�ҲB���WuR\1��}j����xТ;!r�qȒ�Qy�<��}�.vKD�!�qo(5p"	*��]��+ w'�b|ϩ>,����= +�]|v�ڬ�,@��ɀ�����V���\Q�Ϣ�c骾����Oa��pO�\+N��c�48�첢p�����q�3DO�k��Ԋ�^�e$���h9no�l��M/-���A#���0$;M��i֙��X��|�%d:p)�y�=z}m&_N��(�a�Ut���MЕ�p��/����	d�
(��[6W`��6�*f1�0"81��P�.j{��EÂ˾ "�f���q�6�����!�s�OD���dI(��Ƕ�Yy�ә=4�s�莏]��K��/��Ob8����k�-���ɸr�rh	ңl�����|���7���m�e>O�����= 6@]�ῢ�S\��d%ˀ�_���?��3�~���JxnAE��P�R�~���sC����<�3[����[����D'���l�U.�PQ�7�m����،�^��1H���}��Q<�Ro#/m9و:8���ס�s"���mGբ.�^���s8뢵e� �#rwe�:2}�P�L���ڌR4޼���2�����S���H�f9x"~�' ���h{D��R���W�����C�!��K��JԜ��s�ς��o�<�"�K�!i	Q�5�~PR�G�f�g�_�OH��M�\�����$�ESdٞ��������A��90����8a�2�H���0���9Ż��6��A����?[(>/16�ZKy��<��]6��z��>nYp�g�0��f�B(Iђ�`�2Z���RnIf:�d����^ۂI�+���}K�qP�_�� 3�S�I�\�o�����q1Ֆzz��wNː\�AO�����˹�l��0LS�2��ڠ�H�*�juw2=�9��c+�^�&ʊ��;���ce����n��c٢���	ԧ'��n�9��H/ｒ?�,a�c��Y�?iL��~gY������ҳ����D�yHo��@�J�
����tm[-(O�S;���+k����W��"�|"���$_��q>0�%�y������s|��B� ��(_7@��B+Xz9��Y� �?��Ĳ'֣=$�1����\B�ھ8܄��wy�O�1J��ρf�0_Nd3�t˧�njF_b�M��+�oC^pW�C.��(�����`[E��i(�����ӊT����υ���ms�}��H�5���
���������#�X�u�^0����o���M�������$C*Q���ك=f�B{m[č�)ph�BUΌReh�nV�R�wY�8�{��ZU��D�Ǽ�;ɇ�����_6�T��lW��ga��QH~���\��l��)�9;k��R{|��A�����v��h�K�7��/�|��%�.,*�+*���f�Z�� *��R��������|��1�9�qAu8Q:%R�����*�ٚ����|M��E��ц[X�(�-TJ���"�T��%[A��&�P��j{+V���L[b�1�	����ec��\��܋XK��=�hT�ի��o\���1+��' ��		���-/���$E��'�v/o���!b���lp�P���w���L�Wf�o������&��!���l��^��̅|��Q��R��l)�(�R0�&Ĕ�C�S��z~7^�+%-2���ތwȑ*�^���7�r�ͧ�<�v:�����g��1��#Ƥ��&@�z�b۷�";:���T6Sm������.�{=��OAu�m~8��R+�ᩐ�w���E��\j�V`����nR���hͧ�F)�Ǎ��gC���Gs�t�ހ'����y��q���YC�5�_Z}�i'���H��gr4�t�'�2/�y>�k���0@�7�M�H��bƉ�q��NXǚ�2�����qM��3%��p�O%�J���^}g	�T��TFQ��w� d�tuЯv��v��%w�<�b�/7T�d\�gƞ�?� �2q�a������X_.�
v�L�_&�X����2�\���ʽi`���'u��2�8֦�<$��X�|b�^ ��G�S���`��:0-�_�+�y���ŏ��u4��{��b�p�Mm�"Bۺ"�$�C���#����epbs��i�;ұ}�@0�3��P��Kb9A*}�D�8�k�O-S����*���U9��A���̶a��2V]n�H��_/�a+�_�(5ߦ��n	M����ӿЌ�w��݁�&U��s ���Y��M����"gu�!Z��#NCӶ6c���Ϻ�y�o�"���e�0h�&/��\3v����L�B</�Q��[瘑e�����"�r�B�����^gȠ��7y��:�>.�Ndq��@��0<q��Ŝ-Qw�?!TŮ�\��H��ct����V��i n�?�9��HB���L�U)�1=��������U��u��mrh�����kۈChq�;��k�ِoW�]Ya���%�da��T�}|���e�G*>�T�)��z�Pc�������I��*@v��'.!x�3�r�#����I���x30WV��r�<�x�*����p)�Ā��b��W.���A��do��5�?:޹#3���H���D��K5sS�]��r<��Un�0��]J�Z�=b��e)s��rD0���=�
�GG�<�.�k� \c��������В�1�eM�֎'E��2hM����n�>b&�H����O��0`_�8���FT�~�
�U5��.G/y��:l��w|�&r֣t\��8٤� ��9l���p(���׭�	PN�p%t�	a�8�M@HJϕ%�b�ħ�h�R�^�uN0�9z�%iR}A�M���1P���F��>� �����p>�L6�z�P2?v�ȁ��r��~Lg/�WQ�W5�;������D �� R�>�4��J<��I'�G�6T����@��!��*���zU��.?����*INx,n22K�,�)���e͠���^v�:.l�!��ܔ���&�g/܏�l��.��4�Q��9rN5�3�X`���KS���  �y���ƫ�Y��xh�z�y'��c=��@�kM�Kc?媊�~G�C�\�Q��T��h!�w��B���s�MD9��1��B��:	���x��
����1|e��6��Uy�su�����~-C2��P��/���[�Yh���ڝC�ɓ�$�,���s5	\q[�w5O���p�<�`nu�v�����bV��#}M�b���]��%;�ǅvCU0���9����	�}�M��x5U�I�n4'7)��d�̭~
�>.��˳�0�w�����e�i�=�p����÷�L���^�x��=����e��Z���a�TǱ�C�JB���m�
�|�o�/�	L5�11��z�>�A,||m�B͌�o�Z��=7΅�l�u��:J�C�H������4
��ȅ�?�b��<m�9�_�p,�{*+3ȧ�@#���畻<k�tAn��_9�zv�=��*���P��a��عNs��R�iJf��k�Z� ��k6J�{�mI�g{{Ч�8�hфkftp)�?��u5����%qy�LL��RػL�w��8�KArD?-:d��6*O������io�����x6��B�ɜ�<��-�~�~]�5��:m&����A��JMb��"��b������ppa����S�lA�qtn�_g-X�0}D���0���;[�!��ř��rd����TM2q>���U�D}1ډzP��~��K�4]��c��,=�B�{4h���z����9O�U���a�A�xp�}�4/��,��j5���E�ڔ]_G�����ե1���fކ��!o\�ޤ�0���~��7���fN.��.��Ӹ%	�CW�*�I����1����J_֖�?=ݘg�[�H���g�,��bA>d����<�#J\F�kSK���T(�)��<NF��nu9/D��c�)�q��;{D������j��:�%��w+�AΎ0�a�/�8@�y5W�ո~'O��^�s
;4(�ܣn��`�`��\������ �i�R���r��7o��{vQ?2^KخSb(�r/!��v݇m{C��	81�n++L8�6���&U^ at�ӭ���x�)�|�E�$�)�UH\s�s'��~d��7��d&^]�~��y�^��!1�]9X��2\iQ�MN��z�/�P5N�W��B�d��gJ�R�pÖ�͎x��������υ���ef𝐈��X�RbU�	�Q��*3�n�u�w���~]��l��g
IUx�쨷�:'E(X�c8�t���#OsKn�������n�[�,P�I�%Y����#As�
�����Aw��1J�P���xb�G�՜U�&��h�ZK�.��"M̓&ӋCt���s*Ec���emW"�i(��.�m�~t�ws���&���	UxXA��BcS����]<g}d���M����8{�d��o�D�"/}�oL�Z����eWf����L��o	6b��/x��y���F�ᴓw���4��+®WN�YGc��OyNZ <�Q�PW�D��l��f�Y�;�0�<=�؏Sׂ��z��B���:�����&�k%��������C2j� 1����}N��R���E	r>���W[fP��x8(Tk����P����p�ag��}���޾1%�_�X��xt�Ґ8�zx��S���b�-����\�6G��%QQ�lFB!@Y�þ��@�����8s�ȼ��>�
����P,�L���S3���#C�kر�B|叽1�v�r�5�\�G���E���J.��i�?�݀ Xr<�C��1� �{o�Jk��a��G �FCzǙ].��B��֣/:rfυ?FY�d��e���5T��[:'cɤg1k��K�T'#�77�-60/9�X��G���3�� SPYt �	�X@���O�D�v�i	�x�����C��X`���1�e�t���[��Ez��:�����JX̼er�ñc	ఎΘ^/��zkS�+f,�+m� S�`x0C���rM/I�-F
�+�%X��ٍ!a-3�'	5����X;�e�Y�mM40���`�}=�
�t���xx�*q�|��,�qX��qG��gҖ��A���_W
�KYS���j��ʼ�r�f�sWv�<�W���5FSm-ly��m�
����eT�D��(n���1�E���R�EqW��i#��������J�L�W��@9G�{߷���Y�A��w9��2�@Q-��3�ޅϬ/v�Z�#�)3��>�蘳���W��c$L֛����B���dJk(��.υ�c��+��va)bKe��*&G	��x��q��c{4�.��-�ߎq��B{����eמ23���>�B<�.u'�	����y/Aa��{�DI��XF�LX(�����X��*��)�R-y�B����ڍe���_1�ê��8D���{�j�J_��QP��?�K��U[�
sh��ǣ���1*u^!�B��0�^�Y	=<�����KoD�E@j1t���i2��x	��_|�8]��m�q
�%�wĴi<�;�Xmc#��و��B&n��wYrHuIj ��*kc�����r�����,O<
�[ Կ��: e��^���i%�t�S���W�G�Z�Ur��l@�-ʌk��c N/+�!�v��`�s3�%+�6r@3Ye��_\ X�Qr��~�?\NZ?����G?�INQs�e���?�9��`#��2���NN�V�&O'�#?��%����kV�D�E~�+d�D�_��"�����g�ZZ�P2������/~�F �yK��������]f���z�C���3jjX��"&GW�;�3���N3�ubգ}�&7¾и�#����/04G��J@��b"4��٪ug}JkC��/ٙ�;�ꏏ�P��zG����ֳ6'�NOl�|��U�}��t��Y�͘����_�%A�酊uK}Kz �^:��D��ng��h�{a�t.?�*�؛���ku�n��p1� 1 ���(�aG*R��"�v��	�O�;�.��ˊ��2�COK���o�c*�.�	��qPO�®���74�@�'�P�53��	�S��
%��xP�;�a��!�~w{�,���ꦵ�$��"e�z�oK�6���D�?�U�k6O�0d�#\F��o����V�q�����T�;TK�\�;���N1<��K+(ô�Č�e��g�F���{m�jK"Y#����NY����P�� 6:i-U���$��q��x5"�-/���`'�߈;H��Y;k�Y��D��������?g�릜����d��З�/Mr�������S������v�
N�UᠨQ�<A1�çYNE�c@��Wr$�o�HaLgcSQ]�I��-�Ea�������9��臬��,n�29_�^���'�H8�ؚ�	�M���0����P���F��	����fz���%?m;�S���e�`:$eR�Jεs��a-��b9�"�w��,X��>̎�vxO�̔�7N�~wS3�� �X޻��ьI�ʷ)�g/*�g9Џ���˚ཙco�Gwdl0��H��e���(d��Rb}���@*���u��������SS)�q�Z���&��+���B`QV?�z&Bv�������Y�yAe���
'��l�#��שfkB[��Fl�@�T��D�l��0���;��?9��&V�}z���Z�����ȯ�,e����b����>�!;��Z�d�
 ��Ɏ仝u�}/�.�zSA*p��4�Ϳq�y)9���Ј�����jҸYĈW����g�X�Ǽq�B�R�ah� �����*်ym@���2��:��Q�Em�}���ɺ�P@Bb�0l	�
�������u��S�V�'���[�M�}c�UA�S=K��Q��6�m0`|�8Ԑ��.C���Mɹ�6,v껖$�	�V��}�me��s�r>ypX)��1�<u4���n��s^,.'���������:\̌�^)U�?L�Mps�.n7������zKuTf U��$�s�jO�6�ϱ3�҅����h|��Q���핝ŮX��]��J�Nύ,Ђ߶��?�"P�&zH�^�\+1�6H��ԥ���'Jx϶E�(�#���c�.j]�4�{҄>�Q�Mm�"�q��=�B�Z"�R�k2�a����)�������v%٥If�8���(pg�@���W������)�7�[�P�M��?���'�q��7��;Z�Z]��͏�ŊE�'��q�^� �Q��0!���e�
"�vdpf��g]r7@-�G�*t��Y��][���^�,�!�Pv]������>�o`\��ݜ� �Ԣ]Tc��m�`�0(4�����X��N~�~i1�2��[=�hR_DA]lƣx�+���͠�-�x�w���9����8: �Մ��s�2-��|4���6*0���dX@�Ix�	6��D�5�lA0ԋ�H�ޢ�A�G3�0���zf����1{�a��xc V��G���4���d��I�U,zU����|�M�N�A	��ѫg� ��Ӽ�W�����������ݒ�
�VJ��KU�hoӤ�5И���K�b�	�{���乭����$��}/�C��WH���G�9Z�o=�v;��y�J�Q����=I�*�[#`�^�H�Q�E4zrb�x���gw7��W
�_�V��f2Ϋ�ֻ�uפ$���uOB�	f96U4a�2���%�vv�5����."#EgLM�+�˖msT�EH��W�0SN}^��܃���s��q�S-O�%�ȝ}�~�N99�Iw��Gy�����Ǿ�R�	.��.B�V�.5]�R]�L1�b*<�gu���2��I�/��\B�a��ys�	#��i���9�DN��W�����f�X�����ީt���n�x�!���T�;;'�����%�=��il�soW��[o?��W���f|�����#_���{>@��v{uڕ��o:��_����1t�bK�M�􇓃u�ˌ��v�I׿�Bo�.h�N�c����]a!�e^�>]��$�|W�.��ĺ�i&E����݂�C�_u+�dncya�{'�8ۣ`o���{�g�I�����������7�B9�k��������y�9��$ԠS������=<�&��{�lw����熡k@���D�0��^UjBB�?�}�Y.�b"Jۥ��r;C�ݶt��ԋ?���V�@#�zR����>�<�fo;�^�LI{�#T�^�(�rۚ���	~��+�P8N²x������